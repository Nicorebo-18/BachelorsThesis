PK   t~�X˜��[  �e    cirkitFile.json�ks�8�-�W��_v�D]�淙�3�mvg�m�l�CU���)�dKy��~l[��R	'�Be�5w�(�N ����n��?�����s{���������gano~.��?���7_�_������������^�����?~}zl_�kWu�T:�����J۩�ɲ+dWu].���?�t��u�{]�^W��ux=��4���rὮʹ+��2Ng���*\�+�y�b#��6U�y�U�.�2+�Κ��Ek]S�>tz�ݦ)TӄV*ګ�5�׺��*ڲ�RZA�[��(+_��,C�m���:�ބ�T��0��w�V�R�&TԄw��\��"����B�M��w+�H�[�B�ke��&T�k�}�ɢrս���T�֕ɳ�V2����pUE����(JI�[��[�\V
�2-s�U����ն6Em:]P��]S۲U�0<Zi��Έ��F��kZ#:�]mJ�+�g��6 DȬR���l�jى��:�r[ɲ�L�U�/w�ѡb��*�B��)��*�M�w��N���Y%]�՝/�tyS���Y�Pu�$%`��̂t��B�2�]^�z�Ƚ���Ѣ�>4<�o�u�ʅ*+Ǝz�sFԲ�Y^�0kc� �.�-��Tk:�ݶ��(B#�
�j�O�P��	��ig�ɐ�Z�M�9���� O����M�ƽV��'��ډ�8�Y�@�������mseUS���Z�L%��Z[P����&ڴ�����Rਜ-KY��u����*0f�a��m<U�/Z/j�"P�u��l��T_�[gݽ�7ei8ʒ'HY�)K�]HY�BʒxR�Ļ����?�,��B�%�.�,	�WԢ.��Y�Z��0��0�C;��
_ض���o���0���d�h��ԙ�3�+��UԻAk�.��h�W���])�҇�6����P�J�.�V@7u�å*H5.(���dȻ�ta6�`���f�k�|M'Cg�AP��e��&��U�H��
��a�ɝ��w�Ɛ�E֘����~�������hU���AM��Ί�
��y�Um?���U�ذftԻ�b((-���Ļ�jH���Ļ�jH����I
��Ļ�jH�Z-c1��,ެB���<�)}���*'��*�Bjy�G���WN�=Q34sN�Q34�Y5���R��Q5�GxUK�jH��f��f�o��[j~6EQ��D��,qA�A�d>/L��`q� tNդj@����I� �SǪ��Xݬz��f���ޘ�7ɜ���~�xX�`��s�;��!I����U5�� #�7X�^r�	�i2���:X6la�
��ڶ	J���Z��f}������[QFT5�<U���>S�>��\�O�t�$�UM���ƫ��+���W5�W���MnJ�@cͪZSzk^Ք^�ƚW5����,�V+NլE[S�;�`-��RgXݼ�f�g�c���Iiַ�vR�u��D0���6��e�JC@xem�!����lJET�-�+dVJV�*��RNd���/h�➅TCil�Y�ɐO�Qaٵ�	o�K��m&�2N����g~6i�xS榯z7}��0U�<���F�ˬ��K�	�jJ-A>X��gI����UM*4d��2;,�Ϡ�Y��R�:�u8�Π�U^Ք:�αyUS�:~�U�4��g�O�la}���n�|֎R,����lJ�@&��t�f�F���p�j�L�gS�2xUS�2xUS�tvʃ8e(A�ռ�I����,��)}�E���!�RhPt/$��gPP�jJ�A1h��)u��񪦏���{Bc�5S E�U�����Q5R0�8^3xOb���S8���h�HS;70�z��o��0�����I�<v���hr���wi��#�rF��ƀ�W���V[��#]F�O�ש�2$5;����ª����q�ᢃ.�{z;�k���3�u�8g��:� ��2�fe�M�=��z���&�:e��
�����s6�N�%R�L9vsx�AWi�A��pF-�P�,�Qk&x�r�A5�(���2(��Fvߓ�:�	�NyB��g���\��5�ƛ�w C�USn|4p�Q5��gݳ�j&��ؽF�Ԥ6آk�L&}޶�Ɋ�*2p�vUYzͬ�t�#U�F���U�·���j�y&��"Xk�EA�2�(yL��j
f���TM�����yrC�20,�Q����Pմyrb��g`��XU�}r���vÎR5{J�CU�}r���D�N�9}Fzΐ��>�_�8w��*9s��3����y�C����>#�+���a\?{����M�X�����8�â��8}F�vH�t��D�;l@��쌚%e�����@�Ǩ�Q�!�� �WS�-�Ljˇ�M�:Q��]�q����k��y'5^ aܵ��uA�=�fJ)���}Dad��cˆ���0� �f�����t72��q'Ɖ��H��o���l��gNSqr s�#2X�0� �����_�Y�,Y�hInY�s=��`�R���EH�A'x��QC2k��i���ir�������w�_ �.S���C�AU�1G����+�u�Zz}�8FK˱��(J�\{�PF,��S��˺�N�⑚y��953Mи���M�Lf����VSC ���Iv5�c]P�cpb0��S�
����Y�LޱF0ƪ�$�Ajf�6�n���/������+rq{��5LA�^kC�fi�)d8:��m�a���:���S7�`��9�.g)2�A�fM/2������A���6�ĉ���i�k�&�u���Q3���������X��&'!�j�(�o�:<FI�Ѣ����$�>B^Fz� m©�Aj&c���e����,�k�5�ٱ��Yئ�`Ђf�L�`�"�[�RE`�&NլNc����3d-H�0r�?�衴ќ>gMOҐE�`N�3)�0]Lx�U�Q3����c6!�sD��b�j5��E�<FZ�e�1J�paԬmDr=`�$�$YfO2j&�0p3LBjf� e�L�̓�A7b<t���%!cT�HxcI�8U���r�q"([�z�60��.W���(���(�Ă�Q�;�N�S5yb�����Q3��h�5S#�1j&��1b;F�t|�:�с^�㛠�iG�:�z��.hV(�}����>�NPջp����8_�ҩ<M-%X�̩F�J�\w�~�y,y��rY�ĸ(�n�n�їS5�
�����I��1r�&����ژδy�2��/Jجy�5^haZ��j�Vz}X�>���t_?}yz������͹�M>�Ǹ� ��"�������R�_�RL���$�����a���R���Jq�l*� �y���F�ƈ���]�r����Vs.��4�:M1i,l��riF�F�P�Ùb!Z_X��Pܙ��2VL"�F	�4(�����9GQ��[]���)�4y�)���T���D���К`2��U�hH�079�(�oq�+&�)��ꨋM�83\u�0��ĊP\�&�+N1�m饭9�(.L�+��$*]�P�TD�:V�Q�-�5��u�3������Y�b/����h�t�֤1��KS̀�R�MÙ�z@q-l�sV�fSg�R;ρ�9���	g2��.辊uw^,њ�N��.Vu[�>�����X氷���8+�P�z�V��P�MY�v����}ˁ�P\��5�V&�V%�V'�v@q60��:�boK��4���4��bt�e��e@�s��9o>�`�9V1���{^kTܸ�֫Fq,Q7��te�9s�P,��r����K��|���;�ŕ`}�ϓL/�L?�����8�ƫ$����(�����<�F32�oX����[;4O�|��9����_<�GS��UѬ���!x�����R �.l�������ӝ�47Ms;�M@3����}6A)��UeN��dC[���	��6�-���^�Q�fn�o��5�QW���X{k����(eq��$�	JY#4���ӟ���n�VP.90�ihK/���&���cK0����9C�ۂ���M��9aK�i@�O�Д�	�hq��,��c�fܜo�x3A)��Nh��cTX_��f@3k&(�.y�ф��!h���(4e
��L�Kb���CλQ�\��n8o�K���@=,ǯ���
Ms8�3h����F��6�Gp�wќ���c4��|[�,	JK�Q4���������BS�-X�`����%���n�� �KP�X:[B��-�m`v����c.4��B��"�\�hJ��U�̖��E�>�0m�-h޴y�́6懦3�?wF3�͟ߠI����|a�@p�c-���5Ўf暏U@�l%�"�4	��W�ѥh"��SL4'Ղ	旚�4W�|$;��i>D��`~�٘��ͬ4��&I�?<G�����h�_�<D�mAs
%hˢM�3��f�YX�l6��4�˂� flY�"0��BT�G͉���]0h���,����Rnz��O�E.aMIr󛰧�=����"�CS�,XA`��2̀��X4+�|d��b~��d�c�&��aA�H��	!�� 4A�<�Є		JY�Rh���9��`ީg�������`a���)���F��?��`b�ȏ??'Q��y����'��ŕ �u��b�R����l��r(s�|pʂ>��2��V�����i|��Y�����D��{s��{���s/�"Q��_$J�=R�_�_���6�(+���$�^�nM/����	�hq%@I��������(���J��ϯ(�BXH'��R�W�,��G�(a��ޝ'F@it�'PF܅1�m���1���5e�MЖc��T(�����:v�r�.xt@���Pr�;u>��A]�.�t�	JY�Qr��,ޚE�R�"���P���,�XQ.��9nDi�	��t�jfM�Qn�_ ��3r�T��\0���-'��s��̶9WfΜ�,��`.\v�0_Ky����R��\N�����s��0�QNL~)2I)*I):I)&I)6I).I)>I)E�%o�4�i�+� X�A�Ha��"�E�4(��tp�4(�iP,ӠX�A�L�b��2�U�4(V�L�4(ViP�ҠX�A�J�b��*�u�4(�iP�Y�iP�ӠX�A�N�b��:�M�4(6iPlҠ�$�إA�I�b��&�M�4(�iPlӠئA�M�b��?��6�m�4(viP�ҠإA�K�b��.�]"7[�4(viP�ӠاA�O�b��>��"�aNL~)��sb�KY%��_�b�����R�ыrb�KY��('&���~�91��,�̉�/e�_`NL~)��sb�KI�/�� ̉9[
̉�/eq�`NL~)�csb�KY�6QNL~)�z��䗲�����R���䗲8F0'&���1�91��,�̉�/eq�`NL~)�csb�KI3F�k��_����L��D�M�����3A1i ��sb�KY'��_��(����R��Ĝ-��䗲�E0'�����䗲�cC91�-p��_����Ĝߛ����R��('��E91��,�l('�|�����R���Ĝ_PNL~)˫ʉ9[
̉�/e�^�91��,ګ0'&��e{��LP������R���䗲��D91��,�('&��e���䗲l򢜘�R���䗲�/0'&���~�91��,�̉�/e�_`NL~)�K	ʉ�/%M[�!��_ʢ��䗲l������('&�����s�f@91��,[A('&��� sb�KY�0'&���1�91��,�̉�/%�-j)��_�����L��D�M���#Ή���4 ^>�91��,��PNL~)�a('&��e[��䗲l�����R��U��_J�1Z�WQNL~)�ND�3��7z�W�3A1i �6����R�w9('&���5��_�r�ʉ�/e9D��䗲��rb�KY#��_������R����\8�91�� �  '&��e�ʉ�/e٣�rb�KI�/���_ʢ�sb�KY�aN��K�4��aN�Ť𲍈sb&(&����pN�Z/����pN��,����r�3��%�O_������|.no����~������������i�o>���<7n�ct�?�n��ʿ��Yrj&��Q�5N��,�GT�Y��5�j/:�P3x�x���˺���l���j��P3x�z���+�D� ��vU�HU2!0��T� � ��U5���e$$`TmYUs:\���`|�cU��j���^B�A��Wqw�f��5��{�&؅���.ءf��b���,9Z���h���d���A��=����A�=�d���A��j0V{��@'`����Ic��� U�ߌޚ�a�F��U���U�3��Ϩ�\1AJ F���U����Nnl9�sn��,۫f�C9(#�7�`��jz7�j�c��A�=6��-�b�$�ް�2�X��f�a��A��f�k�a
��$�aTM� {���=�l�4+��I�dat8�� ��I;d�a|5m�bT ����	����P��h=CͫZp�Ԟ6�1f�g�>����� 7 +#�g�d#����ءf�Qc��AΊ]�w�[�f�ƿ�C� �	i�B�G�M�����I�	��l��vT��8����
�b,��W��O���DȮĈ�$a1���%#�w���]Vk�+6�[�ao�D%�.7�0�>�{ ���7�׳�Z���>�� ��UC_���%T53 ��2�jp^n��]l~��h���S���ub,Ի|4H��ǲ��,Q��ȕ�4i!��L�ez�� ��h�S���ݜ�I�$�^3�LP>Fջ\]aV2`m��g�r���� �Y� �[��L�ɃM����f޲��fr��o�ĸ�85S(�gD�*�f{ʹٍ1�l��>B�P�0�N��uG�݆20N�x�3�Bé�g����0b�A�N��8�9��&�@N�,^�(�����=Ԝb�MG!`���}#:dl�x+�i�	F���jr�A�+�W��d1���f(+��!�&�;�d����{7ʙ��x�r�c����`��c�h�\(��&��rV��f�6�Ҫ2�� '�_v{Պ�f�rU���0��/�)U��P2B�xW	|�T�;x�AzJ2��dt79�A.KF��ȽՉ��79�D��ib����s˨�&>a��x��_-f޲% ��?��&�2XRuc�߷W-���Ψ��P@�F���U��d�`��U3��o	5�M�a�qe*���#����T-XZ��P�\��B�(�.�*����s�ǧ?��}���H^��6�=�^�+g5�I��o ����.��l8�	e�ݭ(�n@9awk J�o �!v��D��5 �ݭ(m�lޅ=��.��lޅK��.��<߃Y��.��lޅg��.��n��:��FD�gw���v��T��YF #�n@�iwk �O��a����e�M�&i�~}�z�����v�>@�l����v�>@ym����v���r�o ��v�@9ow���s7� f��m����[���巀K��o���s�c�֎Φx�;�����L�4��=H{�#&wo�0)|w���[PB��6k ��~�U��w?/2��.�~����w��Կ�x����lޅx��B<�(�;��=H��[�\���{P�WC��wӈ0���&�=x��-`�	��e淀K.�o�cx�وR�w�2�� �xx����;n�0��6J �~{U��x����6����&�;0��Sރ�x���[�G���.�1\2c>����Y ��~���x�MHt�ߢ��w�������x��m�y��\��k�;P"��2#��$�7�=x���F ]�~+Ț<?ރ<��.��n�&(��n��(�2����0��g�>4˻�4-x����1ʽ��&3�L&f�Ld2���e����� &K��4|�f~����'��@��o ��y�&y"g~�|�|2i��`�;�I�A���C���2�2?�� ��.42r��-�B϶�]ȡ�-�rDӁ��S�1��C�
�>t�	��e�N�6pɳ4�ˡ}e��D+q���K���	\~m~�4��pٶLH.�v�&p���M�Rp�[�e��͛�r��KEy����{�sӖ��۾mr��;���.}v�>@�d���`k��%m_�'����p)�i �����X 8|.ync ��i��Kj�_�����p)�i\/<�fР�i��U_ۿ�~�������S���,���@`� 1N\'�x�T3�Kr(����C���-�u8�(Ҵ�}X��-ಌ�G!y�n�M�&��o�{�᷀��f���{d�᷀��f~o��j�`�����C���wH`�߭ 4��~#�t6�����q�Nn��	�7�7�s�������K���|~��S���y�����|�����P�=����K�������������x����s��B��8ŉ#(��q�D>-�Ci"Ĵ<M����(fF�<.���`��I�X��}
xǺ�8E�gAt
y�bݙB�s *�ꜫ�%�2�љ.�Iy,/���z�>�<�?0��c�o
y��$4���LI5�򎳨)�EÝ*2X_�%��3 g�D��Q�t�,�Mg@�Q�z:r΢��3����vk?�դ<�:������������Z��q��,�Ng /
��k5S�[��2���aS�[�67yV�tI0���.	���	AQ�c�M'�f�	"[_�
���/+>y:?$�v6�$�\��<�ʛ��1z�t~H�xpW�Lg�e����Y�\d���.�B0oM��h1�X�Y!X�7��U�t��L�ǉ��h8q��\���Ų:��3}d����GV^|d��X ~�u
f�G.�ר� �V�n��4��
�G�;0-5��l��0<|$����L�����ذkK^�����;07���j�n �8����-?"49)�4g�Y� �9ig����Q�B�53c�MƎ�3)���;�������
	/�s�aቓ�B)x,�rR��ǒ�Ë#R�܁:�;(&pf�����D�ص��Iq����*nf��񱃲^Ό������1&���)&��tb�zL���?��k7r�IX`m4���N44��y�G�5O�#6Lh�Iy���SEE��)j�-�i���3����G�fZG��F��v�@�ͬ	`c���L��!T��ׁI��=��u8B��|����``Q�,T��ׁ�aG�Y=�����Ű������EK����KL���=�����:0�5�8cw�c����S袦�����¢Q`�W�H�ۋ�T�Ix�B���(��7������䛍��Pw߰ԥI?6�!��Ü|,'Mj��(�9�u���D�h߁�<'K,(`FH4tL�8��h߁IH'}GR`.K4��u���>�`0z)*F�C��>#�ә*��
ׄ�e��9��.�w�b�;j���vо�Q��S������b�6���F�@���q�C����@���C��Enb�'*��+�2J�hX�L�`����rrGF�b%Sf�&�,i�M��T�;�/����#&#DGL7)�����&�V�)]���g(�A�����K��~g�AF$읅�H�;1K�|��X\�ә@ݍCS�L��L�gi(�5��ĲQ�S�-�*"0��jň=�xH,������03ߤ8N����Wvd���INpG�&�����	˶	ox��I��Y�@��I��9��3�����0�b*��4)��}������f��7�X�Yt��9dQEf���XnO8��N8�X��)�jpRa���`��X`�V8�˼
��b��&Z�S�td�ۣ`&����;�S��&�Q}��e�GK���@�jP�L;��u���n:��[;.��Oyx'��Hm'�q>v�wԭ��?8���� �?��ޟ����g����b&�+`&���� �0��	�'ڂr����U˙���[%�.�O�cuX���ت�L��8 �����@FV;���,wD�ә6/B�q���*�wY��u��f�QB���oo��{hz�PෞDa.����M?h����~��P�l�����py�D<�4�l���!�~�0\�n��h��!�{�x���!s����p�!Fm���x�!�kP"m���!8k�2�e�����s8�΢����g���a/;�@��ϰc���/pح{��=������2,��N|�#}��'��cpU���G3ع��5�E�=X���3 r��0we�z�b0	���o�2��t0Ë�@�E�J}�E�>y�E�23؟�n^�Q;[ r�s� �n�l��T�6T�܊��r�����rqc�rb�r�`��?y		���ĚO^BB�'/!���K���o9T5>��8�8ʀ ��H�^�E$<-�"9��b��<�{���L�"�1���Ԅ�
9�m/�>O�^��;�� ��� �W��A.��� 1������'��>�����~0�ۗޖ�{��ß�y0��N������O�]�b]�]��'�9�.z!z��Խ}�^|s�Q�q"�8�Zqw0ƜC�����'9'h3�.v��x�}����}���cӊ�`�2��!�q&';�.Fq��n<�����6E������%����MHN�'�)�.x9�u�0��e;1r������1���3MU��m_\�������"��n�n_����o��	�پPQJ#�ݾPQ��X�����#��x�bù��Y/(�^e�eOI,����p��P����/Q�/aeo�"ޱ���/�ė�$�ۿD�Hk�5�,v>�K�dg�����qZ�)i�'Z��3Zc#�)8�ጔΧ��S#g􍋴�4�1rF߈Hk�5 ���nC���0���� $�:�|Jك̊��Sd���Y(��,�R� �%�5�iB){��њn(e2�noM�F��sanoMD�JJף�4��&�JJ׃��5������ �(�5�ER6;H���5>�bI�b���њ��*�'#�J�t����,S�R� �(�ob#E�b�l��7�eJR��Kd�Md���Q�EF�DVME)c���9��R�2�2�sd3�(e��2(��JQ���d�&�J����'J�D���C��A�BFkb3�R� [)c~���R� �'c~G@�)U2j2��#(֔&9*}�2hJ�tqGMMib���1R1ܐ��4c�Td]Д*��;�"\S�d�c�>GCib�>m{�d�g(ER�moL�gH��ݱ�Y�-�;�1loLD���ؚ���G0cHs�z�ޘf��A�-���O��� ICG�6��� ��o"+���0H�蛈�İ�0u��\ƚ���TL֜rH�HŀN�9��N�,X�D�Kic�M��9�XJ�d<����T���((�sbCE)d�A��;���R�[etNl�(���2�&bVXJ#�T|�Ή��Q&?��"�w���X�^����(�11Z�J�<N��D�ᖵvr済X]��tr済�R� 5#�'2���A�9Fkb��1+�C#"6�#�u�9��r�:��ַ�FF�
G��ai������_#q�����*Oi�5����*O��X�w�#�!Mu,�����z�\5��1<2�icH�5F'���O�1��Z�X�/�hz�{�1�����)M��1̭����������j���进�7�޾|�W��q|$����>R�Gj�H��#s|d����>r�Gn��������<������1�q�1�q�j1�lq�l1�nq�n1�pq�p1�rq�r1�tq�t1�vy�v9�vy�v9�v��������/r�/��/r�/��/r�/��/r�/��/r�/��/r�/��/j�/��/j�/��/j�/�u�L�E��EM�E��EM�E��EM�E��EM�E��EM�E��EM�E��EO�E��EO�E��EO�E��EO�E�j�i��S��i��S��i��S��i��S��i��S��i��S��i��S��i��S��i��S��i��S��i��W�:�s�3�s�3�s�3�s�3�{�;�{�;�{�;�{�;�{�;�{�;����L�Ş��N�Ş��N�ŝ��M�ϝ��M�ϝ��E����v�����n����/n�/��/.���"�mq�>s�>s�����ܩ�\��N����O����O}�}�O}�}�O����O}�}�O}�}�O����O���Z���}�ܖM�T>7�������o/F)�ɫe���/e��o�O�~��>�<����>���7%C��^��+4��c�����͟�/����_�=�������	}��������P�������������Ҿ�������ms����{>������_�?��sM8;k��������c����|}������⇰����l]���L�;VX{���w���.q#JU�Y[�5�v�/��ҕ�P�j���l4��}�6T%no������ �������!�R�{��k_��s��=����;s+�Ѭ���Q���R�㧸���n��G9+���0*/�AL�^N��y��9(�OZ���д�~x���������oĝ�S��@$�H�N�4�E����6���o7ڞpxx*�?���v�XA�N��.	�D�J�7� �g vY��5^Ph1���;=b-2�FWE���k�럚�{�����w������!�������1���fΑV� K���M�վ3Y��U.঳��4�)@ZP��B�x�_�rGէ���7@�����������@��j����] 
1�ohX��������ߧ�<�>A���	8�?���To���Pv���T*KE�RQ�T2�?��34{*��OblB�36b3sĒ~z0������l�L��?��j8j�U`ӆ�t�� -}tm��D6���-��Ȝ+�η�y���*�����M!J�2F时{�b�w�[s������j��?��w���9}ڭ�>r�P���q+�	[���wVj!�����;�ra���y���7M�to��"����Py�]���ѵܳP�q�6O~���zGŭ��� ��iqxPD���R������ۥ砜8P�)+G�Cg)E���w�F��{w#�%���#v�Vg秿�d�	g�w�		���f��g��c��|����=Ac�J�>�[�C�3�$��1ο�ĝ�u'�!F�0Ga�W�v�1wak�''���4Jv^:�����sY���S�ȼ""��F%�w����<�'��rp�989�8jOu��܅J�'a�bZ�����(&O�#ʘ��{K�=r�`CI���NHm
m�f@�PH�YN�F1��`�8-�)(�����Q����B�#�t���0&b�Ԅ�����8ȝ��^�"?Z�N+��l�[�l)�|������e��N��U?eE�� J���>ya�Ť���=�]!�9�p/���:w������
��]�慱8TI�b�A W���#!\q>v<���c ��t�@�\����1����;aN�6~�·����_���M�{�|B�N�}�ARG�ۦ�h��]����U�蠬E��I����PVD��U�/=V;.������SD�����.��<-9���e��A@�=H
�0�~��渇.n3%�]Xs��\��U�a3���5UT��/��	6R�u2�����<�șTo�r&{���?{��쟽#��IMN���9�q��,���s*z|���s���&?<��l��R�d�����J$L���y_hi��uAU9+��݄}JY����MY���ehE\�f�}"׃/���K�S�U�$���]�u��q�W�7;�bo"TS8�w�i�6�}�Y���pw�Ȱ̸��zII�����푉qp�T��P�"B�iF��G=�Ο��g��x-Ҝy|Ϝ�f��o�����gR�Qʱ����ȇ��֟���W7��a�v����+����.��e�h46`W�&,�E��]ЃMX�*Q[!��D�"I�([��?|H@�o?U����k����1
d5aG삁t*X��wtE~�!KY7���m�δ)���M��l���Jl�C9�����τ4��;TH���_�Oy��-������%��z�$���p��3�Ē��O4Y����T\x���^���w�j"Y�H�{��a��Ҝ�b-z�Yku	4뫶h�*�mXht[���mfD+�2`���B$�7b�n��W�E����ah�;��<�?���]��O� &Z�ם�^wa����/�����W;�hW�M��3�E�e��d=��흰}��^��<(39<xR���I��vwt؂�i�3�E�m\�d��,�v��lt܂X�qs>X�����`���G��2�"l�w�ܕ&l)tоa�^T��;�&4GVؖ���������yX����0��Zʝ=�}V�)�~��o�l2z�NL���A���Ƕ�Gkh�H�-U�ygB�<�:몺�d6
��|,����Ӄր��E����񯤤<\ y�O��z�D�%S(�w;�C�`����9�[�;�{��G�����;h�S�������Z���y��'�\o1Eu���t���W]�?Q3J�.�\����]We�Ct�IU�<nR� &U�S�I-mjRR͚T�L8x24��z����.2h�5��D1��N�pg�����:�S�#m�N�M�ki�pO�#~�ύmnf��0�"�z}r��*��Ta�目~��s��4��������C cX��^'���Ln�ڬ����",Z������WJ���I��~��㠱aɎ=0EN<p��r�)M���
��B�L%��]�?N�r��;k��>S���'�6$Pdr.�n�x�����hà&ό��m���)��X]��������qu��s����)��V*,���p�x鯋Ϊ�9d�G�)��+ˬ�I�Е(1C�B�:u�#5�=�}�<�-�~Wg����������Ù��o�&s�b<�m�~wg����m���!����>�۞ɜ}�=�.w�]����w���:�Z�����C�ǿ�����w}��:�]��~�����M��'ǿ�����w���.�~?���o���������w���*�~W��w{��9�]��.�~?�z�~���������w��{X����g�۳������wy�{���,�~���w{��>�]��~���o��u�ۜ���~�g���ߏ�u�۟�n�~7g������������:���~�g������G��S�+�`E�vO_����o?��Ǜ�?�|������Ǜ�o�ᗺT��Ly���%�U2h�`�vJ���A����/OA��_/��㻕�\Q��e�iՕY쩬���դh�w���߫s�'���v�6�a�Й�;W�:������=~��r���m.Sg��m����-�>�.��{w��o�{��۾�}��I�}�o~�Ҝ��,ȢȬ-T��P�׍��ᛀ�ҶJ]t�o��秗���>���ڪ�}YtaԺ"+k��J�ֆ�;v�e)�����=oM�OU>4���?~
�i�?�&��p*h�������c0�<�a���sO����z<�x��s����l�����俟`r���O�/��4��o�g�������t݅�����l�Ǧ���\/���D�4u�%SP�Mת�R�sm0���hDW:F[�����}aa?��)�,�}��\�vm�M�u�A�$��S�ʋL4��/�J�.�l��ƅ�h�V���͟��O�ڗ�_������~���ӧ��?>��>������ɧ^����s{��������OO�<��������}yz������1R�s��-_���_�;��헶~03������A}���C��#H����t�C���qwO�òy�׾�eɛ�3�4��r�SuY�]��邆֒��O�  +�L��Q�A����Q^P�N�hO���'>�s���;������_�(C=�Cɷ�.��w���X��h���y�!J��?�oFk;<����(�a�G��8��ãh�E��(:Gq\�M�I����Z��Ϧ|������S�\�mƟ>�,
�_G}XZ����!�0:ug���7��e�ZʢgD3j8]�m���������j�t�͋0�M����`��`V�CӺ�W�����
��Q��論ϫ���0 /O��n2 �{�f���o�ч���v��??4/?���=���&��s;\��|�P���_���uTC���n�~���s�����|h��������S��_��q1,ʿ9����|~����q�ߚ)�PX����%��z.����M��K��}}zx|�}���PV�G~�����}���"�������?lP^��}����D/p�2:*u�J��H꧿;6��$������+��7 Ɗ֭��Q��(��u4'b6:���٨�r;�¦����բbڎ>�c�ʯx5��h�/l���br�ԅ��:K޴�.y猋��:�7r	�3)%�Uc����@����'@�p-�
o�UQfbX��><0�ȴ+cEӮ
� ��ԇr��J�XѴ�jq1L�}ڨ����ol��z)3F|�¤>:b�0�`:^�k�vU����F�6&�]\L\P��bj ӕ�㊦]hC ��0��� (���$�ҞoEӮ
��"9��	��r���o$��ZW����*h]Ѵ�z(������Ѽ`��~M����k�gE���Ovq4�yʙ�$� P��묄+�v]���+�>>�c�oě��/��I�-BZ��؇Whw�M�*f�E���T���V�Ãl�9�{�l�����g���sl�hq����0u%e��i�݊D���~�X�	��v�s���a���]/Fs"&E]g��] ��@C�x��M�.�^)��6#$/2s�bh@җ+-u+�v]�]�ԉMC~=` 9m��M�*0.��P�P�0��P�_iiZѴ+{��4�ň5G8hi��(,$��ܠ+���ܠR�C�b�.�%���J@[Ѵ���i�iȗ���`�^�FƊ�}�g�s�О�	b@冫�؍Dl�������\Ѵ�Z}gt��R�/������<)WZ>W4��S-�5��d]��bB�������֮	�\'3m�2�J�>w��jktm�&�Z�� ��B�"Z�֭=�^�CZ]c1U��F�%*�GOB�5M��&����ʴ��Һ��*ڲ�RZq=��h��**L���} @(��u(���dy�XhE�V��c����&Z���ڢbq��[��y^�7�!=-��p�v�+v�����y�D��Gb��q{�,��:��|�mH2�5.��`[ѺkbMAac1���-��*�����|u@Ο{}3޴��D��~�K4���)C�>���-[`+#�z�� =�E�^��q���S
巈93��>k����Ub�h�UAty��O|����������#"�u���2b�����V1"���r�=�(�~YѴ�.R���Gy��4�X.�;;��EITNŉY�bt5�%赔����M�z���h���4�=����״�1G�2r6��׎�]���n��/�x5�P#�bŀ]�\q굢i�8�7�z]���9͉X�^z�5Q9)��W��e���`�b̮���e���QE:��{�!�Mx!F� ޴T+�����F5�H��χ�h]Ĥ�X� �̈́��+p��iW�ń�D����8��c�Ї"F���i״�P���nAi�ALb�A���bM�΂��iWE����9�i<��%���m�Ř�w��\]��*��i`R�* A�E�zZӾ} ��!)?�(���R	��&�N_��M��9�OĬ��e���R�`Xԗ!��ԯ��Z�|oĮ��^�ˎ�5nPԫ:���HC�Ʈ�4�i�5��>ͨ���gɕc&�K�� �:�XѴ�BCj�@c,6D8�1)٥Y�}x�At?�ڊ�]y�g ����b�A��4���:�M�P��h$���3�K#�U� ��vE�>hIV��X0��2A�_h��Dt�h�G�����*Ί5ޘ�r����8(!��
��i׵�uw*��q��4�}t=]��rEӮ
'��ˑЯ��rE�'�!ZÚ�
�Ix��%�Y�C�J��Zp#1Eh\Z���it-�B�A�o���]Ѻ+��y�����&*�c!b���V��&r.5�◫��AS�� ���j��]AFl����I��#cE뮉e��k,F*��6�X�f�(�b��堽��Թ��Ԋ�]���袥r�ND�1Jj��}��!v�:Ω5m���~|Cxr��6*w�LD����[]�,t�(!^�
�kE�R�Un2�&�\�;�6H����� ���$n7|�tj��_j�L�e��d�->�B�ˤ琔�hc'Rq�4E�s�R�$4�d�k�im.��f��xA�Jŉ�G�HU?�೦S����L�2��i��@�c.�%C&E�V��&Փ�C�֦S�2��a«�*��ȴw�ն#����!�K!��S��E!!��ΘR�&�YoU�c	�p�c,�~l����a!�)
oN��0*���3�Q#\�N!Ow7�'�I��B�6�j�0.b�-�j�`2��[�J��j9��#���+�t	�u�!O��&u��6�ͦ!F#C>�>�K|L*��i,�#!�|�M^W(ƐȦ��]�1�mɖ.��W�y4�w^���B���P����B��)wMeR",�S}Mx޶dN�m�0�FBq��/4$$�����JQk��[�hK/m"�lK����mK��ܦ�`���^p$E������D�DɌzD
�xe���X��x+�mK��6�m"���K��z���p,%T\�]��R���j�fx������0_�MKŰ�	�c�:K��+�E�ŝ
���} �
1�<}� ^$�U�D+�vU�ҏ�����ܯD�Vjޯ��_�.�` #��+�6�Yl"R	���*fEӮ�aF~K*PtL]	�P엠���D�=��H[Ѵ�D:E-������K�*��0[Į^ӕ�F���k�B|Lf+���"���y�Ue�5s��C�8Z�6 �k������N��P��~�{搀�|tG8��ňLc��-�&%�0�6�+W�-�6N������༼$1A*�1Q1�!h�����Q�I4������%�ƅy6S���;7��@1��1J9]�����6��W#�h[2xl�s9�1��ɘA1�-U1�����)���o*j�M�MK��m����,�ZZ�b��2�\Z
�u�4���-`'+��mKv ��h�Tܽ .�����HQG-r�s��I�ZlB����W�-ζ��c���S\�aR�E��Zl��p&6��ވ�i/jQ�V��s��t�lV6����
_ض�.e �]���m�pf7m	9
�!�;\zK�qT�"
��\ _��e� (.�]��Qꛢ�l��V��|��ԙ�3�+��k��lM�d�m�`�ɪ����q���l<B�_�
���؍y� ���7#苪��v�R��e�M��4ޕ2+}��F�]���`�k����t|���FR��,y�I�n�j���~ű���ֳz��2��]V��gZ5Nm^��9C�
�lEے(�1�A��]�h� )J�=�3ZW�uy��Z�eޛ`�QeE]���M]�>w��I��5�>�%[7i � ��({�@Vץ�(�0s��$%����r�C[��
��2�ѥ(�ƴ&�	S�۹*��?E��Z�T��pi�h[2m���A�C7�i�����$Eh��`z�8H�kL'M�URa�V۬rm�`�t��2�eZm�b9\Ѷd�l�r8�6F h|-�&k�K�n`Hh-�DYQTe�u�gU����WycE蘤Zc�޶dZc��7�6���{���<P��_��R;����b���f�hM�RQ}����L/������+�B_�@�L�+&,�}f��|�S�N�ǘ���6:��)1���>d���i\*Pn;�bH��9�e"���QŝtZ�¬���%�}L���Gh�V\\ӶT@�tAp�݈�Kwyh�I3�h��;�J�;��u)�0�h�V0��i[*mb�i"aqQwa��B�ŝ�ꐰaf�uY�����°�_�[א(�h[�Q�tg/�W��Ց �쯋*-V�Iq���]�Gl�>�>D2#'�j�B!�hZ�צ�ڼ�wښ!���sw�+�I�Gba8�/&l���2'&F�/b���_����ȠT��4��IM�u�-c+��2BiyN�;�MK56mCs2�b�e.�	0#�;G2���iT�jZ(�xB����h[*�m�
Y`P+0�����q*G�E
�Zkl;ϱ�6�P��oW4o���,�ۘT�۩b���Ȑ�G�ڷ��U)OVV�cEے��l�C��B�a=1szh"f�����3(&���˓>DH�p#_	��s�"p
1r�ѭ؁�h[*8�m[�-Ǳ��	mAFb�F�Dޔx((d�$�Yaůh[*��f��@4�++����b��,� ��7c��.�U��6�����8��B�;=+��t�ƇS�Mb�R��t��� *���l��8H���;�5��xے�7Q	��D�D�&3��I�{<o�
��y�D��*��uY@a�AF��*�6WV5u'�֔5�[�mɖ�Mv�����p���Z��(�.�s"?U6��s�X��_�b*�I�y)b�y.B����cKԊc�mKf�o:f�aØ�J�ՀHq'���\��D�p(�q<(G��/H���<��^���E�މM@��u�[�`��n���׺F�]�U���¶��(���w�+Z��P��qP,�ra�t��ag�����}إ�W�I�roj�e����ڠ��"o򰭩꼑��4������s�i �V��j%�V@����7D��=K�	(LA���޴T�vf4�����W���'(fM��K����'P���H�ԶF�ɼ�L0I{�|_�Lzv��,l�Q�P�xM�\�i�ȋ���"�`&bĭ�I�Ǘ<=�����H��^���w޴TJ���Q'�ЅX��u������=��D,A:����v��J�LWaM��a�
�|�ʼ�ً�QZ�}[ѴT�v�at�F�o�L)V�@�DL��4cM�$B�*�Z�}[ѴT�vtr�`¨��Ѕ���cD���Qt��|��RjA�mJ���dZxے��7ݕ����q����#�>�ѮSq~���{"���Δ~�<T+ږ�ｉ�j��6�"~oKТ�Y�Q(��A�"3Ǧ1�ΈX�+�[ִ��<��>Bu�R2'�y/BQP1Qč���D�$tn9K@��)p�E��B��i[*�nRc���n�ȅ�)*&�G�D�h�%��������N�%��!kڷ:t�@�Z_����S��xC�v�8�F*er��hM��h�:��3�m@	x�ц
4���[��A@�����^�q&����^�1�.s+���h\2�G
�"04�v���'sI_rנ�k��1C[��_�_Ѹd������_��A)�.� EnW'	 1
�B_(y��x�!�iJ?�
�nEے��6Yu�}���`�SD>�K�	XNC�S����H�t���~+ږ�ŶI���qE���A#�D>JK�Q`��L@����	�]��ؚ�%SZ�L��V�J�4����4��k���|.�3���᥉��n:�)ĸ�q�0&���vD���~�a���;�m xW�*C����0ձb!]Ѷd�mە��f��O#� ��رVc.VQ/C��*���.|Z���b���c.�q��X��nU3��Ť!t������� �^��&e�Pj��8b(Eؙ��<��B�7�ǎ3�"~r�e2�B���&��)OW���8����[���:^ �(��Vmn]�T�}��-KY�	;�Lk�e��6���uY��m<�%cF]v��m��Q�)�l�Y�T�߉Ȁ� Q9����gA�z�u�p��3WYHi2���Ilˬ�U���ڶ	39)�V�٬h[2mb���Έ�S��&.X���D<v�B
�BѶ� ф�r�Ċ�%C�&"��2����r�6H�xv�!/&�"m*���#�N��,�!Ǜ��Pgⴔc��%X�7H	?Ô�||�L6 ���C4کS!��kE�ւ�RkP`IIV/G�6�p^�i��(@��  E�:8�>2�+�5מ�Z�զ}�x��j��:#��o��c+6H��fkHW��Lx©�\��ۖk�fŗ<!�&9�����ט
�Z�2G}�h��ڬ�e���3/�.3amQ]�[gݽH��W�sk�,�v�FufC_.A����ߔ�gŤ�hm�7�%���az���%Cж��AY<v&���(&�^W�.c�!)x1+sנ�2h�$���ږ]��MWfZi��Ym��mӴFtkx+ִ�<&�D<Fa,�|�1����/V�M�
�f6�;��v������&�zBw���n`��=6�JDQ��E�E���l��B��ReZ�.�TSe��mm��t�H�d��ي�1QD��)6HI"np�bP1���rU�ù��q¶]� %�D�kE�"t�ݻ����U0(8Vq�b�&��>M����](*�W���|-��:Y�&�/�zYѺ��p�5�DF�2ꂬ���⛮�B�@�FUm�ts�)+h�S++XW�h��M=�"F�Ј��b������C�VuU��N5m]�<�klW�EVua�\�֫�(��=�2�� oB׌�n-�F����%)&���gf D���ܼ�G%��ÂSb�B���Jϊ���ئ=�U�@�H�H[qiC�RY<O����",B7o\& �Ƭ)��;(N��O�״���}f��(e����aR�3q�X��H{���H~�����Hs�Bx����$e�.O;�8I��LiD�×�w��C�5�K���x�!bU�'F���҈-��0���M����t�V����o7�{X}�����Ϳ����/����߽����O=��>?��m��?�o���ח������
=�����S��|x|�T?=>�����?��P��)�ϧ�o�'m~n�ۛ���PK   � yX<��)�  �  /   images/04ddd2dd-6c74-41be-bfc6-e572c074e241.png�Yy<�߿��B*!-b�AeK�l)�ޢi���#k� I�H�D�%$��%e�Bb�Kd��<�N��u��w��w��=���9�|������|�?�+���B�\\\B&G�9#���]�˙}��s�$KS[C��HB������YYw��ES�FG#���;p�Сr��R��N�<��\}  �����_P�������c!�z
ߚ�p/����Uj���.?�s}�""#�^���de?y�\[���|ya���SAEMmݛ��O�/�^V~n�RC�M��q����{�?���ϗ�+=c�*���#���T�@�V�����*A޾\?�� _<�,�,�Lt��ѕ�����z���9�3Ø���=���mB�m	!g	Z.r؃���9
��d�l�����v���/�ڜ�O6ZN��|VWN�熬����>ɏ(����L�`0�Z*�WMg�%��QSE���U�)��j���V�'��#Ǳ���mm`��5�JWΝL��F�U�UH~nhU---4F����A(����A�>��5�	~�d����5ޙ@֕������>����Ax_��
��B������e܅�&z��>dV��םD&������?�g�㉙ٿ����ڟlx��������D�5џ�G ��)�S�W[ߏ�'��lI$�ߩ��퓬����������翈8��'oj�ue5u[ս��4��4�0���ߠf$�����WU[�wPNٸ�����B�v%�y�9!{x�݈h_79�?��O�"�q���K������?�C ���q8*.��������w�>e������A��_�م���[ހD�����.�Oy?���{��z~޹_��x�s��WE���5���U�x���֕#�ʒ��_l���&�N�����̟�J����8Q�

�q�����1H�?���,N3��݇8�?����i_~�>�z_���%�mb�g��#S�p�T2Z��.�(_{��I�|��vs�J@�;.T�]�����zB4��`�S���]E%�cɗD�NE�� ��Α�0 Y)�,�ʞ���1S5�YE�W�L�\��:�[1���f��J&��-�[�=�p����Q����%?�S�l&,�G>,��/�X?�%#&�:+u����%J!�L5��/�S`��}8�L9a���V��u�����A��N����Ð֙ ߝt=B:5�<ɸ����c�'e��|�_~��G��=��Bݓo�ڙ��ߝ�1n� �fN��:8~��)�X�B��(�q@z\���}�;�"�CR��RŖ�M�y�Yka�[�ج���'�[�J��U0ؙ;����{Σ��{��?JL�>��r����rՀ/o#���*U�X϶��Bp򷍇2��m鋛�>���v���j����$P�N����d=��IרB<9j��vQ�a��j<j~�SsM�Dnq?Y�#/ �x�f�VI�#Di�{56����UO:��FC)m�z�;�9�:ή�y� 4%4�f�_�z�Z�[����=��*%�4��'���QCg�'̲fI�ȥQ�)���D"n����|��� �
L(��.Ї6BB"���-���@�-&�o��}6-m,���l�,�N/�I�i-�! zsE3�Fď�P²���:�>�:t��C��'Y��ւ��gWD0;�a��#�U�N��7��;��B���Y1�X���ëY��dS�l�y���GMԓ���_/_�g�B?:lQPІذ���%�Mu��v�����O�۬�|X�,�oz�2~�Zv-�[2�H�c��B\���y�3������mk�ۅ�ջe˒q������\��kL�I�Q-�=0���g8ˬ,���Ѩ���ݙ\��z�=0��|�:ֵ]
�1�����������\kc�����؏҉o�	�o$���z��~O��a�|��4�֬4`n������EqYW�0 `���5[���&)u[E9Vp'�%1���a`5�*ӮxhÞVp$(��+��]FM!+p1(Ͷn��
n'+�JB,[n�tÝ���Bb;ֹ��X_�.@�p�$%{�QD��jY2_Dʜ����n�!T��~�Hnx�l�?�(���S�!W\9�v��lL�)�M�|�R�.ggayc��i��1��rt��(���J���oYX��zϷ�e�(��J�	_���v�����d괥q��RnM:�[���-�x��#�A��������H����3�P�Dq�urL;�]_nMXϵ8v�ʗ���D�V0�M�;��,[��� ��$���w��"�����!o���Wa���X���T��[״�<_�/AW7�a���xbvEއ��I,����5��q��F���=ߤ��/�e��j�FЅ9���`f�u���)|����Z)R�7ľ}��z/n�w�����9C���+���
�]q�˹?�[�m9�m3�R�����y$6�L`��Ȍ�9�%�(*��om����ZOu|�|��&G��+�Wۡ�C_���
{$A����E�z�ƭ���ȍ����2n�X*5 D�퐧f|����}�h?ˀ���\� ��[@;������D�sQt��_N�ի�>�jLQ�_E��Ez_Yh4�¼�2�KcPM�/����F��{��Ϝ�=/B��$%���H��a��Ø]�Eܳ�Y���Z�*�q��9��&�a�@I֞:Q�#e��{�z�lDܴ�a�b�8*��;� F��񦨴�\���RXI�v�s�0�Ҍ���8�޴�5g�05�d�Aؤ�i�u�tl+�P���v�M��+XR,��
v6+��5�q���,[�
%�@��H�l�+���d��eSm���s�G�+�e�!0�y��
�����@h�S#���d@�%8���O��.v��+��\�6\��'�"�D�r��_;H��-�DJ��w}�(�>ly_w<�Q�U���"���h��%�Y(��g.���l�v���K���.8?�2ڠ�g�e�>���9����ح����(��f7���tm�E}�����A�"LN��zPE?HV��Ģ9�h5�u.�d�ٻ����2���v&.ʽ$��q}��L�^BQ�������x�n� �Spc�C�2�=�O�A�kqkW����mg��:�:�f,����`�sx�7�� ������q�Q��HΞu{�6����;��]�Q~
/F}�^M�� ��M|	¸s�j�Eq�RDN�
�-�3
�.��`U�������Hsc��n/�Aj�_	�7eze[F�*��;C�]����<�(���7~� 5ߏ8rl�Z�[�[i�y%�@���y˹M2�кz����4��<���~IJ�s�s􊭥��?��΢�[�8{u��)�μ��6R��"#d7!�_��}��.����β'�㧡�=�r >@�T^��`���D"H#��;2������XW=�O�ମ�A�(K|
T����Yr-P�(�c���*e@����Y�йj��+y������㥯���4l�L�*�ۇ��J�VCQ��5*ԙ��� �߉ꆿEH k���R��q�cs+E�<�j����Uкx�E�i=�"��e[f.�h�))�*���lm�z���ۇ�D�-b0�& ��pf��"_�֓�&1��bX2��U>�����qcc}+4wZ�/+�é�M��-�A��T$t����H�;��%b�s�Эw�G��+b��;�QVS�:W��G��VL���)k��=���F�N��q-���v@^���N	�q���,)@�E�-�w�lA~�%�XϞ��,a
�ڜ��MZ�H��ݫ����k�kdލ64�����O��WN��YfژJ?�z� %&�f���k�8(�F)-C��Be�ҷ�szf)'���qI�Ќ�:0{��r��� C��u���k�L:p�	s-���R�
e�:���P�W�q��F	����۽���ƱFz�pB�ъSH�y1*��Y{ �Dϭ� M��{d6m�����cT�����鱣�wo
uY�Cu9ws�`馠(i�n���Lov��d�~��
�J(�V^R��`#�/&H�5E?t�o�Wf�4EB^��S}��C7�{��d-���!�0�٩���ҠR���>��@�3��'�j��i��é��Kց��(����ӆR'W��{��Y�[�x;��rV�\S?L���q����k&Np�ܒ?�]��y�d��π �?�]���\'	ܐ��I����^�������Il}'S������i��9�8��)��ɬ���SĞ�\+i|��ڳ>L7�	��"	�<�v�q�a&�q�_6of�ѽ�=�B�-*# �K��)[�(��c'�.b�X: ���?:0�~�{Wc�j����ՍQ��5��^��)\f�l��k��}�#�3����Q	[T�:�EH+G
�a­�2���n�<�tIz_ʚ�r���h��pۍ�q^���hE�	����nc��<`�� 3�c������+�/��N�'C�t=���z쁞&
l���9(��ʹ}�8��F�RZ!��ć�'�g�����D�G�e(�pkA�j��a�c��a�%�{,h�rLK�-�������H�v���g�=O���;���{�=oZ<�����}8'gϸSO�?w��l5��S�b�QX�5��M�"\��w�f��ĝ�T��VJ)�	��]�X\\���<U���hrc�5Z��o^��|TL�ͅ!t�@�!�����ђ�W�s"��Z��:,�y��P�c�L?��V�RΎ��˟���J�/�C��[%�;ߡa�����j����N�v��hZH����6�NuTN-v�q�;5z�j��R�V�7S���vx�����k��En؝T��l�&m�_�eT�5���l���x�.�~ki�`PgPO��3�Rc��:u�7���]�r�e�Օ�9��sSt+27�J)[��)��jqܞ����Ѯ����>.X�>-����=V\�"�dʳpB��r�h%w1��Р��E.w\�2��ɰ�+��KTO��#����U�L$���X��T@Ģ�\�'I�7����QOs,�YUS��� =27Y��"L�cM�
`���]�!���ݨ�v���ti�ʒ�n�?D�Z��M��2�2wBt���MY�8�w�pZcUg�{�U�r�j�L}�^���V�H�I��+����Nk�X��K��^)�������j2�;�"�VOᾉ���u�hZݜ<%W�4a���~����%�J�ښ�=��g~n:��v��#�z �e��8��¿컼�qx�[ �v�N,<��9����[|��o����������|*�fԗ���C���B\_�;��g�ִsu�&
ם�5H2)��Rki�>U� �ߡ��'OQ�v7nut֡`���	���.ǧe��ח#���~'^S�Tϐ�S���&T�le5#��;���}������.��zk�<���J��?��O���g,)y^FQݴ�5ڥ������~�F�3	�G��<�ym��&5A���q����G�M7Q�9:�7c4�j�Y/G_�7�1�~]�ܙ/�]O��~��d'��j*��G����oǮJJ����ŮA�¦a{�|�<;�x�������}��<�^����5�['JK$g�n� ��z�Pʏd ��=dd�Kz�&іfi��c�,.Q�匊�@��,�Eh��MGg-�S�b ��ORϺ�x�O!�y蘭�%L��>�PK   �yyXL�4A��  ��  /   images/1697c656-98e6-4bbb-a2b4-f12a22fc7906.jpg��UPL����ww�n������	� ��5����߅���WGn��9百�����Tw=��� PQPV  !!��[��u� ��?��h�hh��h��8�88o�߼��#"��#�{󆀔��-1			>9)191	��\����T4,44,b�7������ �DbE�BAb "�"��  $4��-��!$��ވ�����濄f 2

2*�����������hD<2�o5-0݈yCS1�d��H�fa@>Kp6)9%�;��X���ED�>�+(*)�h����YY����;8�{xzy����GDFE��ƥ�gdB��e��,*.�UZV^����������?084��_X\Z^Y]���?8<:�sr
������q��?\H ��S��\��q!����b����$��1��hbX��e��$�M-���b�ӂ�X�g�I������A��d�������_`�7� ��C!HsG��)�ʥ���Ơ�ԸaꘚyD���: ��IW��0pr@b��^�c�NJ�򴔇ׯa�lvN��{��M,����ʚ���?H�V�qg�k��okllm��̾����@	�p_����}q��)ęmR�gU�Hc��g�������"=]���S�-%�R���![��X�g��+�&z��jK��8��#Kr�GP�>f�.��c5�ji�������N^L<c#��$T�z�~�#J���[�d��~���u�r�\�&�V��[��n�'��{���Fh�ó�]����=!�.�@Q���i�+/EYB��о(&1�ŚJf����	Q@9X+���HC�+p|8���_lBx���.�,T[E��JD�Q��9��>Kʜ�I�<so_*�(S��O��D� ����hQY?$�^�2���aS�;\⍮��I�/Xg�W������rTr̹�!
�S�x�E�N+�b��оg9������֊�x�# *b�7�[Rq�A���Ef�4�
�gۑ��*(>�,���;�y���u�B\y1>�D8�j���2NJ�?(�7��K��6�x���t��?O��b�X�4�];4>��>������|`3�x��_n��ɦ4�5t�@�I�F�G>:�Xݶ�5��])�+�%�$m^"��prĮ�E� ��BJ�:��<
�ٹC��ݚ��R�D�PM�j��K�$��׫ZI�?�-Dk�Lq�c���8S�V�@�a��\�ω��G�?�=s��{ 5x�K�X��͡��������U�"RvI���kR��o�P��L$��#�@Zc{�9�8]�I�?��L}I������%ӫ�������k�I��S��x�	�C����[��hu��3\�=KƝ.}r�9kX�d�l!'7l�;#|�.c*e�>�1ZW��%-ǋ�V��ٜ
�Jo��%�a+�e�%�����P��s~w�u*�%xz�	]�e�>���3�
�6�C�	F���kWe`'�.����.�ތ�mS�T�D��R5��DTT���Ype8��	��9�"0*��5�ے>u�t����
Xc*�G?\����)�@xsz�R�����"�e��������������9���������^^�g�N����%'�7�� )Ϩs��dh	��y�|?���Z���
	�w��q��l� ���a���?�17F�%K 6���$�p���K0��Mc��fFy�S�{�.�wZ�Z*��m6��X��ޙ�]�\u�E!�(t�#=d��]��l�"��`�8N=��Ƕ$��b��s�9�/�7S�1@�E#�A"?Į���V�D��d-�f��fjk�K�}�:N������4
ii��,�r��p<񠌲��'��`]$��l�)ҹN�-�]�	��~��V`�飷���Í�z�k۸*˯��]l�[iOu����/�����
��'�
j㐋��.�i>���e���	�N�Y�R��2����x�'�Й;4��<�ǒ������~9��-�[m[_GX�~@�u��9Nr����}�R�t�!S�=�o]�X ��Df�����B�>qT|�����ٿ���#a�S7�W#��p�����՗?�j����I�PB���*Й��ّ�dAƺ�ٶ�n�:[��3ѥ<lÂ��{����g$��O�: �(Ap{�B+�\͘ǖiZps���
�����[�[�rJFV�S��s�7&�G� ��de���7:��;\X�<u��O��Ha�D ��0G2����:���0S����P�E������C}΋�H3���7��P��������s���b9G(D �ԿҶ-ˋ�p��� ����k����13�}��0��ҿ��(D>���d��ݧ��������5�N����������	��>���K�6�_x�_4�~�N��h%b��w~'���|��'��B�Bȱ=���M&m�}��DH>�v���F��y�x _��t��A��䰦`��,Hl|��`Z�͞#���������`Tcx'�20�
�Q}
���Q��Ѡ�͍���آl���X���ճĈK֒,�����;�i7�w0p�t<?W
���UJ�]�jvr��O��ӥ�`*�+�s�T������[ 3�uS�]���ѭ��#�Uu|���;<�R�wr�s��ot�*�H0DJ�͌	��q�.��n2?$K�� ���+P�:�c8�1�,Ҋm��ZB8���P�y�F�W!ܵYϵ0�o�+�S��|�����m��߻Vح��C���8O/��+�v�M�A��Ip\h��@w#�e�ڟH��SE���&�o��3�P1��ׇ�K��N���+ "h�,�H�y1����ԃ�ˌD!N���{�rW\���vW�U�K��aӵ�}ŏlG�ZH�O�y���K|*[\�(�XP�!��b�O����о�Ǒt��{?�=q9VNK�
C�K��dJ�5ueM�X�h�
&ISW�[ɨ�y_1<��Ћ�ԧ�w�2M��aNov��N.ԋ�a��n3�c�qC:�|�
-[KNG�;S��Z��5�?�	���$7<���(�'j��DbM9��"J��4�a�!��.@_��L����7��Hs���f�Y��c{�4����g������_n�������j7���:���M�3��\�Oe�<Djz7~i2s�㜅�����&��.����ڥn�ݫ�M(%�;��{M0�aP��ȤKA��\�qx�k�o�!�G�.��@ ��t6wc�:�(��:
�&�N�+-�ZJ��Y�V��+X���j�ғ�9Ѧ�#oA��z+͜rϗ��c��q�_2/���tk�-y��:�4̗%�abRM2{��"�D,��ZVL�BM����3+�-|�+<��[�r��-�Y��ݗ����0�w�_x�ytD%��p����om��q�}�U�ڈ����K�0��(!&w���p��7g�؞�4c9A�_sݓ43.i�iDJ�r�ڗ�
�(Oc�i��L�{Ҙ���������9�n݊�t�s�aܒ�ȖҼ�P���)�}9[�6�6=���й���\��[�1����w��������pT�-����$�UZD��UD��wz�׷�1Ix��|�zcx�
�G�7MY��
�{DZ)�>Hȇi��֔����{�W������r0�/���:2��M������_���A�����]n�Ǐb񂋣��^��<��o��G�v���_Xw͵�d��P3���c]��g��V� H��m+�qf���y{g���Ba�O�Tj��:t$�iq8�X;��R΄��W����N�&'g�.�|n��WE�^!ٟ���1W��f�帺�(��P��5R&��4�� 
*�����S6�f��b���{�(���tC�] ��&Q>ĸ��{dD�B��.�El[hhܨ��˥���<�ğ���l��~U�R�)�[��6�š�78�k*
��W�4��T�H���֑��11��ˀ���(�ϕ��B�~��;�ɡdJA�y��9�2*>�֭��GQT����zpb��`k�+P̶.���+{+���)��7����x�/ ��k��7����}�m�s��a#`L�44>���
�-���RĿu'y𡳄�'��� ���ҝ9�?oX���Yۦ�8Cs��Sܮ Jԋ&s��1�!hz9�����8'����yO5xH�-l��j��8���ɖ���Ѻ��.�OO�?j��w�e��(r!� �������j��)|V���>i��s>����u�P�!*��(�sv�T���<h�+�D�Xk�jx!Ma} ��.�ǘNS	V��V���ݡ���]r�}�%���s�ZѨ �&7�{n�+x�'�@I�@�*��EY?x�Y��3!W�A���WS�75�-���,5���N%t������o`V�D}Z޻B ���	��w�iN�h��?u5&��o��+	�\6gPR��D�UӶ|���>��`�;���������-Mk,�,T��П�n����q�o��c�uq�'N�͈�&r��g�eC٭3��·N+W���q��'� Ump����'r��|��%���gL#q��S�t���rnOЏ�S��\z�V�̨���iE}����6�cG��Wm5+eגt�բQ�:Sͼ(��}	<���IF^�)����8[��U�.�1�Z���~u����$%B�@��3�z���ܳE�㕻�F����!ȗpяe��<:Vk1�KN̵��d>-�P�HHe��Cr��ٴ%+_veb��$ݧ��ElߐA��9 �A�
��z�?;J���ֲF��T~�f�]����l������K��ӔY��Q���^�?��9p�=����iB��S#���1e���C�cܛr��XCNDW6�^;��#p��&�\J�-U�+�7��똎��g?X�$&��3x�i)>�`�/�-��d3�������;7ܻ��Xؒ�3(iCP�|/���64=�4g/�����֠/H7�	.�k��+��P���}F��(F�g5�j;�[n�q���g��2�ۿ�$Ǥ�p�ۏB<��b�T�	�5~���Z�Ɯ� *���G�:�+�OO�a�66�4�e����"_{)��0�����.*�n������ܢ����ޏu�P���\Pvw����9����P��"[��I��Ll�oݝ�ٮ)�7����m��u6�M)��{����S&��qɄ(��8H�Tl2ߘ@zp�Yüq?ud~?�,�_0ɓa]Q�=��
WLh�WF.���W�\V��Hm���	mE�=�8@�r7D>��c�������ש.������wʠ��� oXu��F�؜~�#��e�~���H.r�Z���ʊe�,����?��m�*��Gv�1S�u��ܿwhΠ�@��~\x�u-��g�v�Z_�} .iǑDqD�1��������N���a�K0�ȭE?mpz���X�L�=�Ń�(;b�}xۊ`!b�� 8����nO*O��2�$i��쭴�?����P�K�ֶ:nc��s}=^��l�n�B6�.f�( (٩+�fۜ�������mj2�,���Y-��m���r>ph���4b0�S�����N�P��YK�;�q�H?o8R�%3=��K2
�v��A��<5×ڥ��Z�*E�Kd$J�$�l񼺅}_ �wA�(�:�s���->V?|��M�ߵ"2xx\f��=F�Z/:[��%+~S'd\��l�9l�j������VK�Ȧ�L��n���@�mPg�7\S2��ΐ��?���T���P��h��C��[a��L!���1���'�qO�ĭ�q��	�|S� ��#!��')�N��B���D��ۙ|V|�P����q����=,�d-�����0NCu$�����Z��@y�v�eU�<��\]}�]����{P5P:�c�?pz���e�Pǎ���9������zV�%�q�}�Yke�Y�9��,�����-�|����՛(��I��
����*���[���$�Ôc�K^���_��.��1��w������i�*{`���V#��6�'s�N�dՔ���Ї;r�(܀�W @k�)s��v��u)���̏�3��7��6���ba��gq�D dV m$"І"F&
S��R<;/�>5�N��CP�&S)����v� �!�<eR�tVt?���q�ȡ�Ě-",s��J�Đ?��e��x�`ZE�i�޽n�[�T3h�����ऌ�i:�D���j�{nx�!/"�O�⩫�/f`�лo\�ڇ��t@rj�W���FxuձS�5�El}�����r��ݶ��K���s��u��
8�!���*����	���)�y��h$�������Ye0XOYǤ�P	S�d(��ǭf[��	��=�Z�\�\�]v3�_�I�>�?7<q��x�#
Hۏ�7�;%��p��%������T�a>�J�jg���۟��L�*7�� 4�SEM#�*X�v���i����b�� �� ����^�9����U�=\Z�-s�66���<�6j"W��"�F)�q��A��++ذ��<���g��{rހ�ք��&U�p��
T�7������Hj�i1��$rM)l�����JHE�U��Ɣ����D����^��
%ZU6�{�2K��ʑ����k�9��8���aG���=��1gd���7��Ft�o:���|K����[v�z����"�b;��"�a_e
z���%�4
�͝G����S&���e��'H��|��q��ݷ}�j Ʈ�����,Y�xR�ٞ2�K��@y�#*�&��i��}6Ȏ�4��nL2xL����[.��X.�l� ��<�m�+T&N��;��GCArV��i�n>ar�L�&
�tB�TfH2 �0�G���+����D��#�s�F��<�Ŵ��`�O�Hp�W����9�z��t=9c�Mw?� %�����t�|��@V��&Ӥ_���n)��Ge��f1̥Ul����nT�炣m���	�셟3Hqƶ�ѫ�����%���������#Fo�Gz^�q���kѽ�9�+g��m-yT��.�����8�r(G��`�ƞ�����+�`B�-���ũt�e(
��'�Sz^��I7Lρ;�D�ǹ7�M&��['�o�t�aG[�5M�����<ҹ��u5�F��Ev��O�Q�!�C��@}�屶�9�6��lET;������і~��Ŵ�Qr�`
앉���s�e��,�/��mޏi֟.uNsc�c����
,�Ɵ����)��	�2H1�*5[z(Pz�6�)U�*�n��un��"�0��_��<�aq;�
w����X��f��U�+ ��Ҕl�S-������8���.Upǎ!�_���p=��Ԟ�8n��bI/������~�w=L(�7�*r��z��ꬵ�Q/1[�ĭ�f��E\�����T%F*�x�Px���M|�#�rb�Nh%5o}�:�?�֗^���$|�QP.�\!e�g�*ߣ�A8�z�R���-��w�+�5�d����CX��DWt�3�Y���d�豊�>��i�Iܪ5�4��f=�r�#6�O8��Y��b�AZ>�*������Q�h�?��OՒ�mP�K�ASR�E����u\�ۆ�v�e�������ߠK�2&|۵ųJ��&.�\��Z�LH���k��j�^,���S�%��/�At�ƣܧ��Ќ�%������V��5�#����t ��#b�tuc�t����.
�]^�נ�W"����/CN.C�a���i��%��� �%n�_h9����M�R�o��-Z#�i����T��qo�Z�Y9X)�w�,1��:�bh���0��.W8��n�:*,�x�/�&��p�d�N!ӵN�Ӧ�}_��¶~W��iR[�=�f��dc�X_s(߅�@����O)����a,���+ wM��p�O��b�Eϲ^e�:6��pa[S�e����?w���#٩~��8���Q��JC]�C�gG���O⯀����V�y��u�y��F�*�˂�7�]�utb����OE.k?����J�1��2���	����_�i�Bcu��5h�s!M% ڝ[��BtY�����q2��O�X�^�^�r���N�����H�7�
��2�� "m���h�I}�X�@�8����a���eC=U%�r`�e�'���R�5����?P����m�6N~�JT,�|�H�n��^�۪�\�a螦�\2Ͳ���Y�����������+���UN�����XE�
R���t��*pm晖h�KP��W2e�^�ι��t���iV@�.����0^<>3�?��MA�{V:��p�>�^_��v4�Z�����Q��1� �@36�m�� ����%��2�E� 5��H?��Ə�/�fp�Ԩ%�n��[#���w?���J�f��%=�+T@@t����;]Ս̌����ߠK���f��W�r��㕣���d�J��؟��!�a��ᎉ!�|����5�~�W�V5�	��g�`3ߔt�.��^j	��y���p����4�ȚrM�?v�^�zz��AD=	3gs}'@m)XLC�=��Pl�?��������@�e��9=��'e�1z���ƴ�F}��s���:s?�[���n�����R�KE���=���'�"�6�
�9�qi'a�O���|~�H� ]_�����)�Di�/�o�8ՙr���5�d�������d*�@CM8ꉄgA�\�|�z׀j��.�N�������)"z)�!"���J(^|�N�۴t �S��4���q���EgD��s�������])�);wΩ�ÚՉ�c'��^�{��X���gF�g@➵�%	�kc�'�j��ۜ%[���hZ}��4�S �ʵ�ކ4���p��cjMɂ�{��(�����D?���-Y��|W`���߫-F4ݭq��1��LX�h�<��"
�>��Nk���\�����[X�lv�ܕ�tlo�F&�� �5~�B����ߠq�l��S_����ʴl��j ���R���ʙ�iz��»*|�p����k��F����r�W
�ǉ�+�_� �?"Bz���r.���\W���R�����.�
:'�L��\������Ȕڻ��m~;��Ӓi�B�=nY�t��M��F#4�/����������/~�,�V�̢����B�� ŋ �\'�2�=�#�����.��B�l��s!�'.�����g��S�*�����2}�0�{~8�Fc�4ٮ�����Qp��l���]��meyd�ە�d��mt�};F��;�6&^�eNO��`�"]e����җƋś�H?�r.�8:�i�lq�K�Ӳw�C�߬�ne��#j?!o!���%�n����wwS�8ܪLzv�N����Z��w	w�2)���)ݝa���E%�-[����'ô�y1i��J��<]�#a���Z�眬DA�6���C?�O�� H��S����(���ǜ8'��P�%�[[܃�3�M�	I�IS�fڿ��p-'w�� �,���ꨀM17[~�o1�ۡ@���77��B�F��~�Ь{djFԶ�1���g����@j�S�Q����0o����(����:[��F��50�s^���&F;�O��IG�$�T�:�e��c�tdxjW�	���Κ~���m5E��}+�����p��T�U������_�9OL�b�𙥸��?<��\�����l��p_{&ݕ���s�m�i�ja&!a�����l�8z,��Rr�Ds��emڳ�'�b7�ۯ�ZMQ�?=�-/\��ꯀ�}��]��O����W\�R[��F��	��\�<�m�Qqt��R�uF��l��eN�њ��+ ,d5�Kn�r��}�ʗ�M]�K�y1Q�^o
�FH��}������-D�����3vӧ�)>�OTt�:�Tk�e��X��X�T�ğ��kn
�Oڀ`+���X{�\�s�}qR�Vk�</��8�T�H���z�jx�S$͐�L�^e��Ƞ�Y���zեj���R�������Ι�W(JY����w��ef�Zә�ޑWVt�3�;p\qڦ���,N�ɺ!`B#TgC
m��R��@=*z��&�US ���x&b�ʏx���ٲ�'���J�>���V�$�<�ڦj�|н���"�X��{̿'2�m��#��01��D[H|lr@�s��w����d^�4c�R6u?b�PB��=bʣ��!�ͬ$\����S�|{Z��*'�6�îD���Fu����J���7�qwy��"M,bbG	�n�Z��y��q�Әui��>�q�0���u�i���ؤ�Xb�Na����i�a��R����s�2R��ӡ���!
4��W��7ɞ��G��F��k1Ų�KWp�\�	G�s[ԊrST#q�y;�{)}9��p�u����F�\ܟ�$���!c�Y]�d��쭙��>��z}��B�O��%V;i́XjZi�=��&���Y�G؅{����D)�Ύ��`_\�����b�"l+�zp9�9v�S�QX���
`�Ф�X/�"��BA��%��:{]3�*���BR6�����%�TG��3��{��^����9�4��fav�r��+��nv%5�{_���I���N@� Ł�Dғ���H���<zsٷ�B0	2R�|��9ǃ80���ҋ�`�@)XŒ�$��5�;ީ���i��^��<�n�ݗ/~wÎ�4v�Kt�Ob�í:�.i=�\��׊��2T�>�~p��л*�'����w�/�>�ssK�5�1�5֭i�X�LQ���t��m}�N����ƣ��ʺW�M4�3�&��;]�-͏�}�W&i�b�{
��)teU�N�S�xY~엞wd�2�K�=S��b?�WZ����VC�ph��^|{\H�qv,S����oc����b����G]��|�p�e�� ���㐦7�����Tκ^|�G�T���^�R��ϴtժ8�k�
�JW��v ��&�>l_7y�H�4���5��-��Ĉw��~��La�gC/$O�p��!�`<5�"ĭ`�nd��47��A|�9.d��|����"�h?Pց��+��D)��в�0���em#%�V���q�']����T�������؟�F��V��3mڔ��Vd�lw#�\�6�b��,i*@2��s	�B���uy������b��X����d�|�wϋ���_�ߜB��s�G����*Iۖ3��A��L�٦���/�_)�9R�,S�>�n� 6+jw{��2��5�a�g��5�г��'�EImw2:���5/!�S�`��ɶr/���R��e��|Y���p�}[���N
 Ӌ�Jm[�����(�[4���\ �>�>1ݜ�D��xW:�p�[���C���D����:k�v���$�d9�9S@)���:��$�NKc��*9�,�vp&��U6MG~m#���fB�,�e��E����RM��)�Қ����U|H�Z����c�Qi�1<'��F'Q��@�}��t�%�\���T�j�!6u%	�:�̓�ˀT� �Y�����ƹY�f#Ḥ�*V|�O$c��JA3�����.��n��f�rs���՞�}�w���Ɍc>����&�5���IS���\X��uI���N�rp�+KAnզ�}��)Ź-ÍE�?���R3R�:Ε��{bW	9p�دO��Fik�eƫ1F
#t�&��%7�|(ׅ_��o�¢��"�P��Z��|�� |L��B8��޻�ڔ�����s0_������<�R�HҨ��C��rZ�OQ��$	\2�&�Ҡe��ceY��q��2��8���	Hm���������k�T"\�br:_�)QElxKЦ�J���������4v��Î����xn��4��s�GV�A�!�V�� {�k�Z�C �;�2f�
m�����c��A/�<�
��VQ%����N�:=��j&j�eQ�Dn�w�S>'��-s8�/�t	t<���__9�=�M%N�%P�%^6���FT�7ϾKV_(MSS4n�yN���e�����u�)�2i�(�0J��M�0��"r�{a����<&R�h�r�v?*�Q�V�6�,繳��f��`'�������'o�S4��j>a_y9>r��m)hNT*�x4U>׷�Oc�mD��^��;���E��}5�7��&Xx,��[��=�{�;�l��o'pt��YP�����!i�����ǡBP�{���2(߆{��MŃSJ� ��'��ݛ��܋ll��t}οg�-�nS�;����|c���z���|}�4�j�����OLJsIdY����~Hi��T(�����(�IIZ�o���0DuiЂ�گV�B�������͡�-�G���I1�8��K�]�1����P�vNk�\�DlX�c���m>�+9k�ql�:�I��������*���T�{�e9y2��T��d	ţ+]��0�^��XO\�pw��'6��D���'��5{�w�٥٦��%�����<��x�9[���k��k:�p��	����Dq7����`k_��B�p����Q�ɠ�o�A��A��_�J��`2I
�h�߭�L��������E>�X�<�?_�ӻݼ��I�מ'��a�U�|b����s�Yb�r�GH�ӄ�42�7�q����:����d��KǳR����ܧ��>�K|�}y��4oz+G�b���Ӆz�@1�;�[��,�JD}�Ip�ˠX������`3k�(Nz�fA	e���Kǅ�Q��xk�s���#�,v��R��d�9�E��ֆ�8��:����u�Д(D>�yt��#���(����ߜV��+��n͋��s���/Μ���9j���B��G��=MHo��Vk-6_R&L�m�GS��r%�K>'.���'�Ϭ�:�,"��<��8���0=/h����V�zZz��L�`��#�"�E���7)�	ɦs�N�.q��qC���������z�1fLs!d��X�:y��%��j&���C�$�0ܛ�W�ѿxX��)x`i��$.n6l�R��Q0�p�z���ب�|o�U�zy�RC��և�n GNW�{����:�E9|��e'��Y�N�ɫl�����TL.=��e�:0�:�べ%C<��x>Q��8M�>i����c%�qTN�MA�%g߮���p�����P;kɐ	7-����=�,�:�W�)��$"�BB��e�ߖ�����4-������g��l�J�ɾ����uP��|���D���,^�>����Vi�}`*�0T�j%���T�q�H���kOz��^J���S��2�Լi4J��\"04x'*^.>��w�+ �M��-�0\"��VDR�6]����[��-���Mc"����@u�|�{\VY3- &�	Ճ�#���P��G.u�c�bp�m�����IY�U�2�{���*�+�n��Fcަ��c6�	��,NZ�\��L�穥�3tM �k�1^����ib�'5��m��=Bx+gC��FQ몤ڪ�4[0�lo,�͑C�V�V�%F�ӡ��^M7�����~������kc� �Tԡԫ��,@��L�[x��8�i�͆�,mJ8�i�R��M��=A�;��wc�c	��v��k^�x#V���yK��D��_?O�'�s���C ������AMzC<��mȈ���rBd��R�nJ��r��/��]�ypg��z��90����Y�`'S�-����W��ݙ�����4PҘ�����/Ǹ�#����-��Q�POa�BBi���F�b;қ'mz�s�(��"Ӿ�Ũ�{�b���ƣ�h@���`��fLk1&�^��9�+����c�W}G��T+IAQ�f�v�ϧ��U���sJsB��GMia5�_� C��n��� ?}��]6�V������í�u�;�8U^;�I�����l��N�ؾM�748��n	j�ݢ�$qky?���s4���)@tӵ��W �X�"���K�g�Ƹ���ޖ[��Z��h���8�E��̀���ќ�(�m[q���w�ba�{�5ɻg���<����~��44��MSB
�	_?��з~W!�L[-�Z�&�M�����7n��ʹ�bđi ���h�S�>���!�_�[ϗ�&[�)���켊G�$�:�
Y��8[w4�ƈ�ɭ�t*G��������!Dۢ��e=.+K����Gtq$ȏi�{�l�ҵ�K[�?+{M����u���6g�X~�!��7�n])ӢU*gTJ���m��N8	y8x��}�`�t�Y ���;��Q�>:�Cezg�!͈�l~��|)Or	��>���~~���P�k{Ο�^͏_j!Z�)C�e�tܖ|�O�=�U���=�JjV�?g'_m���+q���Kf^_�s`%b7}N��],(�Q�c�I��*�!��l�n�S�Od�Ϟ(��N�+l�:�,��0Q�I��V������~e=��Ӵcw�>�}>�b͙ތ����_ą �~h�0Gig��#2���
�i����1�E$=�7�F�M�99%��7�;w�J{�b�=+3�Y�燪o�`Vd����[rw����������7A���ho
.d
O�0�x�s��֓ߞ�x����'�V��[�GH�_������	�|ȵ(�=L������Wk���ۼ��e��傪TWFt��r�B�(S��O��_g�u>�PStxk\�`�?f��?`�á��݃p{v$�ͼ$u���p�w>�=�s�$>�\���bύ���X�Z�
����4m�K[W�Fk+�mU_�FO2������3���5��DS2=�o�(�!(<�x���Eѿ���)��!�U��4�|����$e�>7+g��^g�>�p�-����f�:+LkZ�yU�T���ssW�O�s��?�Ձ&;۫E��ۆ|�Eqm�(N�c'��7�r(�4ě�+&d�	.�0ud I���f�
��tG.]l�oV��:В������?�2�%/R���j	C'O8���2��j�'���+�\�e�~����d�iB�ͣ#�³f��&�Rm ��4��w�ߞ���*uq+�Ǎ���5�V�h`�P�`$���Į���~8Sӌ֒�O��]��!��79O�aB�Ҋ��]a�Q"��h'�g�N��{��K˧�s�|<�پ���5�Xt�~�����;��S�/���4����l�ܠ*�R�]���#<dן���u��zj]�a��I�DOb�sj��+T�/�~�k':��=|N��,��=l�iuk)��$~�р��#\���Ѕ�P3�?Ap����\�7[��u�@��دN�mB,1�N����Nţ�� �]1�E�@|텅��;��Y��b3�����CYN����$	�����nUŲ��&7b��2H*�{�+�\Q�od�Td.�&|7h��Yl6�\ދ���[l|�U����O�Vk�`'�D�)���Z�Q�E���k^�����S��h��ՙ�J���m�$E��66�-�ȩH�v���O�W�)N�C�co�f[�{$�oI��o���|�$��:t��t���Owt�囊ȃG��I��)���y�����ۏ�U�tOCJ����f��]f�����j˗�1��X2|�c���W��a�&?Y9�2�}�Y��P�vp9W�S�SU���`�lm^����X�@m���!�3j�H�]\-Bh,�\:{�鵩*i�ZRMr���d�$\�',r�"X�n�w8�T��ԂN��@����Vȇك�S�����x]��z�\]KԴ��,����L2ėe	,�;x�m�u��wq� f�|9Ժh��;x�.�,s0�4B� @Oj��/)������?�2hCK�e� {�&���@�4�C�̔�	c�u�O*��g�EX��z���ҧ�6w�6+�ny6JӚ��!A�ؕ��FAc2�y1��7����CM�dRʳ�fp�L4-ϟL�r����
0f��,5�g%���e!\�����u����g��JO�:�'�t�=U��3[�Ff�Z��܄@�g��G���3����m��u�W �	�Q7ȑ�� ��` s�}?#�N�_�����}���sԏ/ߗj���əWO�J��}?�g��ţJC�?Iu���f�.�71ǓF��M��(_9)��S�ѯ�Az�Jo򻕇7��-�8���]��ZG9��\���V�^�.��[�F�N�ǀƹ�5j�z亟��A �\c5۩ӽ9�M?toi�V�$��*�4'�A:�������q�\�3Q�Ȁ���k���_��<@ÿߴƥ��	��M����-�s1C,hHQ�;˹l ���:�Lh�~���(j}-m���?§�Ե�]gQҭ�eO��We�?1�#'��I�_ x~���};��ִ{u6�u�ƌu����b��[\I#4��w�7d[Z�������Yٴ_��ͩ�pAs� �Ŏ�x7���}y�wS�Եe�� �-�*c��@r�V�Z!Q����r0Y�J���|;�4�R�M{;�������?5�����Xc�-6�6��Ǒ�����ZG�9�pē��}��N�k�K�z���Lp �Eb U�NF�u�G�;��+;k[t��x6����.>\wیc��~*|2�����@��P��q�]Y�A�G/�d(9�|����)|Ϸ���B;ݽ�V|������-����/�k~+�O�y�+�i�hMD�<�.[�X��и��+�����>��~$��F����M�7'E�>Ҩv���P+��ҵ�jV�������s ��V���R��L��P�NN%]� ���?~��ƿ�縏�֬�K!�� 6�!=2:������*��ֱ����Q����_��=��H|{����uyu{�V�Z[��H��Ȉ$���}��YwF@��	ӯ�|I�]�i��oiq<	}n���Ơ�x���@���[�x�t�@m������m��h͢Y�&�8��8*���s��m#Z��<5�k�ֽ��d�$���G'���v��**F���I�<����C�'�R�b*f�vj���˭� C�~6xw����-N$��#��w>P-�� /�_k�O�ud|���
�3��7�1�|��:�����N��O�\W�3���F��W��#J�R�)��o~^�fU��=)�ȾX�8�=j:��VՎ3vo�H-[��e�B��ܺD�d�Op��n�?��Q���x�=�����yu9kl� ����� �3�>&�{y��޸Pג/mǧ־��Z|8`2�(��?���f	�H{o9��zj�F�Uj���?|/�k�_­;P�Ű��uokR��m�"( ��>�}��T.[!%���K���l�I-�DI5in�"�������<p{s^���b���ş�CV���ӵ+(5�/T�6���Z$��n���p�v`r3�zƼ�~����4���PuK�u�� 9�X��V'�v�oF�����F���,�o������^��?�k��������7^���������*����X2����?��s�מx��ŏ���=����{��L5v�Q�[Oo�#���#�`��N=	Xy��W"1S�Y�i����~ߺ�ƍ,�f���xz�7��HC$����S���M��-�2[m��y��d�	V�w�;`���^��1>���C�$�IrR6�E��� ��s�〠�����F5[�@[[)�YrWvd�q�������rj�:6���cܻ�������*��� �sPI꣈�ņ�hb#0��6���#��׍��\[��:�	�|�Vs��Xle�8$gq�b��TV������q3�o�*��>Y�pT��tbIɇ̸�0�%�ǵ�Aff(=®�8#4�6GeZ�fyJ��̐/˕.��:���I� f_G�FIa��:ym�����
X���������4�Z[\���K5�D�N�S�s�~�W�3Y�l���<P�Rs!VS���c����?b�����O2���(��Ӝ�$�=rOLf��g���\�W�~h�{���C���=\��5{=GN�xb�����Gz�jZ<����;�`x\����K�>4�M�ԯ|I�������^�WeBd���ԓ��k�9<}�S�����پ���4�����Y�����V��(J�� 1�^������ŋMo�f�p�e��q^G����e��b�i�2>R0H�8����:(Q��*s���x��"����w6�ٗ0����Y䉇YL���g�cxG�:��,f�&pJEkg���@'
�����溿|b�g�-wT�'�e��ئ���b��Wj���=��G���><�3�O�:��Z�=��!Iգp7#+u��@ ���|�-O_��zG�����$�t˝J�H�*-�6ec����aU�(�<������ gM?����U���L��������*C�h�b|��A�~���>,��a�|L���wS�u�O���:�
�0���u����~�ZW��MJ�L�f�w�'����� ��;�n	\�,�[�k���<��jӛ�*��N�?x�~���|����m�[����y���]�B�;H�ƀG���66��>�c�\���5Uմ��>�}L�"��6��ߎ���{�ǆ���jZ�^�O����P�<D�|��;���
��hf�s�Myơ��<]��o|����M:�O��͝�9�io �+a�\�u��͏�s��U��O���z��.hZ����9.n�������I����$��5�iky��nH�2#"n���{�k��#��)�
2Ÿ��cpc�����mu[�Pn��&�Y���brO>�ֻ%�c�
v�r܊;��/�70ﲙ.��ݲ	�E%��8�`� ���4���� ĺ����J�R�c�ޮ�k�j�X��R$ϗ����6��W�V�ib� ��Ku[�dR]��?*�������[�����:v���'���j���Z�H�d���÷�#Y&;B��Ű�����1�;,<�~V��+�i�� ���b��k'��A���mus=�pIRD%�
�Vf�ͻ;�n@v� ���MWúN�iuogu'��3i4�"�c�7���d��au�p�ֶu�Ɨ�o��^jV���j6��q-�4pHI��DbT����z�/X�V}�;���KO�,l--c2Kupn�� ~���w�c�X7%;�~{^�jx�T�_2����G��/��U�-�t�	�5/6g�G�����CD�St�̬P�T�p �(nR���"�@�����ݚխ�6��:}��5)��R��v���>�R��v#��R����k-��,I��M�y�����?b�֗eiib�7����XG�i�#+)�npX�p�b0Md�=��������rzi�n�O���Aw��qkes{��x���q��2V���dȍ)i O�������^�|�����u�ܨ�8��FL�8\�G�[�U_�� ���7�.�8K�}�B���.����.��H�` �-t^���moP���W��]�ە�m��6��};�vu�k��e�B�*b����W;�CT�"��N�'��7�˷��q�G8E$Î��ҸO� ��c����,���c�����|�I������P�Ǉb��&�`Y�p�#�qEw) ��0#��ח~��t� �n�4;;���Koi�h��F`��#���<RK{F���=�5Y�� do��x����n��gIt�/5�@T���*.���v��q�_���T���M4�,�d���ԟMYC�[�M���l`mA����L��4�/��n&�+>��9���2�1qʫ�,G��oh�����m���y��6ZlV�]���6�r�Y�.��3�s���h���>Y�-�x�W�����m�8�C��~'Ӵ�&�M!��k�Y���q��ڴk�(Kq�O���© }�o����<���&�0�G8®H!@�\c �����k�7þ(�nn/5m_2��,bK9	����I�V`Њ���X���/�2��Q�_������Ba`|�� xpT������j��=���:TZ����뽏�����H���5]�i�����9��-����>�]��m4�>vxس��p��#�!�oB� n�+��#|v�e�J�ռ3�h�Ǥ[�����Ǩ�,����䱑~u
AWɚl>*񟊬<q�-��;���F�!�k]� �  Ŭd�i$��*M%�άf/괥(��z5��MWƞ$�mc��:7�om���I&��\��ۢ�1��_5���\r�̷�iu��>��xf�4�+}[I6C���$�q�@zv/�G��Լ%rR�;���j	򩉯$u��`+<u�t5����5K]/��<h�����乸V*㏼��ҹ=���>*��89�q�����]�g⦍�t�����V6��n����E�[j��v	��cF�ڄ�n�|��k�|f}�F�l�ח+�Ģ�*�- ���q ������qyu�\j	5�قiPMp��p�LJ�6R�{.T7�)�S�� h��tk�;K����5���r���k��Tp	�\�U�x��剨�N7P�]�e�������<i�ϭ��ʗ6�rZ�k���ǅ�#�	5��M�Y߾ nq�<W�?><|E�'�1�x7E������ƒ&Ӣ�Y�e۞N�r�W����א��s�3\�����5Js�a)5�����8�j²����%�^%��n=>��s�a����;�-5V:��i��������A$���f�����OB�P�i�V�C"�kn20{�V��f��Y�,�l.Y���_2�<{gqC�MT��%���$����zt�[�����[�_���d�||�ܱ�y��Ǚ�iJ��k�=����#}�=y�8�{=F����y�� ��{�{�^��4�});gZ�����5/�n�� ����jְ	���CL��s���u�}p�26�ke*z����������s�*���.;\��e�C5�ݴ��IJ�/��$p�Xp�����w⫋_�����͢"lKW��|��78��{V/���/��^�o��x��:̆=+B�,PG*l���I5�x�G���7���2x7�{��B���CB֋���O1��������:��qz���8;/���;E��-��m$h��Ww2n�&�<٤?x�8Ut
ׅwL���#��AZ�b����Rx_ƚ+mԴ)ܱQ�c$d��<�#9�5���.z���ٞuXNq�����so�D,���ُ����kM���+������S�����e-�����O`�[nY�2��K��?���_�����C���e��y�bo3j��$�rR6(#!Nr $�I$S��pq��;� �>�ddI"YA<n��b���\��bs�[��'�����<�k�f  a+.�8��	i8ݏA[�+��[�����j��	a�gI'i���Z6�o�G#[�qq4p7�r6����\� 0Y���s�?�Ӽ����t"��!�9��;R�į�/)2F��T�
H2��\�eg��`f@ɺ����D��g�Z�n�Ĩ��Ҥ68 �J����;Z��i�Kx�u�4LJ��7S�pXu�y��n�Ye�>�̏ �ǅX�z��7z矫� b�9ol෷�)[�U�r̹�y�$������a_�l�3V�N*���G��v�E��m��ς�J[q6�pxa�홚�yc9M�W�A�z|��;�����&��.��y6w����Y��q���Af��y#'�����O�:/�����~+�Ɔ�����2�O��Y�vwTV���F	�������|\��n���xQ]6+t� !�h��&l����/.+�+���Kݛ��i��%|��O�u
��Ww�y_2�N�Ia�2�R���S�;�?�� g���m'F�io��40��;C`��X�y 	' ��<?�G��I��hՋF<�V
y��{
��j�P�K�N��b~9���"�����t�Ϩ>�/E�Y�M�Y� l��d?g�_BZ90ـd$�a�毦<'��3�6��A�c�M'�x�}�x5ݖG!R6!	a��A���'�v��}௉��l�<k���!�ѥ�b7ف����b�rO�	�_S��W�5������?Þ��9�x^k����K�2����U6�:�0峻�xհT'RU%&�9�xCK���M#L�O�4;@4�8iRٵ��ZT}�l�v��-����`W�����C��Y	j�ڍ�rKg�I��v(�D�de`Hʖ�c>���J� \�~���xK_�����^�}��y�m,���NT���`�ּ�Z�1�]~�ć�G��QҼ��.��3ۆBbfs�p�O' ��)Ú�m3���{NJ�'���^��[�-��5�M�-�kh%���k�6�tۜ��$�l�r�1�����Q���-�q�������xcX��<7�Awpeދ�I3���ԎI�~����K[�.GHs6T�20������ֽ~^���)��_�?,��e����=�[ �%�nWn�|����� ~�k���>ԭ�2�����cWps2qq�p=Go�76#������)!r�'�A�A��⾬�~�U�|I��������.�7��b9�Dj�Sa��1c����q��EΓw�=���T����� ��hV>���|=���P��Л�nb���ɶ<
"b���
w�G�t����U�͹hf���K�$L.W��[�溿xS��-��j�6���6���A��d%b�M%w!�seRJ�k��u�J�O�����RӮ4]O�2چ�.4��!�R�(���8�����*>AC��ro�vjx��S���m;O��ңhl��}&q��\��]�I�r<�,�f��5��� ����r���U47�Pԥ�6*�/N䁜Πo*N*����sxU��/���w���H���m&� �Vc̒����P+��Y�p���z������O��Ʀ!~��� �d�Y��#���+��ɰ�R�}�ӡk����u�7�o\�T�c=���������5y �|,�H�q�*A�Ŏ@#}yc�����+�񷋴_�����p�V6��,�98H�A���v�X�N��ڲg��MY���7���~&x��q�꺀���DQ�K46D�yF�r�pV�;�i�����x��++��q�L�f�o����d˵B�ecÁ��W̾,�U����z��P��=B�`>B�|3D8�I?��	�.c���;��e#qO8^��_AU��MԵ�����k����[��:�Ko]�zu�2[B��i�gF�<cv���&�/�:=�ǌ��:��}J*��MU�2�I���F�����q�$����֯�kR�� jx�ZԞ�no�)�0d`�.�i ����x�_�f����Z��ܪ��&�I��	' �3Wʺ��u\���-�/�7�r����T���i<��7�&2~�%�H��F	S�?�W��_�ߴW�|M��1j��u[��,o$���etkG�rC���� S^S�����?�rX��l�/�g�P��У�P�~���k?ğ�����ޚ�f�ue���M��hoZ9�1iK�(�W\m�S�z�:�+ilxxL���rIٻ����������7�	?����KB��O�/X�i�0!X;(PB�2��ס�>	��n��js��[i����nK�|��V��R��)!���c��v�vx�㇎|y��������PeTi"QnP "
� ���~����K�>��x�;I�X��3�˲�v%�ಁ�1��&�^�,�VS�������^��R�o�-.�嵦����i|l��]/VHo^�9��HbU�� ��W]�Qx�� ⮝?���.�*�R�����D#8öK� !y<~v��act�pj�]�^ǩy�m�\���F%r�\p � q^���Կ|q�k�׾"��]o0�5�v1B�Ynr�' v��}�r��:X)¦�Ϣ���������K�4�.�C��V��x����O!��vܾY�B�FN6�+|�'���2�I𵏇e6qٵ�����N��6��nF��B�D���� 6�� ˩jG~|17��M�R��tI	�Y��%ڻ#V����yo���/]�o�[MZ�Ŷz�����c%�:��}��ݖɊ��c,Wv0� B��S����S_R���w�W�����`1�іw�
H�6��0�h����_kޮ�5E'�z}~�|�Ti73|^����y�����0����`uG�}�t�:����9�ǭy{�|�isB���$��/N��}�CqVR�x*�+sfc�+UfG�ݐ=Ȧr��w�x~�MsN�������;�Ǆ�r���9�eԣ#V�������?�V&KyN܌� ���=N��"�p�D�D��7�4�h������9���ec�� �~��Kx���Fݾ$ӎs�N3_|]�>�!1��{�鄹���u�Ǚ�s���> ��>1kwv�_x��oge�Z�glVK
��t���XF{����f� ��W�@�Y[�F�j�җ�0�T2ci�'� b�|����x��#|?G��n�WM��8n��6���m.Wm�k��$nq����M�J��x{ƺw�Hu�m�[KD���g���&&u$�w���f��=H8�g�birrl� ��������G��v�D^"��I�B�w��x�d38{.Ӝ�@+�"� X��_�yx�X�d_�%�j�vo�hK�ɦ��+�p����h]�hg$�<z��x���WysM�x8���f�|�y�B�������G�֞�鑤�9W�����q �[=� ��b� ��k�Nʟ��i�"����r>VA�d���dQ^��1>���C�����d6߆�H�n�K1�prW:���Kh��X�i�+�	l����w�� $��\[޴pA-��&+$;^6�"|�9#�%OR��~M�}���rH@_�gwmV8 ���A�x�n�@�w�9�k�ؙn�!#p �;�
�<) n ��/�4�Em�	,MT��7���wM���O�F��X��&�a�H$��#s1 g�V�	�5kegђ��Q�l���P�~��N'�����݇�|�v���yc�s.ܡ|�}M}I��1�A([o2�P��H[g�Q��0�v��dy�9��n���u��®]��IT�=Ĝ������c�D~Ӯ���54,_x����Ԝ㰮|C���g�<�տ3�
�x�V�����Z�Z��7:v�koy=�j/Y�Ɍ,Q�����T�3���ߴ��{�߉^мy�I�iVv�w2��I�H�|�1f'�URG�9^k����,�v��mSA��焧����-"���M#e;3���
:|o�v���W���s��G([�+�Ko�J!R�b͌w=��Ƥ%>W������|��E���U�.uG�*�mn5=�rʸ� �p$�n�C�t?5?i6?����Vf�����l�!��
[ �����]R��n!��rʷ6��\�u�wZ����L6�p�K�r@8�o\v�]��Z�έs�� �V�i� F���յ�6�[�t���4M<���\(*��,�+�Z��J�~%��ph���/.�	����'�X����co/�R�{rH�W�� t˪A��'�O����5��v@X����0�{W�E��;��:��P��Ӯ�+��C!RHW�JF�~���H�Vl��Ne�P���v�]�t�����Z�� ������{�&�g]+YU�cu8S"DM�����&��׿�Ěg�&�Oá6��ɩM�	��>&o$�����U���I�xw�+����ZF��9�#��f�T���$�y]�y�Ċ�b��V�,�<.�����Z]���j-sT2���?��k��Eo0F��*ۉ;r��~���nxqTj�U��n�O�����G٧�[-�SVxL��r��r�q�}�t�l0��[�+�se���rwg���#�Ce�5���FC$���m�y^8�?Ni��*�5�nIT~~�~��⤵>�q���ZM��4q�����fW/�����}�� ���qx����*�+�sr'T�1��j�*H�RO���_�z1Ԭ��L]JY�cH�I�S���9c��{WѾ4����5a� x�b�	x��&�t��*��bE*9$x�
n#r�Ē�V<�u�J*Tܽ:}Ǽ�D���Ph��_x[Jю�go�H��ɸ;�Ԥ�UY��FN23� /�~��4h� x��|a���qp�%���Yy8�����-�>���V�%��<5.�w�����K}.�d�Q�f�%w��iH�.�*�6��?�[��!s���Oܯ�l�l����W��Z��\�1��T�����\�b�NsJр��=�Ed���w��3�뺳}�M��{�� /�s�9'�z��}vȇ�3�<���oY��z}��|��NYݎ�bq���׏<m��G�zַ�1[�������
~S#�$=��������@�����ş�GF�m>ݮnt�/Q�����W�$�"�����Z8�����^��]wN���>�iq,�wӃ�CB~�3)u1���ֲ�'/ul|&q��^2�E��%���7��H���x�����s�*��1��kd��:�A�#�5p�P
���� ��]�c�)�Ц���?7@�}*y����� Kc���2X�Vmtm\D�/�������?J�o.L�1f!�l'��3c�O�W�e�~7h>+�uMcPӥ����b�l��s�Is��ӊ����ƕ�g�����5��^����\���}g� ����@:���W<�����+�࢓�N\���l-B�� N��5��c���2H�s��#8=���<-������&�b�ie�a��IՉm�vHlP	�1����iq|��
������Wk�nq�W@L���ۃ|���?1\3A1*�јq��^y����G�-,�-��`2𞟗�Q6�Y��R���k�>��5�Z�1Ҭ������npp\�<d(���x��-S�� �?[���j�f�t�d:���kIdcyE؅#1�	@=��d�]ۅ����v���>��w5�o�@�U��z���������
�jNWK�ߑ[����;X�Ѫ���Bw�ky�}�Cx�������i�?�f,��+�@#��}q�Nƒ��v�$�am
m%�B�q�R� �/h��,����_�T����'���.߻�L�?h� ��!E�~��[j\@�� y�랼TR~�����������!��f\T����k���J�P2�ls�� �W�ðy��8�яb?Z�:k���V�5���r������*�(�3�e{`�q�e�2o�_o!+7��0qi.-7�;�^��h��F�¿�(��t�xN��֑��w�h�Eh�\�=�W�d�8��^�k��-���Sľ��޵{>�<��wjւ9m����df,�ϸ�6>�F2���K� �Keq����s��Uh���!�t����2�*(P�my�;ONU����?e�[�����f�BB��וu�>_�^�<='�>�	��V�
�6��Ň���Nk��-gH�Y�Ub}"_p1�����?�x��� $��g�7}/�e�R �8�dz�����}=e�t,�FdWR�@��7˜�yb�`+H+۴�ܨkq
F�Es8
�p|�F�����֟T������)����v|M�$����("��&�Ō��p:�	�@��I��<Tۮu/���v�n���I6���3�g8�@䓊��&����K���A[no��u���ۑW�[���.��o4�F��H�e
v�q�P�8��Y�mZ��ȇ��n���zo������Ǭ�SA�Kin�p#�<�X�Hʒ6r<�ʏ���Ey��>q�P�'�/1̍aϘ�j� }ҽy#r�!���(EE#ք}�Tc�DrZ��k�6iAV��k�IoR0����9� �Omp���� ԕ��YH�|�2�fu��y��_c�ˊH�D��xެ �8��*�Ьd�_��L��p ez.U98���,j�u�5�Z^N���g���F7g�Ȫ�)�U�`W߅A�u�� #&�H#w��$
��i�Me=�K��tl,s �*r[�:u"���7�VW�V,��F�r7�,�U۵s����R3>��gY�R�-�~�0�����X����}[����H�]'���37W��{@�����/��ŭ�R�g�"E���7ʒW g ���>���� �<?a)VMڞ��$����O'',Fs�W>!^�G��4�/����>Z��	�f<�Ө>��>� 犥�ᾛ�-luH���H&U��7\{���^�����w��pn� f$mr��y"B~��'铌�x&�^�&���E���M
D��y�ؔ��	� ���x�Ź6�� �wR/[��<�>�V(�|7�yHA!���>f�Ζ?������ ����V�C1��A��{��^O:�/�Y����"Ϲ&��aXs��{כ��ĺ����-%Ѭ{�a� ty�;"bc]w�����E����Kݻ����|%�ci��òi6w�l�O���~0����נl `6=3Ȯ
��7�����2��c?��Ҧ� ����� ���S� M������&pT�Z�瓻~k���+xE<M��������y����`�G��� �q���FMxd_�����Uk�I.�w��V_$�(���^2����8�Wz����k�=�[���=��NT��$U�F �Pw|��9�p��<?o�X�6� >�[j�^\j��C|��L�qi�y%�vH�O�c
���>���^*�i_Oy[��o�uۯi��\��#�2O�=O\d�ζ���4�}��m,�w�z˟j�ɭ��H���a��x��2Qf
�	 l9�kn�X�����33n�\���s��A��^���~�r�~%���%����e�|�c��c#�ӌc���T��xX{�ό� �Y�K�uie��g����tUbd8Rx?/���w�Mc�+X���W\�>l�<��5�N����x�N�U�����-/˽�kH��I�#R�ٖL����_9q��i(�I>c
�=�v[���EA��ՎI�E�k�:~�ck������ +�9f.#hp}�����{�#-� �C���BW����M��%���m��U��{+�
�+y�,6�����Wq
����ſ��}��6e�8ǒ��֗V�͕�ƽX�������H�bى��y��߁�9�H� �s���zפ616޹Q���+T����ld�D��J�Xm�p$�P�b�NX��023���������<E�u__b{����%��+y�B���+4`sL\4�0���	�^�n��;�����ד�m�V�Ƒ�)�H�H�.�`�^��L���c�K��c�;�'�Vm��`��ig���8���5K��AAiww1;;��8�Us��$W7S�=h��c�3Q��P��$��s$�9[������~����"��?� =�zW�� �����/�^2�� �'MZXi�ٵ�g2I"f+�x��gwBدV��|��ᙃj^G ���e�O7ϊ����;QU�����q�Euj-���P9gؐ;g�(��H�~��}:����#�#��گ�������?}��f�h� � dk�Bc��wxY�a:� z�8 ��T���3�	_��¹��;+�R��xH��D?�Ǉ
N	�\���Q=Z���������V�ce �m���Ha�������׃�ѭ5�rkk+��>e���hc��8���U�Wb�@��q|�g�-�� ��^�w��Op.����sqH�$�f@u_@A;A�^�.\��K8�W��O�;m���ݴ�}-�%Ÿ�H�����B�j�$��G?\�1�-'�� ��{W��n��Bs�yT�� �/<#`e��ı���Ǻ�?7`�yf��˩����߳� ?,`iU.�FH��c%���k�� ��>u�렁�ib�_4�~�~����u?�_�kw�<77w��a���P�=I''�qYT��v<|�|�
�}��܄���i�sK�.W��7�T	���[-�G� '*3�4ֱ��������� �ڠ��r��FO9�0+͏���Ũb#F���vﱷk�8��r��R���#^�eyg3�t8lm�ayR��8m��7�,7q�6��@-�۳y�p@+�t�g$���K����C��v�@���*���9'��X�h*��O������4v�ڴ:�e-́��t���#oH�rB�b�����֝{*x}6��l'�#�Io�MMtX�Ӗ�]2�R�9ZY�v��!m�%r��Dq��c�zU��?�62�/͊���i���fP��ٸ����Y�~��ٴ�8����6��#d�>��Mz{Z�430�2���*H?��E�t�9g�C�s*^���]SC�4[�F���r�d���� iL��9P�X�������[k2�e��/�z�ZM܅�,>XDm����̤�cЊӹ��mq��&� ����ݑ:���6Ua��ڸ����^��[]�^tm#
��̥YH�e �LU�ԓq5X��'�R����|��xi����->#���e�*v��&s�R�O�M|�W햳6�Y�|������y��3�@���kE����;���ռ���`�H�ø��=+��v[i[O&�{y%����� ʈ��0��C�	�r{�pV?K�*{L9�k��Ͷ���,����|M�a���r01�OL� �Zv �ڗ�.�eY!/�_1N��K/��#r�9�Z-f�0"��$ݶm��
(9l#�?)`f�]ۤR��х�d��H�D�7,o���'#�ꧯ]OL����5��[ʠ���IY�t$d�����5[{x���i.��3���4�4����VIWfIܠ�K%��q�lm.�Mj�6���dϗ�@TdBFw&z�O�i�G;�
Y|�=�\��7iТ��0���m�$n���ZƟd�d�'Utu��I#���W(Ĝ�l�\���]�Y	U�+���,��I�dR�" �p��d�1�xb@�PC,n�y�y�Ԋ;�7 a2x*~RC��]��]Giw�C�,��y��0�<��brrE[�����Xv	���p��rwT��r��)mc�\����0���)$#�W^	�2��m�$���F3$�'�;U�|��1����P5���";Z�*e�]�h ��;G̹!���?vԉ?��u�˴�D���?�Ur6�*J� *	m`�,��0��kv��@�uW�⫕*N9�!r���14���1RUG�X�Ta�d1'�k�آI&��5�6�ub�'�l�C���־?���-��Da�)���ኄ�f��A�__~��� ��2F���j6�kH�������� �y�/���7�x~4-f��K�$)��d���I��q�Z���?�4�.u���e�X/l���%p�]��;�0	��|���K;�K�s\�����lz~�=�?h�k����ݸB22X��?e�x/����{��[��ho5�[K!`�fC˲�y?�p�����r��u�k�F�U��M�j����O��Eh-"ڌw�Ň-+�:��Tn2 %pX��~4�!����ވ�hZ{[}���|z1�k�{;x|�*���a �q�z�֮�mm:0��5�y�i��=j�� � �*dө%)TW� ��t��Ğ ��\�ǗZ��ωkg%��>��_ʳ��1�?.ౖ\��E|�p<�D1������W����,��ox������t��8_N�y�w7��7#����$�hQ��s9d��$��v�K}����<�Nݬ���E ϕq�Y��#�g��\V��=���.#��(�d>f�i
g�91d�ǵvڇ�O��%��w��>�D�C6���Y�0�0��� .�觓��Oj^)��ۭN�[ۙ�gv�Fr:��:W+��HSk�v<�e8�WRnv�� #�d��~���Pj^,�4�DI����#o>`��a�v�
� f�����w)���4�����52���#P�B��P0��9�z������-���_h�D��9��Z�>���VB����O5�B���=r�I�J����Ǹ�� e(�+}6���\�'�^��4��z\Ă�%g�� ���e|d��?����	k6������-��&�J��@w1� �0�����(ɼ���@�M�� Y�
#\�:ȸ!�c=:V��b��eZ4�=��RxWR�/�_U�K���ˬ�]ޫ&9�3�>2[�`����H��Oh�1�i�����~��v����9�@��ϖ~BIn���_x�/��j6���yʬ�m�IS��<��~�� ��_	ͣˤؽ��-�m�@��8ܭ�������*��Z�?��ep��޻���|mw�4zf�`�_� ��Q����.,�Y^EE��Ɖ)��$Gp2+���4}2��/�5i�-nu[�[��F��g��� yCm 0@Ͽ]�u�=+��j� �~����^� ���Dg8��wa`rjݷ�������x�W��Z��5�:��R�{������� �r**�I&���Ʃ�Ri�#+�Y:Ʃ����Nx��m�?�/��J|F����;�2W[��:�c�j_-GX�w6���'.�nI��s��'�5$w	�^��^h�5�Ӆ��t������|)İMl26AF�+$~W*r�M��τ<+�|J�P��?wq���{j�}� ��$dq V���+!�7�0v�������L����=�0	#��Λ	e,���m6+���{����k�� g���^񗊯<}���W������ �Y��$K&������k�c���6j-�����9� ��A��:�0n�����iR��im��>6�����ȇI�D6A|pK6����3Ҙ��x��� ���0O~s	�M}�ďپ�\.��ԉ���y�U�_�v��%���a擳͍���烎���o����������� ɿ�#��/�q\iy�<;�6��t�^����V8�v��9�s�>�DzR��Z��g������+%�&��s4o+<*c�d���׮ipx�RmR� L�k�K�*�U����I��[Im��v��o9r��0�}������2վ�x?�~!�W��]:���'�R+h��#6��k�}���0I#������zXlt1��A����{w՞uu��-�S�<�$�wbMd}w\d��|ּ?|9�/�,�x͆K�̨[�?h\�+�?kO��q���Is�4�l��9��jg���H�� ��������s�֖]��o)o�_��>3��kl�I&����:=�K}�/�;#. `�s�;�pA�м-c��&����W�
�q�܋ۿ1������ ����d�����'���y��d�?�]yg�~?x�Ϗ.��kq�z%���͌ilb1�@� 2�f �q�(8�D�Qm3��0R��QU������v��,d�tox��WR`<�u�)"�6)��9>�n���׊#¬Z�Ƚ��&=�^��� �u(�~S����n��� �q�t����i��ޭ_�_H��6���.���}���{��t��\yJʘ�6�`�԰��Б��]⥍����PZ�j�x�N���qbEiR	#��2�p�7l#w5�xN��K���O�{kp���W(|��T�������oh�&�n��� iإݭ�-)����;I�a�E�#5�i$ϣ�R�XB�eʷ[�+��y���ot����W)v�J���p%ӯ��0wX�s`3�+�}-��֡:�$wFxY�,"����9 ��(�ޗ��w�~!�Y�-����%�j0��!�8Ȟ�jY�"PW?1lf���Y�|�5��T������d��(�U9���y�V*�����O]9�ũk�]WɘSx����#�0��<��n��iQQ�Go�\�۹�{W�R��.�v��m�*G��P��$��j�u��1�'ң`�G<�<�l�[d�6�����>n9pp�����M�����kqm���їqb��H�QZr��3LEl�j�VWv�o���O��n-=[����T���P�m&�����@:U�x!@�k�[;1LE���'�UdL>�B��~�:��`�1����nG�����U�"Ե�DA�A����p��r1_%��������;6�&�E�r6!ʌy��p�w|������R�O�2W� 	�}	�⵳�9%�����Ÿ�Q�`���F8ٕ`�T�{T-kl�$���D̢�Y�r�c"��a�SZh٭��W�S"���T8'k)#qÐrs�"��/����"�����e����d=v��)�p��ZK|�Mߙ��K���A��@�r���[#�g�Xu$�I�!�ef���ZH�`�e �̻�@?4�����k��;)!�M�Eٌ�$�"���� c��9"��ᣒ/��h��U��IcٹZEq��H���d�9�)�_R].���5���'�)�i�iP��0�N0(�Z}�62I�Յ����v�e��U�3�rq��AW3�[(�!����W�(Q#o���RBg=�	=�C��%��^<2�?-��fE�یd}� �OH���6d�#o�� ͜ S8n2�g r@&T]�)���S��C#ۻ`���S�8F� z���F��_�<�>_���8����<� ���
�-�RѸX�h(Ѱ���*��)�����r%լ~i����ی2�RX��_�Cll�`W85JE������.�7,���ό1�nS��^Ƥ���p�+H���)��drUY��\�9��v����.�t�*Xx�5Hȋq_���O�|�~����7����k4��c�%�w�������V�� ^���j�Z�%T�i �q�+��6x9���O�揣�e��_�v1����l98`Z�=�8�{��I�Ī̬�"�-�)ی���ۚ�Oق[�G��Yb�(h׫~�R ��=G�{G�� �u+�2���Kg:�PB��0df9�ך�}�����?;dW���'%B���֜�meg������ e���ZHY��UU�^�Zz��6@���~�Oj���Zw�`�a�f����	�@�V<�#5�_
���U�i�F����t�:i>���*R"f �#}�<z������I$�<HX&q�g������j�W�?�g�W�F�.��-���ř��q0�v�i,r	���iY�
�t���t?t{ɼ#5�亶�+2A�Ak�<!i3�p2q���o��?ۉ#`���d�������v�w�����4G��L��感���drT��O�x�F������^�T��+ہ�5�srW�����O:U�%�p~�uh$h,%ei���qR�k�3��!�/��O�s�ƛy�c��3[6��x��?<+b�|�Ap�+�S��D��1�e�7E�4nF~b��KWh E�JN��W�|�I�|PԟG�-D��4���b�I8,�Q�:�ھ��� fm�@��е�+ķ�2���6\��,��� '�8�
ٖS�T����v�o�t��kC���s�-��U���P��)��n�A�}��/���>��2//��7rW�=;
��3�N�w׍�h"Ԓ�醙m(܈���B�%��z`���~��K�5/훩u�愫��5PJ�#�	��U�֗}��K�{��^���&|��ma�_է�H���ң]��8/ ���׼6�o��N�����i�6���TZC$�� ��:�G�w�/b�͚ɍͷ�-��!����n�uh�7|�|��hEo>6Gy"\\�>
�E��(RgEY6�P08����b3\F>1�Y8v^[�n�ml>B\�׹����Zߋ>�"�W�м��ҥ�έ۾Ʊ���B�)��@�?O��n�1=����o-�C#ζ�G4�� <�&y� ��5�=O�I}�I����c�Eu5��V�n&U�R���g�<|�"�?�p@l<�÷^��k�m��Ve�+�R�)a�pȭ�dGr��l���B�����k���T�F3�yi�W�� �|����k-��^��EW2o�0�9�q����V���'�9�I��m65u܂YB� |�k�º�x�p�R�U�� ��^����?A��a�*�^��O�hį. v�=�t#�lb��-O�����d�[�	Np���8�Ga�^�Z�-�� ���w�5sS��	k��Z���^]\^Ccy���;����F�N���a�=� ��\����|��`�5c���i�^��"q�(��@� �Y��� 
��S�� kD���	7_q���*��<�W�>2<sqq�?��K]�d��7��NZh�c�2-H���N����y��"�8V6-ѻd
���ȍ1�Z�>��|B�Q��/<�	����^|�nm���o�~c�1հ�.�8Г����pc�5O����9Aݗoʟ���y���2�������T�K� ˃��y��S��[عou<
���2�#(n;�y�i�j�=��Rl�|������~S��5����]U�h��v�'�ٯ$��1�j<��%�3��{�ϭh��]ׇ�:�K���_Vqז6���ͽ�Kweu�s�"Da�R}��מ�Vg�.�$�d��.��G�}2I�g�b�'��&���-]Ǌ�I���]"md�k�9,���+���'�^��i1��w�P2�#i�IclA?������b�MΊ�ҳ�����1!��|� 1��}~��|y#7���X�,xIۙ@zs�ֺ-�\dְ<{�|���������}h��1��Z��q���!���E�L���r $YY� �3#������$����-Vy&ӯ��nc�b�d�����6�,�db�����߷x?��Lm�k�$wSrC��Є�%Q�r�8!}k��b���Jm���nא��w1�hn74M��c��5���?v�?�]G�$�E��Dѭ���!`��2�,Dd1��`w  ���G�\�|��K�w H�<k��PN2���-��v!�%�-�嫑 I�6r��mpN�˜�ƽ�uKw�z��%���@@͒Ő��,�O%FA�XZ�{���h��Ӣ�D�F�cf4��#D�~`w!Hl�p�5n�m�Ŵ����{؜�3�@�|��w�j0���(��#35����	 c<�C��A�{���"�enL-����� �&F��nv��s��P���cU�l���{[8��R9��g9f�c�F�a�iێ��-�����i�)���+fb����%	��Ԝ|�$�(�����^v�ٻ#*��p��v��Nj;�%�24�\�,�3��y\}�A�>U$l���55ŵϘ�I<m+|�O�d<cJ�N��R28c�~u��Z+�i����� ��|��ۗ�I�!܅cVp,n��vl���6IT)%��v��r:���fb�lר���%�*�+�*m���1͉6�LRۘnYX�iTr��`w�n����PY ����{f1 2
<n;xی�y�
�j�¾L7I
;�{v�z`�A�� W�߱�Ⱦ	Й� ���)\������Г��|{wn����B0��l�c�x7pI vvI���f��k�F��H0��%��~�sb?�#��X
������ �����4���4�N�w�Oh�ͽ�� o��1Uv���p��Q^��j|`�^��� L�<a��V��^��U��R�h�Q�#�z�� ��n��8%����ˈ�."Yn!Wp���y�q����	�w��"լ!���"����:\1�Io=[$'~3�\�&��xya��������)�kY��0�#j�*�����+j�� ��I��� HV�����<�z�쫢Y��U���6�}�g�*O��0�W��죦1-���j
�iR3q�x��O���{� ��M5ܭ�oxeh�1���>���v�t?x�ƞ&>8��;}Ɇ=X+G|^L4|��#�F��Eq7_������[�\��m����G��q�ں��-�	�\ߧۯH�$�GR	,@ `��M֦��Us�'�ww9�'�&���c�}Ua���n���|Q�=��	l�B��H�m d�ï'�?��Zl�va$ǰ�H?�kܾ#xwJ����ȴx�w�>�-����J�Cc�0k�Fa��F���\T�
��J�]���Q�a�*1�=��^���ḵw���wT;w�Ư�L��c4� f*q�>Ձ�\��~��o7LO:��r~�A�澚?9�[���o٣X���:-�܋[[?�y�I�j1l�c�Y�ܤ� �k��&�M+I�N�4}7X���_$^�Y:�f�r��)`OB	����-K�n_O�k>#ʸ+,g����mӾ,k_�wY}�I��Dr�>�agP�`����_)��kO*гM�_���c�
*�>��+�g�6�%��ZX��>^�]���ȏ)s�
C3��t_�:}��m}�i���76�W C.~���Or�k�S��M>�˜��S�s�G�_`|)񶭡����K]���3�@zt�q<�~�+6�����Յ̽��Uhh|p�!i����N���E��+Kq��v
�r$��C��J�=[�^��"Q���<�;��Vh�7�9��'��O�����t�x~K���#%���ק��>8i�5{���.m�:n�̷EG���l��k�0�~g��ӟ�nw�]��+
�⤹��I�E�I�{��k�:=u�u})���i�&T�Đ�� �Ԕ*�����R>bEy�|?�����Z5���Ky��R@5�o�6�>^l��2�^����S�h5�l��K�-��#�8,� '��>�`��^1�}&��~�ut�����;�D\��%-YRE��Tw���Ȉ)U 
�{��0�UZp���|�����+	��`�fm�������U�d+s��<u�)>�;�_�4=@�>����dh5	,�-��w�I9j� d�s���q${o	�p#򘞼��ʽ-l~����Y��\�7v���o
�bEw�RF1�~UoŖw��>(�5_��� g]N�kq&1�n��c#8�oZ��u���
��Z�v+�����*�'��=�k��ؿ��ǻ����F�o�����b���� �����q�x�^y�y|l���?E?����]E/7��F䪮:�1\����� ���Z�[���[;�hg�L���2v��$¸ߏv�����x����>�f��:lnU��#��ۜ���w�㟚N�/C7,���\���G.>Vl�<Tʠ�1��h|N�'�~
����7��|;q}��Cr��"��s����M����%����w����-K�,a�V`H,	�G�g�kn��)t2�%;x&�?�ڗ��t)
~�~�fE�:ל?�"5ܲL�,#���C��?��_�&�T�n4�յ{xm�V_�<e�Dl�VDld��c�z�'�5�r�w=�p��D)�-��#]x�G��w�=�;\���Mux��p��M�D��#!�t�k^)����l��\�G�=��!�I-����Bg�#��א�T𞛭���/���[}B=*��7��7�ܳ4�*�Ybeڪ2�vH�ʌ�[]�)d�jK�R��IZ����џ�ͧ�� �i�>�z��׆[{��ı�P��vz珥{W����H�۶��5������H���A� ��h����#GO�zX���x�����w�Ԧ���,��f���ż|���(�jS�����9u���n[<�)£Y-��Y�O�I��$u�}��9�8���'�GM6F��R�{ݕ<E�%�[*�ۍ��0�z�ޤ�5M;��i�70��[te8�G5���If3����5�<M3,���X�8���Wh�~1x��P�n�}K�N��Ki�/5�� ��'�w.
0x�x�'�+� ���<0�˥�"���@���el�z�M|���Go�8d��W��
���H�(4;<d��'��S����gn�uE�Q����?̥7�_���wu7�� [G����ka���;6�r1��+���_�����l���g.���Y>��AQ��n$dq��S㯂�?�~0�?«;���=R95�vx����*����6�g�ϲx{�>�o�e�ց����w[�������(+���A�c�+ѧN�H�N��`hW�Ù�y�
|9�<�f���%���q�.�d�⻵IA �*� P���Ru�~�� 	�fo�K�##�%�đ�e�+H~�>�d��p߶6��|'����_X��Qxr�]F;%Ԭ����+�V\�'q{ܾ_�#�\Ou 2��Q[�QvRfX����(Tm?3��k�/�>�)�u�
�7O��;�mmf��7�$B�F�b!y�}�� �(e�j_�m���9֦�=��eD 0��S��]�iNT�l�p5'R�e)]����6�sh�X2ē��6*A�kc���M���<�k���Ì`:	 P�����H�'5�5q�!|�����d�b�c�n@�~�pGQN������wR(WkW\�I�����<}?0��������;X�42�6�&���.衆�����%�7U+�I�e����k}����fɏ�S���~\��*�'�.x�l<A=�����M������;Ac��ճ�~� �U��	u�c�	%��d�?+v�>�h��;^����x�f���-�؉VYm�77�U�-�9���� }o���v�O�u@�����ح�m<�u��ֽ��b����Ҷ����ż��w)n�`c'��t��7�O�M���T��9&��n.�ѺGU��,>P�+
��R�G��f�lVt`�v��~𦏠�9�'6��7�u����y�f��4kӰm�V��:�c��6���5h-l�C��M�ٴ��	-�d<�ٝâ�d�o�|�����Cy�]y,^�&Q$y9
�@_��j��<�_j��ws�Ws�[��ۛ�5Qcve�BL�O<�k�X�r���|�YS��r�+�ַ}u���S��;4�ŞO����op�fx0����bm5fm�MW#��{��zWsy������1�Sbf�dP��UV���'���3���pp1�Ұu#��:5T#�7�yv���%�-l�����G&q��>����d��8n�u�� �"���'��W���@���D�T�ːŅ�>����x���<)���_�����.��f�N7�����w�O<e���q�����Qhf�c}�YgU~@�I�G_z���b=jǏ�u�� ��}G�I������{�O�X�&+0$`r}�濌-[Ju;���O�4ag|]T��rX�:����z/��h�D��{�#��b�D��2d�������˳;c<��ڲ�"�1�0�_g���M���e���=z~��m	q^_��'�`0+�t�� x9�ҩ��K��T��C`��_z��������Z#�n+¿g�����|M�Ou�_M�ˋ�.{��a����z�q_S|7�6�����\Z��Y'����s�\5�� �/v�{k���a0�%iZ��>L���Tx*�3�n�	)��lW����9xÂ5�~�g� Q�9�<��I��Ҿ�����>m{Z��>��f�h������ V�h#޼K�C�}�x/�6���5�x����ҡ��i-��Ȓ8s\Bea���T1=뚎e���8�M�e��R�����W?
G��KXҮ4�4�g����`�Y���u�im�B<�,Sv�t*A$1�5�����O���U�Զ��i��&�"H���Q�+�u/
�~ ���)��`��t�?�=i�-aW#�j�dyX��F���<�Z�s��c��}����e�V�f��-gIl-�;M��8��rrl�m��Sp�lxY��<�mn�{�vo�~�>���	��熵+'���Csm=���'�F��2R���5�ZW���<+��5u�k+�E-���ʳ[I�m���IPƬ�h,�y8�J�6��SY�>%���7��u#𵞳�è��d�#�cN�ט
��J����j*�G>*�E�Ҽ>�_[Gkh�,���\JT��$��@m�ۀX����{x��e�:U��i��E�9�ڿ��ĭ+IԼM����wh/��2w��|�a��6
���"�m��W�|M�I����7aY8�wv�VPL`�y�z^�|���Sj�,Z����Vk�M2�57�0TIwqUT���S!f]���??c�߇�?��m5}6���d��y��uY�	h��:eHNp&W�VU4��{��
8��V��ݽ�޺�ݏ�h|I�$zU���d�]2���g�$�RA�@�����@��5��v��z�!��~Ů��Z��|0�]E+y8pQ� ��v�q����o����{D�>[i����"��Gg
����$s�<�l3`�¿��χ�k�E׵+�4�X�[�RKh����E�B!�<�!%6��5)�Ǖ�n/	UV�*s�������z?į��o�U㈆�i,6�>�p�m$J�Y� >e< �3��>Ʋ�3�x�����-WO�mu+�`�Q�R�	"� Yv�6z䞜׼���?�e�|/�,n�àO%ơc��y~ڪ�q���;0�@�����?��R�B������y6j�"pg��v,0�p%� �?�L�;���\�ܰ���c+�}�p���zZ��_�����l4�#Q�W���{���r�C)VW�n�����^W���ߵ��{C�X>"��"M>k��"�DI uT�@�`��[�ٗ�w�/x��U6_�aka,����qK%©,,���JF�����v��uo
��;���ڊ7X.��Nt�贐FZweP�g��ya�  2y5�HrFǽR�XYBR߳�ө��>�e��Z��k�gD�'��6���P�X��N����ɕ\�*Ҥq���i48nt4���f�Cy$��F���,��F� N��4m��/�m5���lHږm���U�ŵ��AuUR��T����I�~8h6�$F�Oq=�[��*� hW���yw"�e$��>eb�����o���}�>���M�ir��.�t���5����!�i�eۋN	���� 
��W��_2���� ���З*��T`��I�}5�Kx��Ej#Qª� �b��;#Üԣ�KWF2)��ֳ�1ۖ�j,���F�wl�u�h�OQ��>ة��O:����k��d�����?�U�C(�S�d6�C�oZ�.5�ː��?Q�[�n�5͈32�_���5����c&�ό�=]G���$����,1����?~_���B��`� LT�w�o-�4������R���'c8�һ��M��T�m���G�� ���l�Q�*t�����?C������u��V������͋층���Z+�l�����U_wE8��NK�
Z$R_��ܸi��E9�1��U ���ޜpz���rY���e=�����V6����,�{��̝��g��xo)����w��:qj��`�/��ǖ���z��v�t�6�y��K�]���h��FD̹P�nb�g�l��6�>R�"��Q����T4H����iV�E�6���v���rK;�Ě�a��O5�I���&/,K�>d� ��j��?
|�������M���	�d+r?�Ҋ��  �����X,./�$��m��Y�Dp�BH��b��p��G�ek��7���}�#V��f6�t�g�
���M��9�[������f�=K�| U�4���Sض{WEv[�v\�g�j��\6�}�/7�i��M�l��m�W�`{�3���B�����������mc�������� WN�u����7��,��VviQ�b[�žM�g���h�0~��*����~[�;@[�쵭YD<��NHx����2��O��$��wiv�����O��������&⮭�Ѐ3�����ŷ�<0� tK3�"�`��)�Hf�T��S��޵�}�g�U�?ew�:kY�P�����I2+`� �j� <I�`O�t�A��p���k���-+��Q��D�O��g��/��Ƃ�8���?�����|��G�����(�̷�3�+wV���K����Ұ��̓�;r?:�գ��� my��jbaOH��ec��'��r�#�5#����\�^ESۯ�Qҷ(xu�C�9� K���
�������t�Q�p˧�3����/���Ū��P'���_�>�/��f`[Z��a�>�TR��r�(Կ�� �.>(��}�jKtͧi��Q���*��dTc����x�넻�ѥ���m>9Wo|�� ����?m��'���i$��B�|m>ld��9��xw�;�7UK+�%-��f?�ıe��Etacbh;ꔟɻ��Xv����� �z����fx;�q�2k�#\t��k�%|`�H�zc�&�> F|���+� k-�K��i��z.��bF�	�^s���B{ +Ѭd�j�q��f(�S�y�ǂ�!��3���	%���yU6{���@�n<s^��Om�n-"�̷��k�3�+�)^���s����-t��Hc�Vy�N�ģs��3�_Z�����/5��W�{i䉭� ^6_����Ҽ_��ה$ۜ�����
�eMJ�Ehpߴ���Oþ�Ӭ��k��(w�X5̬{ ���z����o�^$���P�Ҭ�N�w_��W�������0î�yG�5��c���P隝֞/�����W̏���GZ�o�}���'�{�ZͶ��K#����ʎ�\��ݷ�� ��Wp��S�\��V��� ��U<O��ȓ���l}aᏉ1ژnn�Ki�Y�̷��P\��K���of�_ơ�)��Wg×�<6���5k�N�y59��z��h�3���m��b$�d|�9�y}���5���ǈ�%�x�uF�:�El�/�6A��3���9��K%��]ßxwb�Z~���(�mG@M7W�R���Y
_<�L0ȗn�!V�Q��bz���Ƥ\&��������¾/���z�H>֖�62�4Y� K���A+�A�sZ� 	f�kK�|A�iQ����s��k7�k�n��'�o�@CH�[��a��m�O��Y�u���8m�l��f��F�Xv���W}6�w�SO=�>ܻE'�s���Ⳍof��y����/v��n�y���~:|L��e�[G��*�wj�]�m�91�w�~Y4R�:�$��~�J���'�g���P�Gּ;5�̑�Y^]����ǚ�X�����x3�?<>4�hzo�t���T�6���:� )���/�'�Ǆ������x;N�&:���^�1@�{b�+*$� >�8����;�����>�|����K�Ɖ�C�ۛ{8��٤�W'̙d��2��Cn$d�:ֵ�|I��,�V���5�;Y$x'��[W }�*�����:��t����~���=?VӴM9�$i ��{�&��,/��T`���S�ij<l<#�݈�ag��� f�yڠ��2tT<(;ی
�S��Gt~k��U����e��;��V��ӯ�j�;�]�|a�TzF�}qa�h�5����|ztR2��v��ܹ���;s�O��f�Ε7��V�ĺ7��[]��v:�._��m�����4�S9`��N�H�y�_�m<�~=�zu��yob���b�D';�t����.�%�k�<����C�u���i��Z�]*�2��nu�WP�l�[bH9P	���$���x�#��s�{��� �vG�E��w�O���E������k��׺�)�"$������ʑ���Mk�g��}�k�E�Z�o�%�x{P����sc�=�L6n )%203�+�O�w_��w������F�%K���M&{�-�@�B"�q��$�a?&����g�:�<����gG�o���GV�,U[�2A� f�ί���H%[b�&�S�`�&�N3Vg�Y�Rq����j� �U����꺥�G
�^����x���[z`���� |K�|HX/��t��kk}w���6� ��I�gp>EɄ�Ed.	�F.���7¾�5��F��H�z����;��"�\J I
3H�N1�?)c�����KO����.�-d�/ol�Y�-�D�\�1��1���s�RPv�|���؅R�M5�֗��m�n� �H�9uxf�ݤ����q$lS�^]�}G�+�� �'��2��(4�0��$��G��5�7����Z*®�xzs����:+�	���G�m�o�4�T������+��	3�Tr�N=��<;� ��O���Y-��%�<nF�g��^�
�)O^3T���U?/���<����>,���k 6�0բY'H���s�׎~0�v) ����in��1�_@x�K�CfJ��.��������ny�G;�:!]Ӷ��>B���	�K�n%��N���{n��>8�����е�7�鶷/& �^bp=K�+�㦃~��!��ǧҿD�=l���픝��ֱ�� x�v��5*jIjwT���������6|@��{�6LEw����#n�=�t��F'�d�����:���u�^���	�i��
�H���H��2m��8���°�:רkWֺ�?�-{S��mk������'�n�|q)���9�W�x}�XЧ�����)��N�����^Q��G �흤��k���rsu>�+�JP����>h��^��/�f��� �zާ�?���o�ڤI�]�U�%�p&]�T9U;�c#5���!��GC\�$���-Gd�u��6����Y/�f�Yw�63^��ڭ�V�+S�99"��Q�gu���z4�TR��ϖ?�V�w^�t�R��}D�9������$x��Eg�E"{��6�9�m��Qa%�l[ [���㎔W����W>�+_�>�����|���RX��jǅ��7]��x*A�{Է,�j�<���1Y~,�6����k��H�6�./,���5yو {���[��nW)�;��/[�_�Vz�u�{Â�̏�[M�2�T��P��	�C`V�����~&�<Im���$�8���<죁c� �ָx|�O���;������y��.�'�u37T�������>(�_Ě���0�:%��8W��NM����rTg��9\��#�T�����i`s
X~T�����!��]��ƃ��i�����j1B��>�b�7�� }잕``C��=k�?h���!�c�x[F�t]?UK�)���$�Y
� )��niX��S�n+�����FEe������ֶ�4�)���+�S��i8�9�����ڃǷ�/��\�K��z?�G�&[y.<��3)���M�c � <�j|�=N�%mZ�g�L�Z>���۬2�8O0��{�+���s3��������c�ZlV���id���ʑ�1����
�m������F���]M˪`����W!��~��캎�q�GzV5���UD�J���<?!߬wz��tW�ߴ��_x��ZV��3C6�r<F�)@g%]��OO~���Sv����R�Z|��N�H�lX���/���G7��X�����W��do7�V�9e��9=�M{�u��!�:���M�V#�S~ �[��x�pؠ��sO	�� G��ϱ���:>��=7ጁ|`����5��E�6 � �t�����s�1)���+�#���gW�SݚKdW��ߔ���ۚ�kdL�s^q��+ =1���;-��'�V�2=���m�+���(��Z�_c����ᄷ�y듊�6/A�xGKS� �VMh�f�9FϨ�_ �6�<�]�3Hp�pz��^���f���.N���,=(��{��X��U�^�l|��]6� �X�ܓ1���5�G�p�>$�=��Z�+��-�+yO�tN��P0��q�y������2�N�+{Hcq!�.Dg����玘�a��m�=*��E�$���b	v	�U#Q�p3Ϩ�Nkǫ��V�
4��5}/�� Cl&�:�8�c���l�^�+�|i��xr?˩i���2��_�{��,`�q� w&+�ψ�5��ց��.KGב�.�覽��]з���Dn�n�!$�����h"�x&h���a�-U���VL�$��Ӻ �W����p�|��Z��>4M�X�7]�f��W��C
�E�����q�b���g�{*�*��=�4�>��-�	�/xF��~&�E��8�����b2������^����e�Ϥj�ׁ�IUwl}�2�k�}q^[�/þ��o,�ԥy|?��s�ߤ7��	#]�X(M�� *��
�h� xs�_ßx�B�]*}ɴ�h�햆6�+��2�p��kg#5�MG��R�ϣ&������7W6�(�g��� ��s 
�H�_��� jk?�K����>��*�X�kn��˯U��>T�_�l�X�����6��k'�d�K�e��ѯL���C,���Ee�N��X �_�/�����Z$3Y�j����0[Bfa�E;��]�B��HǽD���G�S�Ue���^��m!�֗M����;-��<M8����d�fpd�ɱ�Sb��H�30-_�� �W�}ᧃ�Ҵ�X��%��N��s�]نY�͖?y��7���;�<��k�YV��ͽ��
�f�\�9���#��!��:�{� ��楨�R�ޓk�[_K�Q{����A�X$����兹�{�r|0�֮�r�M��t_����
^X\,��⍊�� py:}G�xO��e?X��V�3Z��5�6[cg}J����&0C���&�w��(��[��R��N����I2��X猀@����ď�GX��c��u�A�]����XE�r�YYq�59�q]�-$��"�,,Z������>
��c��7B�<aygo����_1��e�t�P�i4�+�ϖrp9.D`n�3��vzH�He�^�-�s}y;��J�#2����33>�\ ��:]OX������,QD�}��A��̭/��ZVnM��b�\ >�� ��xV-CX�W��Es��v�k�]CW��9�Q2�j�i��2H$d}�+�2U���\UL瞮���^��w��݌�n��C����ZTZ5���rYƖb��󌻃g�	�dcזx3����?h�|2�� �$W���2��N��\4��ǝ���<�ࠚ��G��������8����O\$�Y9]���3������>+�]M?���ٮ��n$FF�FWH*������V��a��F�å��������5��X���1f�[i��ȷ�&eiX�^Fɯa𭴖6:E��������T�JD��q�ʚ���&�B;m�#�2�� �:ȷ��n���ᑰw���y���ΰ� �=�l=T��Zy3��UI��T����Uՙa±�鯁$�ּ��'�{�k��t� �ݪ� k�.�	6���f����/����W����=�~�_�V��\#+}�J��+;�Z[2�b6a�Z��P�v� ]O1�/�xs�Q��5֧=��Q�M��׷ꌽ�\��}S��D}J�������㝚� �/�&�������q�������1ڊl�����a_��5;?��^��٭��uE�8��Y�k}�c+�`�g9�Es� ��� &��V�����w�\��p8y��x��G�C%���M_��~�����gď���_\��k���<�����d�V2^��!�=���?F�4�xoR���x.f����V%@o*t��|�Y�[��*�� j/�Q�1|CםN��Ĺ<�˒8R}kr����-m	�����X�����
v|��ܜ�9�8Z�V���G/�a��Nk����� �*���E������7z���D����I.i<� �.��
�%ry�K�@�,O׌�ߊ�����>0�����r�PG��e,��J�h�����迵�����E�ځ�n-��Y�P~U�p�N>W�泖
�z���1Sw����g� ���Ac�� �ِ[�Ϩ^���"�_0�Fq�ǯl�ώ�=k� -t��2�.�����C�&}�!�VWL#��ݨ�KMҦ�#�0tg��R��w�/a���U�9��|i��5Ti���wz!X��'�4���+��&�������o=O=O��4�@�%��}�j�|���K�-��FF�X#�*�FGt���rJi��˰�<De=�{����N+K{v�k�e}0�Qpp3���鏧z�� �oV������Zj���i���Ězlt�M��F�E,x���rZ��9�=YS��Ӯ\�m"]J��0p<����.�v�r+��.�Y�Ax�Imk��xᆓt���תɨk3�n��G��Jy���rk۫^���?I�cC��2=>�j��o;cUa�p;�Z���+k<�n��E�T����,,
�+��up[;Ge��W�|X��oxv ���3LXz�_�_=/#�LEE'Rp�?�9��N��� R�1�
��H�KQʙ�O᪺,x�d1a��u��w��-(�aJ�2�t���l�q��z�֗ɐ�@╭�i玝j�٫�c;Cڭ�(���~�(��?j�5/>#C#����l�{��DO.�U����_<�њM��6��w��L��Y� v�(����~_'�f�a/��'���7I=ԍ��	��x؟�w�� @�z��Uf����@�k���lN��~u�����C��j�?����� ��및������<�&���~ο^��� $��<�U���� �h۵�X?Mǚ��tI=�_i\���<7k-��q�C%ĭ��'�'�n��kk>���	 �)&9����z�xc�v�q����\xhj��"���I!V�ʁr8�O5������>�ƫyo��jZ�v���%�L�[y���N}3_-,��nU������n�nzK �>g-C�_��&���5��F���B����j�c'�j��C���%����Bp���|���u�n�5��)�-u�r�C��O�-�<�\.0�z0>�k��]wĞ��/,^�F��u��	�]GPq��_/W1���%Zܩ������C4"���<�㏎�t���:�3�ۭdVȻR�
 <���05��ğ�@ڞ��ۯ2)m��$�#e,�D	�$�5�� �����^"���v1ɧ�Y��>{�,�����TW˞1����K��O��H�P�Q���vӑ��^~[B�qQ���뵶_5���:�/�Z��ZNh�����N�J��i��?)[Phd[�6W�q���rCq_�T�k��B��º��Z,�<�h:eĪ,��a~r#H�X���
0:W��?�����@�I`��Lחk:��L�n�ʫcp :�c׶3ھ�Uݢ�?#|Y�[��y]�� ��������|g�Cx���޼�x~IoPi!��2\¬|̫ ����x�ò�|d�u�����t=b��L�m����e�EY�2��F\#`��N�p_���4�^!�w���-Z���t��U�[�Jѹ��l��ѣ���\T�B|J��W)��}B�{ۭ�2�4�Yʀ@A��*���i����[�����8�Ž�����>��K�ᶅ�xGQ��T��n���M$�i �,FA�n*�ARQ�S\'���m�Zx"��TУ�Ю����x�H�p�8�q%�Еڞ��?O�g�U��]�V�"{?���m ���˯�B�C�1�$�89��E|H��Y�x��_IYR�K�g�/26�ϓ!(�Q������I���N.��o�� ��g��o�nW��}�Z����r\!�5B$�&6i�8`H��N���|=�G�;D�wW��B��5u�Y�uG-������>��<U��_�P��T�Y��I�FUc�.a�0$>T>R�� �z���ǟ|=�B����/u�nd���#6�*�2�#eH9�\��ʺ�)Nr�g�0��j����O�t��w���K�x[�����}Zok��}�73M%�1[��H����
X.@'��}��?��-
���&��i�^}�;M�M��eRn%�[͑�d6Y��#�k�o������(\i�� gZ�dY	]��1>���<�o�>��/��ǿ�u[��m�D/�6�ڍ��nc�s<n/��5��ٟS���[�����w�iwK�WźF���Y�rhw��sMh�1�\JТ�,�2�Y�bJ���?��u�|;�f����IF���y\[FSh�˖ߖ=3���ן�Ϗ5K[�v׵xE¸�r=�B���z`��b_ۻƾ>�<'���ֺ-��u��%���]�JG�H`2G��d��,-j:�S�v���$T��+X�����8��@�x�XZ��������r1�t�֥o�kZ��B�(nn��5b2ܲ��8t�.#��>⸴G�$��:��wW�⧷p͉���i��Z��yӓ��j�%�9Ȕ�"���y����h�=8c��� ��r_ge�d�F6�J��[���9Sqr3��� G�ͬB��n����Y�״Y�d{�O��TB�,J���0�<��2� �Y��h+��f�^Amyn�k��hЏ���#��Qk�[�լ7�;w% F���HMĒ��+�6���ʡ������x��P��2>�&29�?�Z�vGm�GN��L���B/���ңF�ݚ	*$��$}6��\
��8]n���b�Y�/��r0v� g'�������_�n�Q�V�t��[k�WxU��q�w��~�mB�K�|nUP�����}N;��֣�#������S�{�lg���`;B������#;�Q�H#v1�N��}�C�{4/%��'I$ʿʮ��H!Ԟ�"ۭ�v���y���1��D
��*Q���V�1Vl����;��H�T���!%�h�pΘ!��T��w#��ѩ��mb�K+�[K[��ec� n\*� �ѫb��<��wT��5i# �$`ĳF��x�[qMQ��g�#2[��l��%][i���a*`� ?�B�wi���A)�@����>eB�@� 1�;�T����Op6�oj�b�ŶJ1���#��1����{ˋ��?�<�.��y2�I����|��1jz��z����{�H��h�|�n��B2�9<�5����;i�g�]�o�o$v$�𛙣�` ��9'��K)�[>��b�؀ǇY9!�6��۷��\V��)�f�� �����c� ���^�Y%���W�<�~��U+��(�y����~g���둾�wh��'{�rw)��?_�j��u��(Ys�~lw=�Z>�E}�?��'��_q�+~�����T��j������m/��[�kZ^���G���H�6��r)��ON��;Fy�[�c��<���5�.�uI��X��\����a���b08ғt��g����ic#l��l�T�YO|~��� ����K{d>���Ke�.8���[�x��u�6��#��g�� Z^I���ėL�HG��t�y��k�S�`��v����i��S�r#�|`��
�P����,�7�I6����LčB(O ,� �}2O��ǘ'�Bێ~I����+�~ÿ~2@Wᯋ�|)�fR�i�K �Ò#�_t�9�W�^+�}��>9�|#�,i^#��d��7�t=��`G��t�uke�j�t�G��ux�6�â���q�Ĭ8��F߷��G�ji�"G�-�� ���wጾ"𮱨��U��ӄIkm���Ȋ#h��,����oci���6�q������+�WX�S�[�m��z-sr X$�Ω+�����?<S�^kV�Qɦ	���BP��X�R�֢��$��� Dz 氼c���D�H�w+�9A�U�*z��O�� �rҧ�{�֋�ιS��r�Y\�� ����},ݟ�k�������u�\[�LbwC����||K]FA����T��߅�t��2��V�]+R��m/�W6�k�����X�*�I�
�?|F�l�;h�m�Zǈ!�m:���ѭm�m��V$��8���{Am�l� w�~�N��q^,��;��.�{ۧ����Xʊ�{���8�P�|n�v&]=�i7 y+�k���Ɓ�h���Md�r2������n@��7dc􅤛�;s�+��nM������l2�%ʝ�;� ��F�fԭ�~X*ΌNy�3��w�I� 	�¥�y1�r�G�s��O7�,�� J�=J��/�5,��UN�s���_5�
��ƭ����O#�3W[+�Iç�k���³���o�I t� ��3�y7�$Mid�o$wN�r� ���?�|�� 5�:��Nc�#�G����q^c�dk{l�U�n���C�pO�^�X�&~O��_W��0oSǦ�{�x�I�L�~�̜���j��C���Plb���߭d�-��m\�s��ӱ�H�ݡ�.���^�PI�C�G�x6��}��1���K30^3��M�ƿ2��ǯ�OΛ,P,���<��J�{��?��ɴl�N}�ێ�g^�E�G�"mC+�Y3�6����g�-���`�^K��l��8���\��׀h���������p�0FA���w|�+�� �����2H����Xՙ�q�Z�C1i�ws��0	��N*�a��g�WK��� $�������9Oھ�%c��R2p��Z��aq��~S�}k���׈����Lt�Ƿ�'�ˊ��S��G�D�A�6{�B��&?�1[<��8�n:��^J��k)jWh���T���*�A�{�4q��O\}�UtJ�)��&s�o5ζ��i�w:�����Y���L�2���Qԩ�|�j��5�c� ��?�c��^���<HF�$�m�=w�q$q���_�W�7��KŰ�>4�lq�k���(�Q��Q�&z��(�+�~�Ü)_BU��E-6��_���>E_���O,k0!���US�����èxgV��{+�g���#p��;{��G�����X� �n-���91$*�A��¨�3���s���5�|o���[Oj�.�N�fc�Υ��,�3'���W�c<�>R�[���w��[U�l��G�?-��r���p3K�����P�7Y](%�Tg<z��-b�� 6��ߗ�'��<y����"������.�-h�k�\��K��X_� }1���s_1]"�_O$0�5�<qGopH}�!�p�
�*�NzW�G�G��ֹ]/�������4�I���x���qgz)�ˀ>c����K�f�5	�rϽ���!��RZN�� Fr�i�9��M.؉a#TdfUvV@\s�*��c)��MZx�-�̷+9V�Q૝�2q3cvq��r:Q��g��o,1�k%�R,Fף+	"-�ۋ)����Q�04#���|�Iw<ae����ͽF���"�4���j4Y�����>�<�$H���  �I�l#9TQҦ��=՜3�Ebm����Y���n(ь1^Q��XlA%�ϣ��K��#@A
e�r<���Ga�����-�{Q���+ ���X726�خ��8 pP<�r��~�+���29�$�?˥A#K�p�a�:�ۓܱ��ڮ��)) 7���8 ���<rzTWOn��l�{�!��ʌ�h����fcF�e��F�1�;~�<~�J�Z��̄*䲎�����kF�A!�~c`�V�����<�u�A%�6�J��<m �$g��Nzg� �6�ܕd�
�'ҽ��_��$��ƞ&_m�;�=ԊJ��<���$��J��>��IJ�ܲ���_O�^��=jW6��F��#��$�xVUU��g�;Fݬk|��J4�Ӕ�H�� ���E��߁z�΂t[��VqZ�z`�,�3ȱBX19@\��,W��5��[U�F�q�j�w���k��,�I=}�����ù?k/��Z�l��jńr�\C��;�+4�23(V��ڿ<u�M᷈��i�f]%����|�z������mE���#j�?���L��~�7�ഽc�	�(�z��0@�8����~:߂��K��mt�r��|;y�Yĉsl���+*���1�� �~��#���K�W�%�x;�����l���t�ူ��'s2���X
���3V�/�_�7N�n49ud��o5��!��I#�c�ny$PH�m�*gm_��wМ��O�<�ྒྷi�x�� A1+�5�ݪ�
y�Ѹ
�!�1!��SY��g�����b[U��[��[��?uU@۞�df��x��� |�k:�I�~������9nF��_��#6�0#9��ڣ�T���/�Kk�3O�x��d��<Q,s���d�p���lyq�6�D����9eK�k�cͼ&�u	�`�b�]������$�>�
��W��t+��9�����ܤ��d�$;W-�x�d���\?��l~\V�zsX�6���%)aT^�>��}<���A��-�5����D�\����?�}>�+XYDq�/��'�j��sۊ�cdqʍNǰh�"�9$q��l�oolH�Ny��-~)][�1�^�kN/�Z����2m;�ZwW1tg��s�g��?Z�Me�4�>�rK+L��澍Ҽ+��ᗻ�J����7���V\�p��5��m�����|-�]R�M���D��I\|���^����)v����)�.c���i>���n����v�^%Lf*N^Ξ��%�ݞ�,=8%��d�����^� ������-ɖ�ʀ��2W;��q�1�_>�b�[}~����� �T޸��3��O~��'�<Af,'���ᷴ�Fb�'��X;��خCM�4ojwW�T�2�(�a9\ O�#�;:�y��/�1i�ՊI����>$�J�_Zq}�����uzy�{���n��G�����#Ek�DŔ���2����kڼ/��|�9+}:Q�9���5pWZ8�7wX�R���H�)��G�\�q������G�Ӗ�/��g�#j���p��/�����1ڭ����������Ꮛ�?��]Z��uX5]>P���q,ko&T�ħ;��(�������Lc�Y�xu^�u	��y9�{���G�_8��S��d~}B)t�V�M�
S ?�Y��v^���E� ��v����� ?�S$� �V�7j���a���s	#�o*��K���Y�B���		X� |��n��Y�����>2ʼ���_F|K��l>�R��t��B��ch�.�����\* $À�8�5�~=�ko�+�:�k�l���#��z�\�;���@�^c����~W,ʌ��]-���8 ���;v 	�f� ,x۹'�F:Wڟ���v6��@��0��˦�8����#�-�B�o_ezm�	$z��ҽ.d~�c�XLj�O�W��x�u�+��n�dM���@ǹ'�W�	_�8�Ǘ����u�n����������\x�m^xuH���[�\�v�͓�l��9n�T�K���̪Ɔ�Y����t 7�q�¦F\�?�����}Ż��X�s32eT��� �O��z������2M�/����L���K�\MoߑayWw�v�[������t@q���s.��t��/K�e������u� �P�[���6בi�8ekHa���w!���X��oc����绅�ԥU�NqW������o��+�G�b�?h�^�6#�=
�Mҭ�unnI.Tv�D����Ĝ�^I� T���Z����-Z;-?�>WS[bT^M,�"@�$kB��|��=��?����u�[o�P�Y�;	�mXm��>S"�Q�ӯ�G� ���ώ�����-���{O�j:$�v���pD/'˜�e�+����3�_�jB�UBpw�_^������9�D���G@䏨����� ����x��n���۵���bu��'��$(�]�k&�T $�9���� G���$ڴ��XG�dN�{p
��]��z�`��g��-�M[��I�\���O�E�$(��8���s�V�~��K{�6� �B����'H��.���6�kՉ#���29�����q�|3���&�!x��(����L��r2� ��� �1�����W�,<}��Z��J�U׈��j%c��[�,%9�-�q����!mh�I$:���W�.b��@�]����yd s��4�|�2�ҩ�r���J��fU����4�"g�@�P.�/�U#����?���-]�ٔή�U��R��،1ݰl���^hHnYqb9�+�>hbr�М��;����]�jW2���`�26^&
�t���Eb7v�+[��kq��|�m��0�"��bW|e�Dʂw�����C�����{HK=�ْfg($1�2G#�2dTx�� IRd�tVz������V�(�F�XY	.ˆh�z`(`�F�D�B�.#�2x��$.�*meh�0U�s�<e���s$�:��"|�C,r�W��9�0}NQEX����kw�����Iybd�1FV9���/Q�pPM�Fh����N�3(Ǩ
1�c��F:dt���Q���)�և��I �C�󭈘Ȯ�
���0�d�u�#Es��1G�7;)�c��>��RQ����L�18%Ÿ
T��2W��s�d�r5����"r�y�,	��� ��N*��5�Q�B$Q�����t�����yf��%�1���?^ *4���H�T|Q�2>2ۺd��� g8�� b�7Iߵ�x������X��|��׊���O'0��S�O�+�����<�5�q!��Y�ް��M�����0�{]3�>���7���-���lR��\� iC'�9c��̑󑏙	8�	�� �К��-.��G�^�. �~�um�kfc����NUH9�~`����s���c*��d18P?*��F���N�`��������iU���py�&6��ף_�?I�6|u[�` ���@�@��Hc/���pX�?�|tPN��~�O���x�Y�&���:���*C���VV�1�I��5@N9$�Ok���8E2^��pEmxYD���s�]�a�|��֝IJI�K^fx�^#R�\���椏���:/�l%�ò�֒G���]/Ux$�.n}�-�(�R�qR��a�pu���]�ze惧�������I�5%K(���2��r\?1��a�p�|߯*� iv�%|ͱ��z
v�3ɪi�;�<����r_*A���S��=p�R����~ަ/��}c�W1G�+��3��tR8]�"�U@.�#������ �W�6���=0�g"\�~�#)m,���AZ����9�i9�k6���MזkI嵕R@�B��� G�b�'֜}݌�d�d��s����լ�_���J����%�H���H�� ���x�����R+ym!��x�ŕ����o����2��<��X�Ɗ�o�kjMJ������u4�ڤ�Aj�R<#{���f��'5���V�+�� �r<e�K��jv���7�|����m�Y7'!d �⡶��V�~k�N�}��:B����^�{�t�J��e�����ю�&� �! `Ts�a��Z�0�/��O]_�\�\�D�34�#Mꉸ�v� �  �����p�������u�U��qKk� �M�X>T[<�<9���/��`[�9ՙ�`f�b�5���V�Ԯ4awyqt-��[x<�Y���pX�'�Q��8�:E�M���&���3�_��d���&��U���=�������5����<?��ma��f�"r�q���������_<��N$�H29��mZ�\���\��9�s�>�F|�2�\dy1J=�/�h�'��g�O�_�=��R�t߳"j���H�_��p@98��M��ݗ�+�`t'�rO���|���V��Q��T����8������;�B��"��
�08##����K-���wA?3ϭC�+4����_'�*t�$tO����x{���s]<�N���hȈ�6��K�߂&d;eA �d
�Ѿ|G����][ú�d��X���6�<���Z���BY�
�{�ּH�[�S2��U6��,>��Q�I��� �[��Tg��� �3�����"�_Y��������#8[��-�φz}�gr�i�so/������Y�m.�S̾z���c�3\ƽ{p��O(%�O�y�U{�� �'b��O�^�� ���wZ_��RuyuO��Đ�i,�*���I8�I$��Tf�G�[�Q�Y�l4O!tn̠ǌ�Q� ��3�L�"�XnGJ}�/گфF+��<�=+(������Ŗ^��';w�#�� �#�o5/�z��][�������fx��HQ=y稪sY�Z��_�*�`�mV�ܷ�I=}+�m�4��Y$y&�7gbK(~��j�f�My�`H|���b󎕫����OK�9������ �3��H��,	?�!���р珕����V�����KC&��_K�����+\<Me]�b�юrN�3Ҽ��m�o�?�H�OL 01�;S䳷:�H`���3�0�s�\�JM;���&�׫St�U���8?�H�C��c� ����㯖��� W����aĒ�� �<E�#��.&��6�l�U_��ǵs:.�d���i9�2XĤ���*Y4�&��;r37R�#�cM.�w�ņP���T��g��\�o]�R�+m��w@� :c��5��FC�xU��spI��ׅ��w���m0EF�� 2�c �8�MAD��f�BUd#,� =��*|�:��]�s]������E�x�OKY�?�I�47v�s�b�cX���r01�>��3�H]&��ĝGCmYb���j_���*-�,�s�C�A$��4��K0U�/!�s�\�*��j�r��(T��F�03ӊ�7Q�g����嶆�T{r;�g���f�d]|C�@�f�����HP2N �zWϿ�.�|D[������h�)��������2w���2Hʌ���t�)5�^�݈;Ah���J���vQjP���@��,J0ޣ������c�Pt�UAu�]��M����խ� g	��K;�`մ�X�F��4����̏ЯN@�������bDH�f^�b�b�ˣ|�́�nM}=�@�7�Ǉ�o���mZkf�)C./BFO_Z���o	�+�y|�_�a����3�\ 3�+���zy�Y}:<�־�����}g*�4d*��h�����e� ��<�sE�א���2��$Q�-��b�U"0��y����S��x(��[N�oޢ��U� � P�>�zV���o�	 ,:��5nB)��_@@J�=�Z�=�P������ePw��FM�2�,�J���%����[P7���_9a��}�I
HF,��$�v�[uٷ��5�.�ăt�9H�y����v�(�E�v���7%Y��X�BH���kƷ�I���i��ZO*]���.P�Շb:��&�����y�[L�WsܪJ̢i�,�X�������n��PK   yXv��^}%  �)  /   images/16ad4ddc-6952-449b-a843-6c6b0f91f705.jpg�zTSݶ��(��J���TQP��JQ��
J�.HED��"�A�� - *�K轅�CH��_��;��OF�H��{�9��{��FB&OG5U5T** ��� 2
x	03b<�����x����Q.����GϜ<u���9A����_V�"|QV������,T��M�+Z�5�un�T�:D��t����'/��>s����M �!�ا�:P�QѰQ�[�2)�~]��5-=�.�Q�������������ė��e�;vV\����C�s.�Q���K?s������5�����S�\�/
	_������v㦊�������{�F�&�V��X��ڹ=s�x����2�U��7��1�q�	��2��g�����TV^QYU]S����֎������?084<2:=3;7��������������P4T\������������*��?��ҝ�?�������9��C��Q�������x���t�����͟�~)��	
��R���?��G��4T��ѰP`����{0�D2���m@�7���]u��`̭�B�(>A��� �[Vz�i8W�=�Tt���L�1�mN=�jHC���!��[�p�F��/��Tه�U�X%�1��a܇�>����p�C��+�>_��j<�=��^�����&2 �����Xj��A�
�3f��d5
yb�zK����I
��hܱ� 5?U��ϳ�u��w��% &nоQ`�����D��J�4g^?խ�krɽ�H����]�暃Zo)��9C��vtZi������`��0fc�ь��u9㗵l ���7�����s����գ͕�+^�1,�[��b �o4@�,�`E�a!��uʝ���kL�.E�?D\��J�2�VK[���'���]z�����BF���	�c2���oA<Ѯ�z��uImJ���i/��Ѽo��!I��y��a��Zl�Ъ�ᐖ��uZ��|���a4v�f�ߪm�W�#����+k��D�O�g0T�0�@�I�g\}CȜ�Ͱ�
� ��������X�4Nf�7��R�M�hcOKK�OH�zQ������v�[���b��U3�p�#�y���E.�\����^w����]mBˈFCr�������`n�i�R"�feWa��
L�Y��/#��Ծ��S�0-�75�~j�=�nq
J��(/����@4��k�x ��ǘE!�����}��B�3o*Ǽ��'�S,sj����\lB���_Q>��9棗o>|�h�u҅u�����[����,J�,f_(*Pss���~�������Y�Ӟ�|
_$�hY�Z�l1�Q6X:��dc���(��&^�o|��;iM��*�if� ���f�p�f/ڶ�A̖�C��)��t��n@:��t@�4���q)�H��7ɿV�Dͺ�E:�J���ɀ���������Bl0Y��x���M `�T#MJ��`���]�8
�[)�e���M~�v�����X��~U>T�O��j��o�n�&�!B��(�1g#!x�A��VA�������&��J�rq���-꒾�z��TG�;^)3�_[�����( m�"ٽ|ܺ���#��R�~K�R_��(�e,�8�Q+^Q�Q����`����3s�M��,9R�u���^M��E���*��u<`���������o����m�mj�b-��+*=��� �뾆��<�<{�@��G���[�aal����W�-���-���!����^2Ь>�C������ d��a�q����	�`�o4d�\�٨yr��A���*5��3P��h'�@	�C2pٌ��,�)Ƴy�>B����Ӂ+Pu=U�[U=��4��٣�����:,�8$Fa�hC6���TϜ��Y�Ao_4x�''�._����zTA��)��\�Geo�ܱêcgo���FR�ʔ����x�Xb��ΐ.ݿ�'�+gl���$8�cU�lOd�Й���s9��Z������E}�c��tF�7O�������x]���H$O?(M��Or'>����LCH�"9A_<4Dѕ�w�.���ߝ�:0� �fp�3e�)�Sم���ߌH7�X��w�~-��Kg�V��p���̬9�y���cI���>V���~�=U�슪2�>i��*���"��Ǜ�W鍢VV�4�-^�нi����2��Hg�����"l��;��*���w���ۺ7*٣�5�;�>��J��xN�<���:��s8�1dзΩ��0�mK�	�t�x�e��jŏ��4���%�Ĵ3�CK� yJF���:bv�W��z���U���T��O�ww�U�e+�}i����
/�\v��4G����F!@���M	�C{�N	��X˺�1�q(�p��{(�lRr�Z�L�-��UҎ�v�J�[8c*�˖L:��Z�p��j��Ju�[F�\[� V�w<��LL�,��Qa�M�Pak�6��)�ʼ�8��қ�oYjz����9{�^'}��s6���\ץ����j�Y9Y��U=�og?�N�rt7TO-~P���K�A�}�����u�m���$t��+$�BS�]�)�b�A�U"n����R.)���D����N�j(^aa�+k�J����'���ߦ�2~M@����@������{�͌E�'���#�"���Y����NH�r�.��,��������*���7sN�ŕ��QߗI��ѯv�����d�	�Rf�,d�<�p�KąR�S�֏i�4��h�U��h?��R��x-�8*t����s��,U�/�n���l�x[{�\��oyfȀ��u�Է��ru��䘸������d_��z���j���G_(���v��Q�l쮠�x���G�N�{�1�Y��Ƌ%���k_�Z�����T/�\��Y�[�ِ�r1.�5���0�;�6����v��QӷR���;��Sl�C��K�_#��"�?����}u��;�2�q�1��yw#K2�N!q,{�]�TY��|�pC9�`�S��C�쮋���>�w�.��<V'j��pVI��]��X{Htil�;�3pY�����VW�CV VS9�L7��h�ʕ�Zr��a��K��@~W>��R(����;��y*��/�ѐ<HT8t� ���ge��|{�^6+���1�"�ђ���w #_�� ;e��2��恦� �=��+>��I%�͌�_�|�����ؿ�z�m� �c�:�
�����24�N�X�$���h�}�ݲh��>;-�M2�ū��3/@�9��`���Ն׿��`��ꙿ!����d aM���8��iW�!��جO�
�K��J�=]�4^C�
���b�0�_����L
v���m���Y�z#�Y��9f��e0A);�۰&C��(v�pme/b���ٲC��n��ն��]n-�C�O�����_��E8�D]�d7y��6'~�Ee&����~gqB��F����`�dc��,q���G�,C@������z�ڧ�d�o�_��<��l�;䴾g�F�FE�Uu��Ă�a#g���^Y=���5܈y�;��:�w�������g�Y�,��z�ڙ/��W��Z}���t���&*'�#��V��|��(��r�� �	
�e�� ip�¶��od��6S��˘5Х�Մ�5sD��@UNbxv[^��~Z�_Z��ٜ��'�c�Z��<�I��Űh�����E|'��ݷx<$��!q�	9�S$tb�W'0�����>+GH��'ӹ����tUO_O )O��C�nG2|9&0��A�~��.]:�}���{�Wa����������/,n�W�����
ߺ�gE_��B*�H0����P�6[���{��n���uQ�*��
k{�hZ�Qh5���'�J y�!�v��f�J��8���b��"�l���"h�f�AW�b\�
��md��)�s����:�<� Ch��֐�U��$�!�者y�͸G�)֥g�z�J�L�:�j�&�lyLP�zq���ca�~�%�W�Fm���1�~��9S%g���V�q��F����c��^��X���T&e�ڑ��՞t���_s�o�-��I�u��"���ضy3��GZ�k��H�+9�wl3S���?j\�v��T^���@ً(��d�*ݍ�M�{��9c��^w6?.>��,�x��g&���$Q�9d�c�o�Þ��gɼ:�;j~s��#��r�2�h��ngF ���G �X:V���c$����֜Pw��k�b�\�jjX�r��S�[+��o�M �se�رk�4�����ڈ�2`G�z�e��
9W3���}���x;��#�pYe����3F@p�H;ج5Ս�JE̷�E��w���gB���T���t��𡏖��a�����t�)jo\���5̕�'::n�,�Xt3��9�k�������c9i�Ë%2�eJ̦?�����N^��|���>�TX`?�� 9��t�.4�����m��o������&�׈������"��V���xǹׯ��\�N)@�Z��!�C�3�%!]�h�,ݯ[���mO9X>�ř��Юm�n	���8�;��+��!B^�*�sF�)���>%zyM��c���2�_�G���na9P`U�y�j��������)�J����@y��y�}��Ɖ���g���Ow~	���G\�;u�'�+ӟ�8#y�V0�:��5;�y [#�+/�-�JhW$Ĥ���Q2E{8����Z�4a;���J�o�z�W���I�ևc[m&����G.W1��,��a�8C��k=��bR�.�)�p�Jw�$q.�o1a�nY��L\�#��-Bw���������v�`���սϝq{�s�,�mj�ɘ��QI�V�ԍ����]ν�xtƷ�����5���/D�k$�27f���*�X���o:+;ɶ8�𸠍$�.%Y%���[O��F^T^�dd��WW1,*
G��-y=���â@��ϩ^�%�tri{̌0�N�)�Sf�����Z�7�f�n.3�����WZ�^1��{OA�åo���To�U�~'�m�:2�D���!Sr>㪏k���
i�i�n8��=xf�dQu
3�^�1lbdF���߳G(Ι}ğU='��I��ftuf�q~v�AoF��<6�<R��>�:WpF��Q�����$nr��b�U�ח˴i
J�b��وY	�+��W¿\�9�2|PcjS)��}�i+��_�E���E��N����y�>Ժ��1�%v=&7x��vs�g��.�E���-H�n��8D���804z`����#���D.���D����F��j+�kX��[�x۽�
�\wD�Xƞ����g<1�ׂ&9����U�ow�>]u��r}��[KL�Z{ݳ��J��Yj�w
���e&��9^�%�ը���W�A�|�J] 4D##3E��Y�ğG6`�}v�ee���I��}�ߵ�rU!��@/��Jh�A��KT^}����VdgZ���b5M�BX��R�`�d��R����u�nr��
�i!
v���4�#�݄��L�V��,D&�^;�D��MU���t�K��ƹy��4 %�d���DS:s&�;�F:�z��{��N8���tS�^/{\�B�|�)�$���{�����|Z�Po]�҆���J������_¿DĭDN�X,mjO��N�5�D:u���>N�Lք��Bl�N�9d9�4V���)��g9�F��e�W�p����tx%$���7�h|�Dx�|�~]|1�n}ԍ6��ׯOT[P��Iy0L���F/wۻߟ�7�ҥ7t� ��Vd���:�䣉J����?�U���թP���O�]��k�m� �ޮ
�
+��(�V���s�S���[��X��K�t�ۉ6Bc��j���A!��Ƕ���V+к���Y�΄�ƲNʮ�����m`���{O�ȸ"KQ�����ǉj�$��z���HĘ5qE�\�؛�8���y���۽�z�ȓ�4�{{߬<��*���_�{%�3'UΓ&�!�4�	�R����c-א�PL����m%J�_���~yKm$b4��;z��1��U�;��[K�#'����y���~�A;����	�hA�0�kD���O�'�Q���P[u�;+9/���u�w[�M����?���>�(�����z��:8H������N�e4'���� �َ����}�-��`�,���X��V�L�hA�l�צj4Ϩ�d�iH̏��s� $Hw�>�f��L����+�����D:�:S�&�����.4
��.��糥$h���g�6s�4���T�������e�C����at�4b�Vq<��(����ͻ�:�z�}�<V��N�6����\?��똎:���pOsg�ʖ�,��Y&	� ���Pc5և�J�Id6H�GA"Ӂ ����9�P��~���K`p"	���y�@��Z�2.@R� w��DZC����3,n��&20S�}}�ަi�(?���]Q�W���@Hj����@s� �8�E�w"����j�	#��2�փ���Ϛ� �m3�;^��k�����:�K	GRc���H��Z����l�ǈ,
��M�]2&����2��)X��pAT��仆����g>�qAe8�����M��W`��@�پi����[�1?��x@�M�[��(NgG�&�5h��%�M�?���8O�3�I�iV��n4�|z.Re^Dl�Y}κ�ծ�wr~��������y|	n����<l����ԙ��LMf�a���jՔ=�WT�K�e�I\b�`���1W��0���}���žv�������7�fO;%	I
q�RݑϞc�1�EV�N\3uL��t~��iNl�V���K%�`
�5�غq]�b\ 1C���4CsB�������� T��.=��R��hV��}���X������c;�U�W����[�,��J�ݪD���uh��/~�ʡR�ml�zKZl�z�*�ۺ7���}v�"'����ٗ��N�+��|�hT�l��Lw6��SB��}�e��D�!yK�����{&����_���:I����8l�,�bl8�g���qfxy��W��� ~\�ޗ_�tL-6'�*Mi�Έ��Pfd �=;�')�,X���N����4.»� ���Ǘ5�n��H�ǆ"���n��qS1'�f����U��T󂋴��r��RZN+J1?������l�;0-�|S���t��ݬ����+q�_�$�狜���c��U��%�p�%f�#f>c�����-`��2��{P�37�h�ؽc��ر�
yX{a����	���d2p�l�8�M��?�g�OLt-��]�v`NM���X�uW0��5;	�d�.ɽtZ[�����{�ﰰ�NE\��3�ڒ�Z�&n�����\_�j�To�:8cF�-�2�x%��bf�Ϙ���tv2���{R��"Nn��mE�4:���~ك��on
�J�O��>TBf�$B��|"���;E�a�n.|��(��-z��Z��Q���v�p����7_�R3�2���E,f?�|HInpO�ڰtq�a�+c6O�6yQ�"�mJ�6��uqؐ-v�W}$�iB0d����*���nY-�b���Ff�I��1�s��Aؖ���μ�`��� %�q��?�������'��O�d��#9|�	Z�E��v�����E�9��_H��؋ ����B���$eچ��,R����ɟ�?l���W�A�.ʰJR�~�ǐ����N�	�s?�p�֢4E�ߩc�K�Wy��m�y8գ��������N�-\Hę���
��I�'7JTS�'��9���{�����b��<�>9�P�f�_�$n��|U����P2P��AR��U�wSd����	��z}�l��R4)h8�$\��t���.]�:S��-W�uz[#�Ψ~�y��<;���^빌<h�����$:�c�8����I�nQ�4�^��t�V��1��[A�7����A�Vz�}5�0W���=��,G9���-}}������020?D�#�@(Ͳ� >�D���~����?d�zC�!P��O|
��&=��`�ؽj�C:;D��%����+�n<A����Y7|��C�V�\y���5��m[��K�����t�gk�gk��M�tE��0c������N�3��癱y��6����5�Hm���G1��bjT�r'g,7߈4�9���M2�,zKw���j0��?���.���.�^�hù3���:QIӈ�)�
+��E��1�*��1M�h���)2�[���iqE��OЮ~e��X�"�6%1˓;��}2�:�2��\F���Ug!'���Ta����R=^��K�T�!?���"d�s�7\�����ek藭�?�)��m#5@J���_�\������i�w��
ptc1���lx�O;Gص��:���Ҽ�
^S��s�$h��ͺ9`�~��"�P
 >ѵ��]xދ�BĿ+0$�a/�W��L�-�N�!�K��b3�E:�+GJ������/7���]����x�j��k�؂ք��پM�?z�O���?F�/AЋ�7����.�^1����x���b�<�x�i��VU�R�r9W ���[ǔeM ��������*��,jm���Rv���V��ϵh�����z�>{��s�����[E��
:c�Bn�7v$�;P�8o���
u(v��%��֔��Wt5�*��;2�Y��I�;�s��63�U��Z�&v�mL�递�|)k� ��ԋXz`A��!�~�1y������D��o�R�l@�gw��Š ����#�@�T�{rI�S~���t�O(�!m�� &o���>CI�j	�Dq��(����g���|������!���N\�+�D9�O�D;��2��%����"}�Y-+r�+�p��������1{n���P�8�����o$?�V����t���J�{���H�uq�>x`k�s�	�$]�͎e��$�⿃����o\_d�ܝ*����м���i-�������*tz拠�_�9#�/3�_%�7�5�g���_��eɔ:Oq.k���/��{��fCįA��׭���m�������~���1���z���Cl�|g�#�}��_���ڞ�_]�2�eH<�L�%�p��އ�f��I;��
u{������{��MIy#���g|���,��g�%`���O�w�<�,�-$t����Qn�:<�3SE�)�>IY�����Tw﫽9/Xg����B�Ǫ��"���%MLZÁ��Y�2��N��KUMN�w���K���s���.��B�r1i�x���]J}��.�QW��M5	�Q��ӼR��"싐`��f���;z׃3�C!�t��3C���T��챷�ڼ��?����4��T؁����23�!R	����Ut�������x鄎�-jl֙��}�0��|v���Y�cI�7V[Ur_=?�Y��!��q&���e�"kP��A�乏��!�_���ީ������G�PK   t~�X@�Ǿ�@  �@  /   images/20309cfb-f1e5-4537-8027-12bfe73d577d.png !@޿�PNG

   IHDR   d   k   ��'�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  @,IDATx��}x�U��{���5ik�M](�
f`��u�1`p-#�0�(>���Zܪ��-ikܓ��׻��$�$'R
���ܻ��|�e�Z{�͈P����I�Yr�!�L��ʕ(W�����#W�\��N�O�Z)�/���'gu��@���E3�/g5���u�\��kr 0�'?�rx�^��d��h��� <|a0�L�(��p�@�V��I��ɵH.O��`�)a	r���r=%�Tՠ�/�1"c��E##��Մ�6/���p�p+j�ڵNYL
G�ɅÄǧ�19�&0�A��&�a����a����-(�<~A�q��KЈ�&�ש��)�"�n�k�4j�ۇ�.=>W���QY���htz�?�I��&�|~��_��(�G���N��b �h5��9��)�1mD"LF��ćvyfim���ޒf���������XMS�ˡq�3�/)����r�\�*����S�+��X��0�Y��5U0x[�3}��sq�4?����n����͸��X�������B��'��W����X���
�yz�W6�L����k�AJ� �<%w_<w_4�_ٍW�*B�h0�<-�%C�wR��C ���ڍ 2��m6^�i".����^��{K�bXT>���"mx;�f��_$��cBIS^z#��=��?	+�:���n<��~�_z�
ۣ.
ꠀW*55]%���٨�+o����J~���uJ1�s?�c]R����>�:z҃���'�t$�"�,)�叮B�o����\'�,>�(ĵ{��l�c���x��8w�$��$�T��˧����/�J�ur=M��hȠ���Ad|z߱���w,GL�:�nL)��^x�F�A���Q�|m�cLj3Ƨ5���O�Z�/7����'!9֊;���!"�pǍIBe�E�������u20
��� �,�23/	�*�Q�;ar*vj¸�qX�����h�g o1:}\
�����*PT�T��5!�E�ԉ�3a ����)�ᚶnHQ�BX�۱���a���-طk5.U���v�Π�@����b��&�axR1]���w����X����lO�o���Z(�o��NѝަUa��&5�t�D�Ί�Iw-���U�9�Vt�.�I� P#���"10���Ңݸa�n���?�ׅ/����6Sw�H{I1V�:%��s'R	�����v�y�0,�� 9�Q����� �%���&7Vn���s3P����"˗l�����c���5����2T
�qB&�XQ�;����������g��EJv,Ι����V��n~ag���Qp7���2N�w-̵�d�%� C(LZ�W�\�rE��9�<�'ϣ,~\6�V	���6|��<�K�(�I�� ���l)��+�Ć���`\8;��3��YY�h60l�~L���޺���+_�����(g���?�h�&��A��0��޹�y6�_7�v�b{~C7�B1���js��Z�j?^�z� i�:l=Р�#�#�yr6v7�M؞���	�� ����5hh�`Bn�}'���1d`4�6�+�7)��&(cd�<?of:�SAk1D|����5VƲ�^���L
qr���X��߯pF��M��]��2<s���F�I2�ۥw��8�X�st�G�������H��t�@��׸���h�#"��Ӻ^qF������iQ�<���T�E#-�������g~�f��"2�v����X�a-�ޚ�G���O������V�6	2R0iH<|k?�c�ͭ�y�(�U�WPު�9F���'"��	w�ɉÁ��ʌ��J�7� ����]"�b5Rę�~���2��+]�����kd,�NAF����o��f�VR,L�>�}i.P-5�Q����h�_��[˙���;��3�����r4
��V�|����C̵�T'�xW�ucJ��ґ���5�ަ:��b���::��[gr���Wֶ��J��%�K�|��x����Ṙ:*	��i
��|,���ߌU��T�.:�W���~Sd�x��{Y)bE}��0~*���)���eAZ�C�@� w� lʰ�!!�j�%ǧE�{faB�b��DF� ��+%=v�Oq��m�(����p��Pik6�aY��5��r��>3n�}aǐ,��V7R�®�K�*p3az��<'0����N�MĲ�%s��3%��r���kb�s�+N6*�V錚/@V�M�3<Ov����BjT+�Ai��V�o�����ɭ���~l*�"�g`��n�Z>���{��u� f���A���(�� ���@9������w�^(�F X!zⶳ�*�����Z_�1y�H��`����t����//C�|C늈��[+mN����x�b�ڽ�bU�?���-5�1<�U5�L���j�� �(k����kؘ��q�v�18�MB����"�O\N l	c����0(9� hf�az�2����T1m���'�BaE7?�U��g�r7"�{��x�N�-{�������ׅr��x�K�����f�)��b���E�,Q�B0:@��xWt��4?qB+�(uTX�Wq���;� MY��v5i��!�p��	�N��mA��'����\YV�Ή"F�XY�����w�e���Ս����`y��q�=�clRř[`���x���(0�zS	~����G/c�I��#�E����F�0���ߒ%�垐,w�a��/��Y��D����-�q�?��8+j]�dw��;�5CM��t`�!"j�vP|�=SH��#)�6ť;���⛕i�"��c\��m���N1�<��{��#w Nė|��?�T�i�.T�W���*�[.����hn�lZ~�g�J�c+ӣ[�ǻEʎ�4LI)�Ry��a��y�P�"2ۈD#5!�P:�fA�X��:�a߆8{ݞ��i��Ny�}e��[��Uf.}>l>��T=�_�"��V��FWKh�� 0���}(��X�D���T�^��h�na�^�=�7����,�d���hG�5��i�g*���+Dt�
�\0k������D��b� ��j�ɽ��bݾz��z�6ؖ��4 J����Nr��@w1��s�_��1��+�q�%�/�}��B����<��3V�T�i<J�2f���ms�zmrz�e0X��HE�S6:DA;���}��������0��fS�[]>����f�$;���P��T��=��>�?0�j���b�փM��-�4vy|H���"E��/�)��;���@�8���M�����EQe>�P�,2�����,aݒ�.���w��C,:D�$�2/����p��\l��L�E��P
�Qs�>X4�PYV9k7��G�����RV��3B:�u�c��5�D�p8A�#�N�,	a��.��v�fV�6(�`$� jvN�	��@� �؜��8$���i�Ŧ*��&:ɍ��V���嶟Ś���qI���82#/�u�D�	����Q�|��8��4ԉ���8�a�H���>��U�2�8�V�I�7MƵ-5�t����b.X
ge�2#�	��9a�_�=��GN���L��W���y���������v��DjX��>�奙�����.g��������^��d�c�3v{+
}��|�w�H�/\r� �KA�gߊ��c������q�xJ,���%#J�}������&��w�����*D�o�8�[6b��g2����as8�R������i��LIoP2X�q�����,��|K/��`�������3�ѯ���09X�`M��a�E�"԰d{5.���{�MǱu:�W�{ͯ>��[SmxL���,����e�����$�*A�,RB�ۄ��l|*x}:�oK@���6T���j�/�dk�z]�Å����	"R�ډ��fF�H���q�͢�L�Z`�,�y����Ux뮩X*~J��4�5r�������т�K��{�U1kYi�UQ��Uc��'�}NEgk��O� }2N��|W+xˠ6T���g+����;]4�����g�/�y�[[���-�j�T��g����X ��=q#\6��U��&�VM�!��i��v��������=e�+V�h�v�A�3(S�#��JE�F��v��u�媰	���D^]R�*1�9IDǒ�L�)+v֪q�~QU�E���Ӧ���ee(�w�BOS��W���+F�1,�ߏӆ�+��c���9�`	����(0���p:m�7�~?A�d�~CZ�i#���%q4N�����'L��C_)��vk�r�Yp��o����%��ʯ���x���j�E�ŭl�%��v�t��R���49��iV�b~��q~�"�A���9�AqE�w�%�ފ2ݪO\D�f=i񩠡U�нF~�%b�����bU�;�K;ߕ�M��y�2���~C�PN�?�����<(c�y��ojP!w!�!�O��/c���Ĉ�A��j#L����n�9M`����C}J���Qx��I
�+�U�i�.4K���m��N���i�Փ�+= ����˥��uq�U�=I6m@��<�c��[?��-xi�<u�L��9�(ُ)�HDa�H�bOu��u��hT汊��;�.i�}�)���3q��n�f$�=D�C`��j������&��ńW����l.�!IC/n�`;}d,&\�L�_Hs�I�������7�]Q���'��Uf\9n�aA5��B�s#��@d�Gc�����U'aN^<�ݺ�6���c��S�5� �-T�%U�g}|ξ���F�_8��d��e.�C[U V�1F8bL�Jt׵Y�ʎ��3�<p�0�����{�����R\i7�[&���<�� LOޅ陵����k�[���8�Xrh �|���阔#2r5�6FV�}�cSp��#t_[R�bXz�[5���S��)Y����Squ-M)�Ǆ`4�7g]��1mʘc�X�z�8䤞��KAN�6�˩@J�[¯���t�fEY*��������e��'�(Gߑ��EN�0���['�c��o��mۋ�R�k@��*x*��V6%�͒��f���ss��`�ܼ�b�~/d�R�����!��]�2<��I^���TM����i�C�xNsb�s*t 'ʻt�I�Vq�&�MeXƓ�dS���e-J�G�P��ĊB�׬�wת1-�m2�=�S,x^[�O���!5�MC��׶�p�)վLL�0
��!bˏyX��+{ԥ=f򃥛*1�����a��#��FcŮzQ�ub�����C�݂�yq�2/I�b�Pp;n�����
�����`=����O��jw��� �
�\4'C9S�G&�)Z:w��8�^-N"�u���[u���*y�S�"��E#���O��n�5 ��&����ԄSm���awM�BJ� r֝��Wҧߟ?������U�U4)��D�1$��H1L�{H�F�Ko�M���&g����.eipR�gb2^:7IB���9�V)v�F��o��Q3�*��|�:#�}����^弱����=z��c����/ŋ��ɖ�F?>���Up�Zw?������	����q���@�d��'����veIA62'n��맡�9V3�E.���B��8^�R:��NNBZ� 5���:�g6oya��(�նk��>���\�i:_⼼!��_+`3�c��-�0
��|�"�;0��|濼[�1n>k�d�(�%�jT�Ŭ�:|���~Y�B*'N� ���т<f��wa ��ԦR�2����e�|jZ%��EO�4��12����J|ɰ�٨�u�����Ra�Kc��?I��di�k0�Ҡ�S�sR�ԽA�/�>���#�gH������~��#E<���G(�D�b�3�Ŝ/'�0�H'�\��g��y$"�<o8JE����L7��]���Н�4��}�N��w� W	0�	��{e��ћ�"��h�}�Rt�@��9���n����]M"�`�a|���ˈ��w�^���|O:w�XD�{�"�Vl���xkiIϢT�g{� �1� ��н�g"��}KU���z�I0Gi�wCH���t��w������{Ag"�=��.tNSm��QC@�81j�栃k�4Y�Z����g�e}-1���	8w�~0v� J����8Ԑ�ч��;�r%�3�%�Z��#!�c�Yos) qz�I(�4� �!rL��틀(͏0�n=W�(��!^D�	�-br����*g�HQr���w��	J�F��%R��`���4�q6ţ�����)�NᒽuI*k����@KB�H����B�4���+�sa�Rd݊|Bz9~9v�j� �/k��I�Q����a
Ddl@��;�.�q�t�\�X'~ϯ�oB�Ƃ����cV�n��],T;�WC� �ʡڌ�����)��8kX>�-��;��a%}��`^;'N�-�W���A��)��W�&�,|^��FC�6��B�K�N�}^���1�E�#�
��nŊ��j���"u���[��5[��%��Ţ�	΢~�N,���ra���K4������k� ��py� mF��s�2�ζ�QY6޵�W�,�5���-]3�����J���H�E� ��������������!~���5!r��J]]�T��ݑ,���% -<a�������S�2�Ղ��(�&-�_��Q��i���N������V���o}krC?���߇��t䍞.v�R�B��� ��-1�>VG"�T����,�� �m݀��DD-Ţ�� v&��		�G���.u�'$�]]�(XGBb�j��F�5V�D�5�}�=z��:�D������bq}~p�BL���_���Ѹ��w���α*8���ZG4�< �JtL� �X��-�a5���[��Q�N0��"�z��24��)���-
t�PeB��K����h-)�B����bD��qt�0�scp#�@��L&����>��X,�wJ��0&���1�Zh�s>(�E�tR�|D���U�����[Q3��{�ibޑY�fT!m�I��k���z-
�&y�sդ老v'�V-�m�F:��2Sl���"�~�����h�fy!'�
E��S^/���<��z��U��Lx:�F�����^�CHf�1~��8(ط���>FX��_�!l̯�Ek�GpxL8fP6o1�[���hiEƠQ�j�)8��k��P�(�ȉk~ZR�������G���\B�בc��ގ���#�I���%*]iޠR�[ѕi��
�4q���̌���($���^���1�÷�UI�������6�]:5ʕ�w#j�/109
QV�����a�=�N]��EC�	A.!w�$�z*���ǟ���Q�q�lBc���_���/�nJ�5C��6e�x۰l��~���
������>"ܹ�Q������euq�H�ܸF�Z"���ǃG>�-�š3m�A��>�߿�o�vv2�0�b��e9���HM�M<��"�m�{�)��ޣ+�5(/~Db-���������!"�s��Z;�AS�,��"��z�,\޼�7!�2�[�cbؽ!��,��Ɍ���(ϯ�(��[�m��e׏���[cЧq�& =�����|Fk7��Wx���I�qF2S���*�`�A�x&�Vע��U�%9B��J�Ý2�󦈱ҢRTX��}0�����ˏ��8�c���z�]G�_��oޒ��������|rHUU�2���M.��ֽ�ٍ�VH������$[��n�᦯Q����㣆�*2LK��)߸s1�^ђ��v�F;�a��Y�GE)��u)���zx��1S��^lز�Z�,9��v�,M�Y��ϑ{"
�l���bRL�h�8���n\M�O����zhل�(�?B�/�n7!Ş��Á^r�;ˏ���ײ�Mj9�����X��]�N%)��)�k���	�G�/�S�Z"�'�6���1b#-(2h���z2�ȟN�?������
_������+�}��8#:MZ���>3?��C�\�KbBZR/DQCmX$���h���Խ�.R�z�H�נЕ�q�X���:��"����"���?�����/������jF�`R!��*�m��Ĩ2���/&��K"����3��]�3��|H�/D�
p��ࡵS��zZb�_*�x�+�y����ţ�2�
��zT6{ÖH�P���4b^Z	^ܞ�;�����d�{����fNr۷��c�3"a�z�/-ơ�(4���_Mwaܨ�B��r��Jb1�ъk�9��6-͵x��*��3���˄#:	��%x�'L�L,��TL]�6��s�����e�
/Au{=2���nǏR|�vL���gꜶ0 �>���BJ�5�eh�yPZ\����g���=��1TH��޺��ك�.ܬ�3C���ЂSO�'�n�G֋�OAt|f���#����O��G�/��R�4o<b���a�4�o��͊_?�Q��Y��8��Z���9vf�OK�K�-���nEGG��oo>	ﷵ����[�8�^�9� ��梮��7���tĥ���BO����^[ڑ���v��c0�Y"��8��邯�~�oI�,�)�$"����,�h� �{�S���&0^�k���o��'&(���.7S����@��-T!�8�S��K3Ut5�;����'2��O	�ꉘ�
����D�D(MB	�x�P�����n^7פ����f��b�Q,+�{#ڜ�(/�-�;\�ʑ��Mr�8c5���b��*DKk�+��ʉ�s�В"4��\6�-O�� #���}�����BHB|<�R�GY��$�P�ߵ���ߚ�Z��v���hm��v���l��~ǐ�`}m)��ۥV�z�cB�h顭(V3ߎ��������9S7+l�GvЭ(?2�P��G���}
��Ş,9-0��1���U���B}MqDKR��@L��aN= �Y[��S�ҳ�)��$�v_ͩ����󈃃�`"�ߣi=��tG�o�=��Q��6S� ��o�O� �h0�0AE��x[)���r5�i4#'�k�Ue�MT�,��O󗢧���bbR�M��aJw�Ġt��uK�C'�#���ҢB'V�}*�#��)2�}��xc行�I,DFQS�z���zw�����U��T*5IՏI��T��K;�u>�)*�|�'6N���)H"B���?�c�1``�R�aE���ͱ�;�sJ���*�����.M�KZ�Qq���^���`QuGx�}����&�^������O���&��W������~_�2�fʋ��˒W�a�B�詇є��� a�͂Q�f�ȹyZT�� �T6(�Y��6nS�*���42QK�;А����bZ0P�jg7�(�?<�AY{��c��H;J�q���<���*?j���Շ�c�Ze���]K� s����x�/.��%�f��Kq��hv[���c�l�a��*+dq�P|.�#��L������&�?� ߊ��Q��]�p��(�`�d��e�6�=������C� �ٌߕea���[([�"r�ӃC�" r��1m�&�w7]�W!y���g���7�hl7�5Ӵwh�ɽoe`yq��(~��6"��wh�U�k�{؎@�CJg*i7%�.ן�"��TȝTn���Q�J�h���{��:� q��d� ��\���Q'�D3�@�B-ZjR�w�,O�;�""��LD09����f.�L�|n'�����a����*N�*@^r��z�ݡ�7�v�:���=�Q��-r#�&�j�����8�p�����&nw#jy������]+	1E�~=3>��n��JW���'u1b~�bf�hw�
&{1M1��s���/�|-�+��f$,��{`�s�_�FbJ*���jvr����l�SRƊ��1��ڃ��/���l��zT���FN\S��h�A�h#��\b��ߤV:ir��d;�4��B!1����e��i9�V���@�ͧ%��M���ŴcB�Aw����(i��A��񱚃0�۹O�GL�8�%/�V�4`' D�;���f�%f�E�>�J03� �V'���,��v{hᛗ�ރ'�DS{H��|�)��S7�K�*��9��8����T\�����y�LO��6deg㷿�-<�6������mR�	^;%�D�OK/�qU��yj�{��o�L��91qI�-Mu��R���L{�t8[PY�O5�i����xv�d�GH���$���뀞�l:8�A�����¤�h����iڰ�2�(��xH�-ڠ��b�!1u(��hT��PWU�kMǻ5m�7�p�1�O�Q�o4��������C��E�%b����x�o���1�B�Z�O����؋�y����P���B�ǐK��^��I����b��󺅦U�� d�O���g�x�����X��������o�Ag�[wtt�#'r��ǔX�Y��A6p�)�M�z=���?�a�O��6��n"���������?r��	5��n�kz�{耔29�$�������X�2�U��5�-k��JC��A����kV�z��SʿAͩ�וFdqe�����YtoI[��h�;�EV#*&	��6X�s��f&XQ�����*dE7�mCq�:凸��҄��E��SfΏ�
W���'�>��q�Vӫ~��ۄ�U��{�^*���N���ڄ�A7��o��:'�4��7G[�4G�{����Sƺ�����b�f�%bb�
j
�@c�\�����-��M�q���K���Y9��Ch�r��/���;j�7�υ��P_�O��xL6")-m�T7$4 �Z�sғ-h�9�8����a)+0�:Wmq=��������?�= �n�;`U��,4 �>�-H;�f1�jlc@��C���]���rV��cb�pS7F��~@����4��N"x���L�T�ۿ^�XŖ���1���t$�1�׌����Ȥz�-��[�D�1Z������-%��ϣ�O�;�>S\�6r<R��������v7�26��͊��|^� :N�#$օ�S�N�G�m<CE͑w�s�뵠��#f1ꩅ\ʬ6dva��vEV��޻t��p><0\m��Q�>��St�3���{�b���;���V~0+�#FD��"�h�w��7��Sp��&�������+ۻv����S��F:��/]^���d�f�8��C�!*I���)��j$�,�g��)\�8$#מ:���Mn�����M<�{��,���Y�ڡ2óc��*�8����z멞�Q#D�����ČA�UL���ؔ<�y2vRĎَ�W[��sG�:i��V7*	q���ϑ���O�5H��iSU�{@�Cx֤j��YyIj����!��(�!a�����FLN�R�3Hw���e�(��}K�ԫg����Sa;s�1�t1�59���;'
z��бъۧ6^�W"�Ǉ�N������/����V�YK��_�.)�����!$xn�Q�78&�+��f�R�9,���7�`B�������O�Wb���=vZ��@/4�c�X�n���Jm����F�f�B��f�'�r�����p_E�՛��p��M�2{l��a�rj���z.��3s�C���ɪ�m�����!2N���6�)t���N>*�\�"b�AzLK�L�B����+�n<3W�u�Qq��������SGձN����"��#�)Xw���6��/�Q׽޻}/�9Υk˱tk5�Ң�YUg�������<{Ċ��ĕ�j"Y�������3{��C��'�<�r��&� nC����]cpy�n�q$m�oJ3�uQN�y, ���m�BCu�:ԋ��V�����+��Xr�<��~�y��|����R ~A��qQf��^>N�L�]���ύ����b@ps��{&x<R�{�p�ȿ^�ױw}K������	����j���\�����r��.��~q�=�o�HW٪9�av�pهk+���UnQ������d|��'�LǬ1ɸ��mXɃ�l�^��Rʂ�F���!ޠ:��Q�JIs��^w�d�s|%�q���B�����|\�}lf�sN��\�?��+�]���c���5W.��J��E�����0�B�Ν�z�k���ʷlT���o����
u��8�'!)ւG�9��zgǡ���Ǌ$��`B�Xbť͚3)��S�\�$�sEL�!z�Q$�ΓF�hD�"M���v}�V_f��1=�>B/5Q*�ɛ�hr���ԣ�Z���M�}z���Ε�~�CT}w��W�7����ғ�J2q�W������g>.�Df�a}<�2{����I��@��Y�ë��e��sDg��; ު�K����/N�R���(eȜ��z��Ȣ�QDD�=�ޫ��5�5����b���u���2Z,����l����'Vֽ�&[N����Xun�W��Ӥ���P�Ex�#ܦ��Wv�XL�>;y�c�x*��{�g<ܲ/!L�[��\&�_87C��CizC�j}R�j���NMS���E|qC��:f�ox������-
�e<b���)l��sE���G��ڃK�f��y���m��`�B��[�n?�x$Ξ��g?)Tʾ׾��I?Ǌx|���"�#���ġ_��X��=T�ŏn�G|D��]T���N�Ν��p��x��Sq�CP"T�/�Gq�YC�Rjq0���EQ��߃�$������@��r(���D��"ܭ9i�"�6���?(P'A���)~~2q >_WчR���S������4uX����^�/�Do�@�H�Z��e�,^_�7�T��E��<=a�B����NIU�{�P��<�e���R�H5)"����Y����0_(��]mDKKs���L���#J� �X�?z'� ⣬hi�a������?�����DP�(S����$��������~�@��ߤ�I�YK���Z.�C��R޵ ��S+g�O���N��~�ډg4!��[����T�Â{��Ok���-�q"J�r�"�����>#�D�F��E󧪾��5��ʞ���|�B��G�Dg]�/+�CB@;y�+7״��Av�]Ln1�mc�O�*�-E���(C��~����l���"����Q+
u�{���� 7��O�'.Өʯ��q�dQL}"�_,�~#<��u��6������>��싳Y��[�QZӮ��#G��'�x8r�E�KBxz��0�D#��s�~����pA@��Fp;si8T�ҸA�/@QS� Fˀ�����kb��}�ܶ�Ym=�����b���!fU�y��S�4�lK�v�@��r/0J*B�)��ͣ�e��ׄa����
�x�(篨Q���u+r��6F&�)���-��_��v�E����[,�ʷ��*�����P�(@/���~�6�60����^�ݯ�)�޶���sfl��N��6�v�����jp�9G��sH��|�۪Vf�6�iS˽��G��b�:v��}�6�B$��:n�ʵxm�n�����.�C�=ԃ��L�����m�iC�d\2j�hp�f��M������a�2�����f�?���3K��4ɹ��&pzj{BZ%��_�[\�Ib���r�}EI����6A�z��{bj�Jb��b ��72����"��O��~ä-�\���6�czz������d���c?Z�F�S��u���~�V��c����K��u�FEٌ�n�J���<����#�f�B����ee�ϡ��{��u��]�¶�:�ߌۡ2J$M�e��:�$>+�)j=y~˔M,���6뛛U�ʉ;g�X�����r"�sI��O:����g����<���Hs���^�C&�#�H�*�Nۨ�]������R>)�귎\��b5	U]:z�<$��G��������8W�.=4�s���?w�!��o���y�c�ԟ!m��F�n�� ��3� M`�OD�W;}m����<vɽ����������~B�{0a��W!�>%OwK�'	Bn�>%���{FG
35!C���*e_T/֚�t��5�T�X*�D�_���'{,��� �爨 ����Gl�;t.�zΊמ_1�۞�K���>�*VU�!L��ѐ���m�guWp��Ci{-O��+�����Y���|�B��J����춾ku�������ᜍ����$��H�]3w�y�/?^[��H�f�����!A�q�)a!0�������&�N~k&�|��仯�/ф�煹�%���Y%�1��A��E->-u���kֈh�r�\��(g� z�P�MQ�lQ|U�����r�������5?��:����e�S�<l4�Α�CB&�"mO�:� V�&��Ƞ��,h��Q���'I��
-�ϣ6xOo{M^r��EnӰI��Q�T�NA������b�>�/��w����-��˙P���"�~-u$r��W7 ���*���;O�)�뢯��]��F��}aK7�ۻr�*"�c�nB�{���AKח���3&����>�c��R�R��(���1��`���� ��(��~�w�y#́����uD�C�UF��x�ԯ����7<�1�ʊ�ߤ�[J9q��y�x�Ad��{�u����:J�N�����"zy�/�"u4ʳD������
-H��DA��w=�gޤD�j[�#���?&BVʵU�I�'/^}�x���D�j���|H��V@�w�B��� ���P6�zQ�K�Y������5��R�(�Rw4;����U�G�E�>A��iE<\���pkt�(����]��������JW��w�>��]zV&�(��`��mA?/D_�-��!�~��?��$�k��C�]�t5�qs
��sF���W���pM�R�*�f��-aܥl�k�=��&�Zm~����i�-l)Jl�T�������S���P�i֠�;������C�jB7Ei�s���%�g </r�"Aj���CYḵ6��Q��-4+E��#ʒ�i�;�v�5�-Z\0L|��x���ɀy.���DEH�7���b���ɑw�K��u�3�O�.�{��/��~G}�6�V��ľ��� ����R��H�l�&��A?�c��lHraP-�RNݵ�"��3��v֦X��_ڞI�˻�q濠[Y,��u�\���)��~�Z1M�Z��]�?ΑA쟓Q�+�x��TNN*� J#+D�Δ��Vg�NqX<0ܟ�*��.m���P�a[��մ���eb�Ӵc�*}����o���6�y'3xP�g<�',� �Ѵ�ju^*�����a��4�� �|)��값�7�Bn����e3{�W:���S���Xi)�bQC�1�߄a��4:����e�B`v07�q��lD�#l���Y�A��A�zd˔7��+�����q�#���c�>NR�<T�J��#��$�.�6�o���3,r�~i�X��a��������!R�5�S�s�����7;�M#�޿�(-�:S���ů�h���P�����ē��'`�I�J4���slc�c)0 ,��6���<i!/�o�*nTC؆|��a��@H@-�1|'�*�SA���CV��X�*H�\b���o�r�U<��uݡ�)�?�~�J//:(�����ceFJ=�.޲A��)N#E
�Kf�(DUQ$}.�]�éi���,C�r��$�Ŵ���:y���U�}�vL��_'�<&�	-�cD�	�u,����B��>Bt ��=���9I�g�Ū[�40��1令��0�.��'?́O΂�����k��5�Ha<������AWĽŃ�Lu�XFy�@(U!���"V�������Z�� �E�~���j���։��~Ӻ�9�~���C,�H߶I;���)�ȩ�Ү=�[�	�V!����HHܾ*���a��A\h�����z�'�t��m�����r��{��ۃ�J_����oXb�7�|�q#^G�6�M�L�H������޹'q���&g<�A��Co� ���M���1~�rTߪ�Qmo��3:6u~ ��"�%<��#�h��ﲬ�[3�L���ťP��$�g�	��ſ��&�̾0d�t?zU^�wr
Y��^�k�\��5K.n����#8q�U�o� W�\4�>�w��H�`�����:p�    IEND�B`�PK   t~�X�u�̔� � /   images/266cef04-a032-4603-9423-684d401d8b46.pngL�T��րҍ�E��n$�[��Cww��tJ�twwwww��r����w-��{ff����=$'#����B�Q ��@ xYDx���p�_��BJ����5��J\�"m}��j���|����������7����wS[=�o�6F�G�� 9HB䣒c�����O�;������XBX�^#<ԒH�H3<3SM䀹��ћ�ԛ~�Á��}�$�u�D�m���r��5�K���VmO�M
я�D�c�aJAs�w�;c��H���Q��_�xR���������"?�P<a�nn�CƗ7�`�}�
L@�Z`(uԖW�΂� c��a��>8�h��PA��塤�<�WǬ��|��&����l�MU�3��B�@e
ݫ��U<
�K$�3��g��_��R��=�`�b�hQ��m�������� ���G"�[�g�KY|?��K�٫`�R �Bi�1���E"F��͢�N��e�c�S�c��`�7`�S�}ي�a�D�^�K;��;�w�>/�r9�#0yuX�7�&�9ф�5�زE Lz�ɮ�Y�ZP���qл�;0i>{j"�<���`����tY�>N�\�Ƭ�F>� b�юh�k�F�I��$���߲��T%�����n��\H4�ō#�,s�{[>�q,C�'H4c3�q*(���剫p���s?�����a-0�Q��گ~���QX*�@d�Y�����Hu�������SBn�_�[�B�!���֩87�Ӡ�v��j2�YŃ�@��8��{�¤*ay�8�^��3�%+�A6�"�B���e�*�c�L��r��Nv|��
�-HT���;������`Vr���oL�C��D�[�9|���I��G���˅6D��h؎ψ�>�!o�ݘ3$4q��!izP�梉"�%}M�6�EW��ϰQ�3�2�Wtދ'4M	j��1n��z!](~���`��@�{����C%�2�_�v|[��@B~&MW}���$��ܠ	*��E?�V`��pnh�q}�'����Q�z�ݣ���i�j��Q���M����4�l��Ռ�&rȶW��$ԨK~����w�(�r�m�?ϭ�j����N��v�4��W��7A
�3�M4x��~���G�ĿPńst,:~��kE���y�㙭�]�zf8���S�"�l�ċ:��fKH7k��_]������o�ĮJL_n��I^�UvQg��@��I�F�WQ=�-���K����ۀm<�|��ם\d�����;�5��/γ��@w� ��u�-����G�H�p-��K�8BG�oc|��U�+�%�����X�Ӥ�X^>r���!?aD:{�C���������1��>��4֔���K[��}��Ji����?����e+KK�ՒrwQ��{���G_g\�*PǑs��KM�+Kڟ�p�v�=b�Zt���-��Vjf�wc�j/լ�!��3Yw�=�1��__�<_��Fx����i���z������57D��0���2f���)t�vG�:0�-0��:�BȂ	{����B \�����&4��]���&+q�n&>����{LgSt)u=�����8� ���5#�
���	����yEk[.l��]��b�W�ȁЁ�$���L��H�t��B"�d�!T䣥�����CKPF��,s��%�g���DX��ȬA��<�ь]3��H�����"'Zh�<��'A!���񍁺?�#	4�g@?�3���:%�		�Bc�Ʒ��'E!�����6Cmcd��el7;�b��y�]��y�����eBөY8�J�� !���[�S6T	���Y����z�I��L��'?�x��Yg�d�Þ�x�&��T��ڠQA � 	�|F'�*F�FzҐ�6�'(\�����_� o=�z�zcx~�i�:!7mbe�5������Gn�X���T�]�G)~p��%BKw�|D���'��@��To>�S~��Y��Ā��	D��j��!� ~��15�R]<
���Q>�}���]nnEFƔw_]쳖���ʗ�Ѕ1��D��w�,�Z0��*�\X)S^`�½�A�#���[>m�,���D�Ki{�/�7ҋi��_�B𔦾x<�!�7��T�
�ȧ��o�V���Ǥջ>���&	cd��9��
�9F�5�x �a�w�����/�h�}��l�ɾ��l'*u����7���H�O���\�����$�5H���)M��x +�=��K<����}R疠���kÍ����ǿ��:�
�~ds#��/�=}��%�:�9YO��$������	��-0`����xߑ˝���̮�DH�SО���n 8��s8����X&�֕�"y�"��������D�lsV�Hd'�OM�9�g٨K*s�EA�bh!��7�I�ث��f,�� �+L�S�7w��c�o?��][]H }t�A�{@��o~��!\A� 3�giA�=��Dh&�&�<?�7�D�q�1��ۡ}:����F�X����]2��8��V[9���U9cW�*��H�ۤM
U�´�a��-�B��i�th��G�[:MLC�*��G;�`�����8�6QK_V��8�ch�M����]�#�?�q�K� ^lc�0�������j��<��h����ʌS-�H�@��K�ۄ�Pa�5��%���@]"�g�x�^5>	��ʓt��%�q2�c�;�(�����m��M5N�R����wt	���
�EK�W��MvB�~x3竾�F��I��!&���![`Y��ebƩ��@[�*�v@���X�4��Sn�Q��!'�_�#?|-Da��J��
5���1c�hE�8F2?�t��C�̗PK���.3�'�+���EDw,R�3	^D���d������/�������!�׉��S�Z�L�ըۺH�n�<�'P�9Ņr�ݙ��L��J���y�d�qt@X8�⍫!������Ð�"9���w�,E1��r+⪲��/.�lS��t���"�(�!@>*f�Ջ�ڸN���̸��-4
)��-��SKQ���\��÷j�ˇ��C%���{�F��;Q��@���8!���{�vht�Sd�"S[��e�~1�����PtVj�+N9+��B�T^�ӟNϝ"�`�����Y��CQ�|�~�s�v��nI-� �Z�#n)����`�15��`,��V	�wD���Ry����/{�����Ȏ���:䍥���]a��8C��/����EAWD��KL���ֲx��P��%�9&.r�F����7�n�9�����<�`���E���T.Z �5`O-��$�m���e+��?�*n����08to7:�}n(T��ͷ�H�(<�A����Lj�D��s)>Gxˬ������{�oqYN�����˗Q;���D�2m��H�F�����qj�9(d�|~o�G� ���Y6M�_�pBg�N�s���a
W����פ�h�Z��j��D��2�;�p���I�;-��D��NG�+��C@��P��<�� ���9T6uee��8�+�і�(��7y�9�Hb*C��lI|�2O�����,�w�@�_Fŗ�z�5i��?T�F������09zkN�?���k*w.%c
d��=��m��i$Ք���z��O�m�)8?�s�`;��[7���/j��E^^~TfdT1�Z'{u2��{�W,O�M�$�����g�|)O�]��\�#��J~�x��7��T��ţ���I�R2+JN��!;���G�~߯1��O�}��ķ~�Y��2D� %��h6���2���|G��y���z�hN��?@fg�)�!M�k�`���v����}Ɍ�����4Ki���G�Spq�q ��M\���O�U�n���۾)^?[՘�� ��]�2ۦ˘^�H@{(�tb
 �^aa�EJ"�b�RЭqw�yg����?.z���RGa G[��a��6�h�̠��s�%d��Tdɳ'l�]�|��{���L��[� �dp�DrL�}k%��o�|w�{�ȧ��͢)�`���c�i0X��W�1>�t���L��ɝ�9��c�-�0w��u���٣kЯ�9�N�p_!�:.h?��X��ܖΪ;�u{����bE,c?�H��G�7��>�X�[��M�PD�SjJdV����>h.�(��}~�+�aν;w��$��i��%���a�:ld_�̸jݧ2�dam���\���(�А�T2дoIa�����.��S~�� ��:�shz�w��>�E�0Z
Y|���"��h�X�2m����ǰ�|�T��J��P�pTA�ς�%eP��b6f #���6��^�b�^	C/����&n镾s��SںL[״=NE�*��,���0��'M`��N�R^�qa�}�1p�E��-M����;����S�|1Ck�>��8!8�";j$3�ؓ
Qzw�w�����G�\_���,v��
/k�V�>���%�Q�!�c9���i�@5���I ��t��na�4��2��X����rh��o�o��}r�N6r�N:����Ffi�nF��Q>,�n�_ b�u6-p济
� �+��La!� ���E����Y�������T$�&�5�B��v���O��j�V	BJ~'ˑt5at�*2�;�] �e��/-�}߯�w�r�����MS� #����_�����3�i�����.��nB8����qm��g����40D�Q��Қ%q�!H� 0}}�i�x�/웇���mZp�T#o�1vi�;�g�5�񲃧����)��7���̬5��0C�Y/��ة]�s�@!+�-��5e1y�3��9�$�
��[EhA�N5�R�D4e���W1g=#�n^���a�G5R08�(h�+)d�w/$�u�!�9�V&��[��{��h��ϡ���?�ߥY^��?�c�+ +d��-�,j�pQ����8�����'K��RBq�k;m�����|Kt��4%�zX�׹hk��K�TDoX]Q� 81(Ψ���]�v�"�x����ą�Kw�^���e ]��k��@Z��[ik��^6<��p=�~0����7��F�{�o]t����g&U$��/\T���S+�p�����I ,QB����}y#zz27����K���.��u���=7�9
���Ԭ�C���
A+<F�C�3z��Gn��!	��G��\e=��Q,!�g�c�wq⮫0��-y�8�jA�:^�$Mgr����\6
�0Ǉ`�7�W���Y�ԉ_6���������v���'�z"È�	�Bh��Gi�t Y�Yi���. �����/�8��be�d �Z:H�of	��p-��,H�O�\t�ra'� l0c��m�����O�@�G0K�ֵ�^�3;�B:��X�xb�x�o�=��Oy},Y�/#9�`���]��Y�!*5tx=uD�>�#�t���l�P_��Gu0\��庩�A�j?�U�oW�R�G��w���MB�����3'���@�(��g��`F�A��E-�)����O��+ac��o��ra5�J~}���Ι���H��� �2��ys<��M���Q�ۅΣ�0��C��יXV����7NO��^M}���iu��ʥ�A ��aM~�EB>j�);��`4A}Dk5ޙ|2 Iy�:�o����M�B*֜�0j��B
�s@)��=T�:�r��pAU�ʐǱ���Ͽ�IH8zm�E�s~�C:��4u<X KvxB0��X�*��Z �brv\�K0�}h��^}u9���j�91��p��?�ip��v}�i_�'1͑n[�Dά�������[kw�ExR��9�U��x���O���v_���(�q�_:w߅@_��l(pv�ZW�{�>�"Ɩ!l���Hl_��L掼D�P��xS�V�����p3GB#�Z��e�?@=�H���g�C���\5���3�;�d7H0�h�	�6����}�#�+���RK ��浯�ڛ�Uʀ�7����|��_���x/�U�]I���^x�q��Bk��{pHZ�)_8I5B��[��~�$�3�6$b��_�����*���g�l�@�#W.!�ST���������U�#S�e<��"��|�"vq#�m�[J6AHҳ^�TC�{�wG�-��1�A�I<O&-i��$���F�Z4�#4�X6 -6P��6&ֶT�����J�_1C��{N��<�_�?�O�^�>	�!��X�iT��қ7�ϻߞ�1�頚�qo*�QZ.I�5���3�l����썂KX��዆������B����i ����{1l,�ٳD� ��ѱ����>Z�X�*|*0{���E�:�{���a�e���O�w�������c�F�l ��v^x�#}�i����g�K��Yj�d��r�Z�(;1��g��b4F�x�=���e�[����_��,y����\���H�@�	��E�Ǐ�s^�� �̷�����a�<�q�5i��VWM`��+�߶�\#���|���VKq;-;$j��f�;�01��Jte��aP�z�>�Q�0��GZ;��x�EP47|��LW]�\�����O��ޕ~5�R���e@bn.R+RR<h,E�V>�ɓ���ԣmJS)��U7���[ډŖ$�5���#�|���Px=��J�V�\,�=mqA��O�{Ң�&�m�Ƶ�����t|��)�T[=����xf�4��^
�^�<6�ۣ�� ʹûn$NgB'�Ě 7��l;�Ҽ���G�r�[�.��6��y�	������@%Σ,�����t�Ƙj�j-����������ОB�КB�d��@�)3q����JX��������G�@�_J*��h"��2W)KW`�]~�����՜���G�\t��U��^̃��0�w�Ky�Q8�\�Ŷ��V��<��V1���rqL��� �}�,���'S{��&�8s����)�|#q||Y���0�G@��t��{3��B0ȩ2�>������[I�,Ɠ)�Haed�(�����?����]~��:/��O~\ d�_��u��
z���ҕ��y�"�ga?�� Q�i�xV�C	���?� �ؿ	�ȐRcS.�"��R��S�0�5�fE WS�N�rjc����X��~��^[U�b.t���}	~4_��m\�UM� ���@����OPy���H��ylm���@4��@�ܞ?J����e�Si�(���M&3@^ύ�]����� �|i��,��E������yh�F��j¶ÚZ�:ǡ7N( D�|����5�ڱ�3 ������C�O�1�*,{g6��Ǖ�������v��Ȅ�M��!�ư�,��g��;(:J�({2�S�aN.b�C~����z���k���C�n�A#���.�j�����"@v���{Z��qJ��M�O��i��L)5�B{#�X�T��\ےh4rc�ʫ=�h�Q�VJ쿔��A"@}z<1Tc��Zz�ƾ���ß@V[	}1�ֻ����Y#uOS3�I����vD����ʺr9?n��̴��p���v<a똹�5�d�Ŷ�Q�r���~��4����n8̦<�i�Xh2�)_6��w��k��A�Z��q���3e��%
w�kJ�c�lJ
57��A �\�u�����Q"羺���$�a>N��c�F��ЗiU����j*���h��i �q�j��uZ�����eW~��|U��9�V�-�d�h��=�b{=g�'�e�]��=NY�Z�F�m�\��vƿw�FXʱ�(�G�)�EG\h_�~��T��j��������18ݘ�`SR���stw�?�1���#��'�Ǭ�E&�K�� n@T1g��mM�y�@��F;�������d��:	a��ߪ�2��Ϯ��\:)W_$�����n�ԏ��� V�\�&��y���Uz�Vh�8��C�f�K�
�=�Kn�q߭�&O�λ/�b�Fw��q��������m��T��&��>�updX�oU�GR�,����>��*����BA�Q@A.B�
�����}�EnX�SJ��X�B�n�h��^卾08��
��N,NO��YD���:jF�Ї�ӚS=g����o#�����?'�W��W����d���ME���I����0��%���p���O|��n"c�R�x������3���|[�Qi[Wj���O���}b�fԉC����؞jaCOkM`��Üb�ɸM��<uj�U}z<�{R�
�������:.K�i������[���r���w���X�#���Ϋ�1Ҍ
�_�Rƌ��:O���K����Uѿ���p�+t��s6�q��77<�V%���R/6Q�N�@��G;�)'vw#y���07�by�a��-�7(_�i��J;��0�؛W	F�]�{������n�{�ly��>��u8!��[�'S��l.�����6��K�y~z���JP�zDKEȊp��S_Wi�⽮n�z��W���jf��bA���k]Yb��\� -�MA<
��~8��R���G^�Vw=P�*�M���E��oN��QY�՛3��s��;hmT'L�.�ڝH�F)3^y�f5*d*G����a��Yp�+L ��*gL�o�����!��!���C`��VQ׳A�1�/����V׉�s���#�z��b�<Ʌ�	�w��L|ʚ�1C�����I#j�Qa�[���	T�.��ל�ԗ:D��\̒�G��������I�j���j�Q�L���m^�uҥZ�M�ˬ�Xn����ݩ�B�yA��3sV�c��o�Qb�V�eޙ耣!QI�J9����)/�f-�U<H��Z����E��n�I�g(�"�&iL�GI�XNU�͘x��#+Ҕ�~�G�� ����VY����F�Iӄ ���[��}��&B� ��Ne�J҉��z����&5!g|�*f}j�j��cc���)J8m�Nt�9��~���Mx{]4��1�ͭ3���U�W^7iٷ|(D��NN�����C��\߈��7�Lpi��6CZҧap�%$E��bq7\�;�7ŰT���MT+"j���@�N�R��86{��D���\mL�};�c���s����� aʲ�����k�sֲ�gI��a�EJׂ�$�7���w1�y�79>G/�G!���(2�I�Տ������-��F�ڝ����|U-}��/
ةI�����4����n���w9k~���Z�}�ok/9��v�*�|��4%I�Db+�x�L��D\=ʱT�-2��_��L<����q�����(ս��
�,�sG��Ma<�| �������C�Tw��qeQ�ģ秵O�QY�;9��E5��"y����
����@`㝾�|C@�q�' Af��<���K�j1��q3�k����-տ׷N���% ,[Md�}��;�A��5o��{�lZ!�Z��N���:Q��Sq�����*9�r�Y�$�I�w>����P�y�1ߖ3�g���7"M\[ܓ� � |�0��U~�����2�������ݧ8�u���a�T����1�T�xK�v_62i��>�W��!fynB��w��z�|;�1���T�:.�wB�a��%��6`s��S���o�Mmf�7�tU��4���W���d9��J������薿LAE$����9������yǰKeWWiuH+���;���K�WoH�=�B<H����~�A1g�>}*ү"<Y�W��F�f����a]j�`�a���i���\��B$�qQ�h�P?�����I����gQ��xT��`g�'�DÅ�^W�&۴)�	6��8���t�W4�+��cV�3o⊬��:�,�Mim�'$��ǌ�硍�,�X��2��ޙ�G��f�e��6�Y-P�.��6mM�s0�ś棗B,����3^[PMxj��5��\M ���������!	̷y��/���4�W>~�2�#�Zc7�K�!O�BB����"�W�,��7G�{��5��B���ܼ�����Gܵ��#F��.7K2�~]}�C����=r��M8�?����'%�z��V�����9���ڛ��s�غ+�`	R���?����1���)���QNz���jy�3"�#U����QӒ�^�ze=�/ǜ~�B����Z�*����:�!px5w�`�a�
�]B<\^��o�Ի�k
�]�|�����?�o��;`�[ $�s�[�i2�*���������E\��dN�i�`$#
�n�ʰbҫ����ٍH"2���:,�ְ�����I��h˳��Q�,��`@��bD#��8��aw��!����x,����2��8�_.�~�����]z��>��v:�F�Q�C=\�ݹ�v/L���tM�՗�>�֝L��2:>s���=��<[�m�H��`�*��O�Z��d%�b�F\��̴�ڜ��&ѫЖa�Jg\�w��ѧWv��}�h����(a��V�$2p����7�����[h� �y� s0d�dg��ټN�������V䙾�9®;�d;�vķ%��㕿6Ӟ�x�V�,	���R�T������ò�W�Æq7�m��έ�3$C�Vs@�VQG�1��j�ʹi�������!i�^��?Y�/y?�]}�ǃ��� ܇�9�9����٬��'�I���jdՒ���A.*�~�a7{�zl�MM���ɤ��"���0�W.L�Ii��c�VB2�f7�V��Z}|Fh��w��I~��
��}��B���c)�SH���U�#vv�9YPq�$��\��[ӡ�fIq��ٝ4g�1�T_I���?YnXN��q}���Z>^�F�����0ȐX�&4�RW|�����4�`��+���V�G=���`�J����L{m�@��p7G�px�Y:�|o�MS�V1~�'$���I�,�o]67�mc¿�\M٘��D��D��"�������g]ע\o|�}\�?b�K�8nN�U��7/�#ɚuQT(�����v�:�V5�0˷y�ߝ9{O�OҚ[�iyR:�Pf������]ł�m*�f�@��Z]�%�1~�xd�N���7d�!?��w���-�Vn�*�)&U��<���|t���xNKZ�=�47���@��E�2��jА�L���_��[�bt����/7���/�Nߐ�U\�,�Ϣ$SG4��_���9m�xo[���2V�>�'�NR��L��m��賞�L&�P|ո�|�r&/�$�Y"��B\��Dtu�9�?y����~�#|�����G���t��W�W�K�������.əmoA`�D������Ћ|YuF�<�փ�<��F���"1�})z��ɼ� ٻ:�"�=�1�;�.5�A/���?��;���X���'�O� ���_]���u�`S�2�"�R�/q�����X\��
2~�	��~�$��]J~']r��㔡���5;Qa=���؇�V	�����ƾ,U���:yF�O��_֎E�z= ��U�4��?�;��s�k��꯾�kx�y�-�tf���0T�Z(����U��h�������h ����׳����-�.�ZMx��y�l|�#����V�|]|M���T�/�`��T��v���~m�~v��y	u�ʫ���s_�вS��?]#��E;vSLĻeh���-����	�?Mj+ZM��<����F�,����^�N���y{���ŞG['ƈt��@û�@Hu��7�f�`_1xc���b��\�c���77��v��)$ɪѣ���f���fL*��Q_A�R�SLw� T���֝Dbo�^��e7��ܹ�̱�U��9^�Ї�O���9TV��C�w��v�&��i�9%�;�v�o�M�/9�(�Z$S:���v��U)���I�<Q�k:*��C��Ċha�������* @.�*P�� C
Ha`����P�g�itq�B3��h�R�����(����"��W��b�|���:R�i�>���|����U����a������K􌯭P��[�F+��`ۆG�,���8#Uܜ*g�����ˆ���f,#����&���%��4� �cW�԰n�9�p�K)��D�� ޥ.�X�\�O��J扖��KDrz�er��"�	�Yy�*����G�^�����q��뱕��)a�K�� �%�F �ŏ""n\^ň���4��4`��*�����?�)�M_B��f��K�R���)��ӄD
���]���U�����z#�[��5���o|v�A����>Lx̐���þv]�$	�Q&�@���k����J򝶔u�}cC㥡3�S��]kGrFZ!�V�u�c�]Y!��seg�f�r��j@9�I�N�tc)6���{z��g"� ��uk�ej�_I<۫"Q�S��_�*��Ѯ���|�>{Ѹ4x��
T�w-�)���t2,�T�Z瘚o���(w���f�?�ůNoy��;�t�|���Y���l�qE=5@,���8��1�9K�����HP$�g���!��g1 6��T�C��GJD�[j�"�??x�F$��f�+����0[��1���-��	c��?�$��6ֲ5����rq�1L�L`/,�'����`94W�[�A��|P�4��3��%6��щ�ڕ�_��*Ax9��Nϡ����Kc\w��WKu*�;��>��4�w��?�m��J<�"�u��O��fu��g��?�u��F2�}>v���J���x�W�C+��@���p��X|{T�κ���p"_�����n�c�d6�A#�����������FD �,i�@c~�����Y��3iH�4#��/B���M�+/����*s����䒲�n-J]��I����,�H���X���D��|���Ү���u�O#����(�����ڋ���#	�='j@�@?oL\hRt����n�\������/��Z���V�0OOx�ъ��Fi��~	��̙�Թm:��".hC�?��00|�^j�켺�"b�GP1g��csUY���x~>��5�GD_Ӹla� ْ��6�Ը�L�h�*Lt2��<S�m��v:��tt*���=�ьI�:��eM�{u�3wgS�`!(�D�Y�BJz�"V�Z��S�z��S4�`a�r�>���L8�����:2m[��K�8�a"�&�$W+K�Ϥ��c�V����Za��G'��O$����qǱ��:��Ϸ����q3yj��<-���Z�7���^_s������R~�G�����T�$������	 ����|<;o���̜x�|,��d~M4C�,
�rN_�&��$��=\�0�젊_G���F��\��q2^
H�pV��z)��V�V�/4k����,���e.�^��E9����_�J׈�9H��})���͙V�a�&���(�)��T���1���t�����<�h�Hق�Qn闐��ԕ�ϙ�sL�2Xr�5�t��+$*;ԹЪ����_�q�Yô�CJX�{�e��i�cA/�WC�b�9Ԛ6]����&-��~'���x~����z{��*������a��V�7��,LxE�B؁V���,Z�^3Z7>:����s���Rf��Σ
���,���@ן%:�TZj��oku�#����43n�j��du���]&!�ZƋ;��K�,�
n������:^�D���(��j�����AtN69䑝��i�6����#%m�]W�iH3b���K`v�Q	��j�7�^�Z[}&����;���z� ��-����kZ�mNl�G�Wz�K���|<�����և��I켣Yի���S�v	�)C�6A@��踃���)}8Mzq~�k���E!{�B�U���������W���$(Y�v���P9|��n���i��e�>:�N���,�M� uѩa#8i�5��9�dS�)w��}�sxC��'d��Y���	��~M~�%��}��Ã$|G���T��~����^�/(������s��dQ�r�Uv8\(�`}����)~���t ��pz9�ٍ����]����V���b�B��ә7�ˋ�#<9�:�ݨ�sp�핐)����F�:�DXD=�H�ۋ����i����hk�ߦdUjfh��<���\�+kЃ��=*���&�v��Τ6}�9 �Q�.p�����~m�s�$�r���m\���Z�o�W���L��2/���h!�H�U���`��(��z�����e�,��ר�45���"4n�8"Y)+N�^�F@X�G�Z�;�m�,;M�v�B�h�\B��>n���mٯ�Yo�;2wgd�IL%;dC���w�׉ݎ��6+:�W�:0�}��
����G���%��vCw"q�zIW#���2zw�U�kI*�F6�C5,,�٦5�~=��{9�Np�A��-����V��M#�9X�7K4ʾf��G��vQ
W�I�6,�t�.��"%���M��k�~�j?Y�z��7�>�mI|�9��/L:%�l�߶�|n�k;	^�K�pܪKyɉ�Ż|�V'��^��d�ȍ��2w��Ɏ�7-��(?F�3��)�բ�5֖֬0$T�q����"�qi��p28��ww����b5����n��[s�@�qia���@q����`�z�+��9��dz���`)~������9[Sq�euX[m��k�(�T)-7o��D�h)���xw�W����e�]H_r�A+Yt��=/����8�,��y]l�V��E7��e;�h!݅��ġ�?9�u��N�_n\�Sw\��-QB�YC�0\�;�-.6�MTr�
��^���TTշ_ ,�ڞ\U���3��e֐ײ�$�
�
/WH	��j��!H��2��w)k���',;L�ًV5u�_i	c<�ޭ��ݶ�ΥҊ:X��V\V���@L��|_frЛ�I^;���f7��[�琞�,W�"�w�֛��֚��0�G��y$�uY7�#��_|\���3�?�f�}�ߙD�v� ��Z���2w@���]����iJ�+�m@`����-�G���WP�.z9����Wy�En��mI��"Mmi\VnsPY�S��Q��<s���&b4/����:84�������/¬c*��Tb/������U�y�:�u��
���̣6#Ɉ����R�NԘͼ�~1��n�u�.�!!=�m	'�yNf�I�tf����a��BZ���m1�_�lP���4������zM��W�αO/��#��F���X4=Y�,"#��Kh�w�n��O����s(�t,�w%�}�IUuQ�����F9"�}�<�}!}}�Q�~iݟ>k�:V�=�6cÛ���=�6�v��	 [�x|�w�O}o���4�%��*�t�K[b�����(%)�$m�2�`�+Bk	U��9k�iaw�gm���֮��>i�Q����|9!��VT�C3�m�[�j/�s���eMc�5=��?���=�.��h���Z.�[E%�V��.�g-nv������P�ޜ)gb�c�w5__���U����̈q����?̰�LB?ة���:��ۈa�����Ja0����V
��(#��@ȷ�Y��8�T��ن�[��XU_=΀ti姾�� %)���N��S4�����V=qR���ָ?QP�R,O�J��?��)����4�Z�-�Ӳ|7+h���G#BS�6_�1�}`ǟ5m��K:o��[B�etu�fq�b�_Ϊ��2�!�ۛ�Թ�����?{���q�?)g��+�{ �1����w���K���*q`��,'-�i���RK�ځ),�H@2�lky��i������E��3����I(���~X��v	>C9� �۾{��Ǡ�E���ne�-�.Ϣ�VJ6m������@e�傸� xi+����er�|驒����)g����
��dF���\�:?��U���v�|���Z7{�����/���П���|[h�"\"ꂺq���<:<�򣸔�bwU�R��S9���ɼk�Ĉ� In��Ҩ�g��f��+��Ed��*0��ucYIID����Z�2�l��p�5v�
",��^O.���M�^���r=is�V(O=E�"�TA��{Xۧ��L�"���r�����y���PC��U��B��KJU�VZ���ײǡ e煟֧4�+�O� ������d�Kex��ӷd������Zٜ�b)���X���{H�IW*�iW�����O��%�?k��kv�s���u9�
>�?�9,��+�yj��^�`I �c`%\���~�jL���.�D�X+<�\�fkp0\)��%8������0U����O���###{{���ۓ��s�w��[|���9A��첦���s�����+�.Iy����c�/����=t�X��zҝ�8r�a��c�Y�p���+���)j�f���1W2��'�oxT�{�G����:���uz3Bg,�����n!�,�o�q��.�g�8�q�W��Db$E��$�ݲt��T3�� �s;u�� OFg��f|���pLZ�t`�3Z�����rң[��Hv�h3��,Tv�����]�r���ΐ��Fn!��Gv�vAw����A�J��(�!�{���*�+�hn�`��<t�T{3������u���y�mk��FfW̎��y+v�GW5���G8�~�rt�>�<�q����%#��C��@<��[b�{~��L�w�Vݙm��}�����u�8>NdM�w��$n�R��'Z�%���y����|�c��6h�2��G���Bj�)=Z��mm
\ձ��Fk��:j�P`*=�Ts��aK���rɿ�K���#�3���ŵ�g>~�*cp�G�-'O�K�бo��9.�����4\0�[��h6��:�6
�I�4jl5�ݨ���'���nl�6Ol۶5��w�_�����^�Y3{(t�P�l��e~$��kz9��_$��s;��?o!�i>���)�%���ģ<��*���?OV��jӉ�@��	� +Bt�,d"�r[��[���<6T;{~|��A.s���ʏ�T%.ލ�2�~��^g6~GeD�^ks���/)q>aL�`�	��J�ط���`T��$� ��d��+�2��϶�7/xc���ИSdg0�x�e,���$�)��q�6�1��[P��#F��kS�K���5���Xp�U�����a�ꌩ�%W��1ZT@���C�n�c��Ɓ#����c�� ���;U+�Y�4}��v���7<9/�s>-��#�^�6u��\sז�|�M̸.�{�oA��vT�%�Uqc���FA~-z�֒� :z�AFt��RE����3v�p�gرV!�}�����E��ߍ7�f���G��g[Z6&W�M N?Df<�x��ac���%�-�� q�B�J4�-��B��ag���=�|%L�T��zC`c�)��o����b��^��:g���'?7W!eWܒ%M����Z�sT|��Q���T��E�to\��0{<�,�����_o�5:����D�<��$3��k�(��`�὚̇ M"�8���8)w�#���g��0�#:(c���h6�Y)v��D �s��΢�?��BM�J/]���U�Xp%�HJ�X_��Lw��5�R�?�^�^�E_i;Dmt������[�����g/���'Y ��Qe�n����m�k���U���խ�����z�M��7
S�7��O[�e���ݹ����$j]��hOϻ��]~��OC{V���:ܽ{�ٓWD:nm#K&)9T����0T�%ϊѡ�p4S��I�P�ҳK��Q'���	27M���4_~�ѦPƟZ�j}d�ܸ>��ş�ba�b�����*�c������3�����6_� �J��
�Nj��Lo��$����#�j�m�g��X:S�~l|s��㉐��,���=*�&�d���[�Ǟ���͉����~"l�qB���H�D���(oѫ]M���ͯ��[����B�����嫛�� �_5��LW�S̅s>B�`Ozة&����x����DxP��v'��~;����K����j�p��J��*{E<�s5v)��!QM�r�ה�����5���w��!��΀�e�S��r��,��K:!�ۤ��_�=�<=�474���{dp�|���n���p����-��`���E2<�2�}��Wvd51��ճ�J��L���y�,t|{���E���~���
���R�r*���f��
)��S���U�Jz_̟Pp�����0g;*S�=�}U���5`̳!xP �`����c���rW�b:i�C^i�ɻ�\�{FX?P�D�a`����k+^�\g��qB!��"}�_=}��tA~zG��,壍d�u�}�V�P��+�ʲc�@��]��5Ĕ�ep��V�xV�𔱩G�~�T��tp��&���C�0\�>�$Q�`%lMo���EؽZ�T��,��	<��b��1�IvmQc�Z��V/��'�
_?r�ÿ��V{r��v�l�3���$N@���%�� 84D�����7�l�e��嬛��Pr�u �c�gL@�H�Ղ㉵=d}IQIۢ�V��jΨ9|;^��]"��JA���{
㤪dO��S�h���݂�~����7��,����Z)��5	i����a�
g˿�V�3a��D~k�������9��8���6(���� ��sN3������͢Mp�-@�tP-��f1b��k����U�tS� �]v��DnU���nƔq0`֨}��r #�k:�$%��	$�j�H\6������ߜ-h�fejׂ6_��@M�u��v��s�u�J��5���%�`),顀h�M�t��Z���X)G;��E�:;�N��r�i��"���~���ٕ��R�f��z̦1�.E������b��9qdF+������ �3��k.���V�2EĴ�dA���4���/n(�� (L�Ȝ o>U�h����\�߱X�)��!y��Z>`���\p���}��U��+�D눣�%\�,���-�����:(^*���(QV̣l���	�� n���pm2۽(&���H�y�[I'��:�li�-��wsO�/��ͬ 5�m�^�`.�A�;E�|n�Y<���)�6�Z��$���l�'�����8�z������-y��ma���ˁU�=C�+��!�m����T��H�̵d����bC�'���|u(��t���d�2CNQ�1��	-yq�q�ѥ������4��:��0�(�4ˆ?d���d����*�Ri���	c�1Yz��?�;�ڦ�*����V��h#�,�Lk9�Uw���H���&^ ,��*�F���I�=��w�l��X���$�/I� k�?K�O�;]����ne����������x����x~5!����낻�~e\��ݐ�G��a���&W���Q����M фK4}��B5]��&K�)�Q��9����l�=�8;L���r.����Ǽ���d�p���-�O+*�K�h=� d��1�����m�DCe�d�<����ti18�g���sSl"��O��V��}/�+��`L��ѷ-#��0AW5�̩M��:A�n��O���;X�7I��r�ЎM����)U���pz�ע�>`�ۤ���E��Ʊ�
~�>�)_�cHm}ɜ���i���G�0�w��ǅ!�%��|x�a �L+z�,�!g�ϤP0zJX$5��B��nD��lm��[�i�ǽJ>�+�u�V?]� �ʒ77a|/M���1��(;�zθ#k7�ɤ��+K1i�����T�l���	���Z�ե���R�p�C�E�-at%锈��y;���y�	��'��(z�D�`h��/�#us��Z7�}���j�5�Tn������:+�~}�d�뜽'�˥U�]��GR?��mu�b�p*��@Ud���G�#�gt���P�y��5=}?֒�*�Jʄ��r���aQO�����m���UE���ޮ����j4s5mO�N���g�����`)�H�Ui����)�#�D�����h�>���(�,�_���DR6b���s��e?�؇�&��v��ݟVql��HRC���VG'��c5��b�ی����<Qк�K�����U2��2Hz�|"��F�M
���]��	�Nu�&���x��%k��t8a��r�In���VO�WsA�Y��Ʊ00��d�)1���|١�ū���0D�ލ��� `��MU��~(l���E�� XZp�c�[T��2w(c����K�� ��4�,b���s̰B����ԩ�j��\���K���zC�Nֵ�������H���`A���`�p��-�l��R*���[],�9_��=��P3�C��C���7?ʵ"�$�mݨ~�+eF�T��4��C1� ����dEȶ�N��}���������+-g��Q�ˁ��+�̤{����l2#��vL�?��.�DۙW�<���p�a��b�����Ž��;J$@޻~�程��v�%��3-+s�3�y#�u��bn�טJ�V`̭�s*8[�`Uaɇ��.�;lw$��ݹ�^Ñ�!����.�`_��L/�Y����]�Q�S�_����� ��5<<)�Viذ��K�/P�7���9�,����6L^KJ�k�]���T5���)},��bu���6i��_�4��^�E^�h9��9LZZ�?7@*���A����d����z{����cH�M�|z��|�jB��=X�o"��L����F��[P0~Q�~]��f՗���7-$���}5�^�)�!�3��Y��R��܁礽��H�}/>Y�i�+컏�n^/��������}M8�+�ט��dB�(/�)�E�Z'�N1s�X�M�1���V�=�~���<��������7v��+������i>�-^4;�\W��7��>
~�.v�)�u�T�b�YQ�wJ�09�F�9`��J���8�t�A� �ݚw��R�1|��۱��C⦍&f\O[�2��Tۨ|�u�"�)L��C<S��崄�F�^<����m�>� �{���5��e���p܋����+��l��4g���j���D���[�<y�����ٛ�[��'䥪��7f�2I���Fp�E_v��7����kF���J8Վ�"���x�W�үU~j����v��2~�"��+�D0�O�pNβ�~�_�1���C�*#�V$��ԓaq?xn+M��3��V�׋��[�VA�iP�d�vt]}�q��/�Aa]��xX�����fǫ��gL�ߛB�umwͿ'�s�׉��U�!"/]$^)6`}���ݶl����3�qcoIN��3����Ɔ��[��OqQ ��SN�!�_�����r^��D�YK.c( �����i�;�����^.O$���w�2՜R��Y�r��Į�k�%������9��� ���w)\b���"k��6şr@'�o]��w�E!=Ńx>�>�I�-z
��j�<���-����#ql��cI0a�U�������D�u0�#D(P3�n���ޅ=O��)��L�1�͏�R�:�����l.��C,}Q�h��؟��5ޯ�NU���������v�FD@n���X�i)u+�Rqe֍^3�`0��)�~Vc�珕����gq�b����vn�?+��T�Y��ڏ��8��}�u�2b�Et��7l?3�}=i��wZd+dS{WĻ<#6=z�e�
��+�?L�+�8�jx�9b&�/���-q���UE�X��1���%�Qo�d[: �\��*��BvI�m]����oO�Y2��m�Z}�/��^�����}c��L{9X`����|̺/g�����?�aN����z47�dD�x��=�p.��9�`��Ɖ�S�����'�t�9⶿��U�i�1�jR�PMӤQ��<N����3�a_�C���a�����дrx�^T�@�kX)fAG�|h������:�jP�9�B{��'���� �2k�= ���wT��i�	�����R˜�SVZF�d��#���{b�Zc��F8��LD_);����/�ب�n���*���E�.;gp��;ic��`�y�e?`O��:�Ƭ� &����kbrc�>gk��8��_l����r�hnw��:�/>x�f�R�����f<'�o:%�F&b�������������6ޭ�H���ʡ.�^u��v�[~9��(mi�3����5��#?Y=tT��o<����.��uח�����i]لK��{�q4A�G즔)����|ұܿ����"8�����O�����^��ҏ�*(���n�"Uq�GX�����-8#���w��p�}�O1ǫz7�����Ui�qY����nE~��h�"�"�Q�j�֙�y({*����?���4��	��:����7N�ٶU���B���!�1c����3��6������H�֔>Fe�3����M{\V�!��r�)$4�r�
bm��uyU��?T�:o���jv|�7���b�:ݗ��c�}[lkjS�z��=��TQ8]���yt�lb���u[IMD��W�z�S�( m���E��R?�s�b���y�uu_W���+����0��%��G?yK�%�E���i�C��Ӓtϸ����d	:hN�x��̮Xm�e��,O�K7,�)�#�ik�H��o���A�t/㼝6��D�% ���ds�=�II�U��;�雟M����C�a��{=/vӿ_8Ix�(��	ȖM����KI����k��|����%v=��.%�F둪m�j��܍�n8r�����2�T��OeΟS��"��h2�ܤߖ� X��w}�n1�f���9�a�w./!�V��{��^�.=4�����Ji$G�-��(��봜>_�\K�l=D�Š�e�L���+����gĀ��P�J�R��`��	fT7==M����,vX�}w%A)�uP��������xw?Di&��;�q;$�?P��k7:�س��hGC����c0����0�ߧc����K4�eB�8�,*Ã]o�'l��n��e�3sj������w4�-�RlX�<n�d��L�M��xs�%<���ߜ�¨Q�/�)#�t�M����C	ۘ5+A��+�]������VV�i���^4Z�i:iDW[%���;�y��e�����F�/��d�m.�_a�:Bjމ!C�1�sGNܞ:��]$�Y�?��#u�����HH㈔�[L��:��^2ݦ"lk{�R�Rq����I���g���Xb��V��	�)�Mr�)wzCѼ�>d��Mtj\=����]ש}�@�e��~��^�P�}��G�Њ��h3����u����3��Zc� ��A��Ȋb8¼���|,���V��}��I eGv�F�s��&����2D�E�l������I�n��xT%�69�b��K��F<����Q���_,u����a���,�v%��g[�5�[_c�P�� ��ⵅ�Y��o�u=��֏���V�l&�c@��V��\2�5�fsܔ���s�Q�����q �#��6�=�Ƚh�)���.rKj�y>��>�9���=��%��X���J�:���_ͭ/NIɢ��@�S�5!D�|I��: bU5�k�-�F�^��� ��8��RI�X�"z�Ak	(�16��	ք%�����`����h�� �5�1���� ���@�+���N��o�|Ŋ���E� O���e��� �2���%E�Ŋl�e��7@��[ tFDaLYw�X�[�]����ss��w<����
w��C�bj�~�����*6Cԃ}��5$������s?^!$%����/Z��C�����?��{�c�7�4J4������_�U#���r��V�q�N�Ŀad���9^[*A)%�径zmG�����?���d3�U�_=*j,+��zn�(2:�a�ڂu�^����4E�������.�<X���������xߜl�� ���� PV��ҵ����v��t7O|��<��'�l�}�ؕ��Q��L�+n�,uD5UB���8A�	-]2�Z���K�a�����%.�/�2~�88��}��w��JΖ����(�R�t'/�\^�_ϳ�~�s����Mr}.��'hs���E��YԴs�Dz�������]�ld��W��h��Lf���p�an�f�W�2���	��M���6az��E��H���2)�b��t�e�M*����}�d��!���J�a��ل��%�J�e�93aH�N"��ڛ�mL��U	ڢ��G��E�%��Hl�0�.���S�ȓ�l�eS���5ڪ1��a����h�,�U�Ӵ��{�n��V�Ƕ�{� S�`6��8Aѽ�S5�J�����QI�tG�E����d��G��F��܋�4���q�Y�i1c�c��
"�L�I"���*�d�&_�V�ټ��������.��5U�(��+�A�"_W&f�����A�yl=�?b�TƁ@�"⒂����|���h8�+h�k&�ßd���^���W}�S�"�̤n(;����f5)$�d���e~0?V��5�,�m.O'�	}Fk�/l>[ɠ_���$�l�׍��������r��s��<~g�6*�/����u�/��5��-�����K[�.6�*�q�Z�1{���H[�t��(���e���@��x���B���Ai �R0zN����@�f9�,���i��w���E�L��ڠaG~'�al�����R��욭D�j�� �2z�Y��h4X�e�S�ޗs�U5렀I�aM�/��K$i+H*c��������y�4X0��F/gL⋐��@8E73�,�-O]�Þe���DĺDa�/����SX�Ly-��Xta����S�n#gnt,�,��8r1�%�ˊR	��k?=@�)D�a%��\f�p5��}A��a�O׭��n�W���I��oxr�I{��)5���T.|��ilf�G�RLimze�B	��D�Id3$A�?M揹�/�o�ƽ�`����<�"��݀�����=�#,8p$[Q6axm��C[�Ow u��cf�&�Z���ʒ���H�ᤢh6���p�ĐZIK}��;�W���c�qI_X��xb���3M-��An�{
aXA�i���?�2�<���K UqxOʮ�
;�y���񥱤#�m��ʾ�Q��P���u���y��!,�����1m�VY��蛃r<�$��Ғľ
|���\ks<a1�VJu7=Ѳl"��@�m��:om��?x��ݑ@�����\��2����K����J�]Pt{�Z�CK�W���sfA�ݓ>�V	������4qI��s��K�V��h�@�Ɨ,§���i_��S�{P�t)#ŭcٓZ����pS�j�� :�(�/�O����!�y�sā�x$�A	����}!zX"A������>�����H���n힘��L���&�g�LJ"a���Ь����C�d	d(ˏVy��6�{���	3 k��'�#�vC���]������5��{&�I����+���_D8�XQhj�^�O���P�'�I:��n�*_����6�_㼾�9��b�f��݄� ���D/�C�x/;�jeg֙��=��{a�v \�;p�j�/��&�]�{�_����$�T�#������g��kzf�w�Bw(�	�9���Q[t ߤ�U��NeY�S�,��k~��[��k0xՂ����&W/��pw�ֲ�����R�c��� �Rn��g� �ꐎi����"��rV���	�I|��@q����3yЗ^pcF���s(�m_S]���z���|�Q2�oA͏����:���_�����.#�k͠�{�e
z�=d�yn|C_4y�󫳙}�����%@���I�4 ����OL�#���
ǊnU#=�ŪC`��T��Z;P@lJ�kT��a�%\`�-�)*��rxݚm�Pj��{!Z��N���O�#>����Bv,�B��x�$��д��"s/j����>��k�!3���\�8-Gmo����PQ�d�e5;���,��G�j�q���P3C�F��թ'I/��.�N4��\E��nE&uë������#��'�]B!����
X6�c�kʔ���ƭ�ۛ��W�'~J��&��V��D��%!A>�a�%5�e5�������hȥ��.��.�NUY;'�z�-fm�d-��w  �(o]�JA�Y��Q��"��e��(�ޙ�[�����N!�i�	��d�Gw)Wi�f-q)`�F�RpÒ
���V�� q���$�t�G��k��NO�SP�P�1���g��QG����62�?\�0ng-���+��;5���o�U�xm ���?لڢ��k�'�ֹ�o(f���v�>��QKM����o���B���Ur-�7��PV����,�[�5��XH�~��k��p X�x]&x_�b䈅��J&�AOE�d�A*J�cA��Od:Z�q,�Ͳ��^�δ]5�N��MO{/Xg��<��i/?kR��Ý56k�8)�x��nC�*�>�:׼UE�n�h��|U��O�>���w��br,T��7���u͆ݯ�$)�KWh��O✷��Z9
.#��[8����`ߒI�B�]M�$���Te�8۔0j���B�'�}6�/?��#�u{�H���z)�o�f�|U9��������l��k�8��_��U�
����\p����x<,|����ҟ��`�r�r���Xu��\9\�ŴJC��C�U&ᓤ�In�]BOk�SY
w7����:k^�^�����{g �?���rL���8���)T�q?�"�pj�Ù���Ɨ�����',lEh����=�x��*��M�R��ɲ��b8
�z��OQq6���K2	W�r�s=�0GEK���`�}٠}z�k�ⷎT�?s���c�o��JV̕�(F���ɃVR��o�|x �л�M'����IU�������\d2k:����0}`�lo0vS{����G�.�60W�ђ���6Vz~�Ma3&C�^��v��H@"��E�Nu,�T-xYc��!~$8�0m�2��:����޹��O�O��I*3�#��i�l:�������N���z��� Eǘ�D�zZ��`���5��=a������p���7`<D7�@&t����Er�n��6nA�j-�翣o/	����v&�U��F�� �Y6P��Ep~�Rգf��	��#j^&�Zk�qf�/��&�6�Rf��h#����Y��Mh����L�2�IdGy��1�kU$���>�U�	�lʿ��;�	��|9U.y�N�'�:b�WJ��,F�m��9��n��������*�px��9�b�5��R/f(�����	h�ˆ5�v�$~&H�u<;J�4'#שx�l�=��Y��'���G�����M�ɚ^QL��y�漸�\kc���yɐ�u�u#���c�h�ɵ&7�����ͽs�aW5�?U�<Jt��^@?JFpA��u��rD�����G��̤�%�����[�)}]�1�����ի�|�~��Ti(^�&��M��'��`z�)�YJzX�+7���E!F�>�?�E\,<�^��6�,sTE �w0�Uj�y�[���5�tX}:U�Zz�ɉz�DC-�.y\j���}��a@�M鿑���Я����(jJ�`��n
�=�z��ݛ���0��k�'�~�kXM+�g(����]���r�(l��ո�Aɣ��֨��b�R����q�j��`�S��O�/�^B�g�
33B�:�i(���7�~���A��p3���nW.�UfZz�@~�0#� �j�o�z�j]w��,����<Z/��y�e���m�k_v��Vy酣�3>�R������(��z�]�"�W=+���'�A���$��1nEe����zTp��Si��Ź^A��%�~icT�vv��o]���M``�X��~˘ɢ^�A1�Biɼ���7�/����J����{���0�ln�+X7�0	����/x~Rp���m�PT{ɝ�c&a.C:�7Lۦ���&��CR��#�0�������e�����=�dԳ0��O�+�Ay�c���n�^n�g��q�'3 �jMO�[N:�7��@�7I�E�t�ibt�i*�]�W ��^v���C���&�O�5���r͸�����Bǅ�
m_����m��	,� 5��wÉ�����.b���8`���I�\]$�L���[���A��t���ZV�s�r���&<�3��葖����oRV�+-h%�L���.3n5��-����慹NɧQ��O�+UG6��v����x�Ӵ!�s�
��ğXN���r�j�D�E���[*=��0X��Ԃ��.x{�++��BW;��p�̖�:�H�Fg�+����K{��pΏ���ƽg��'-�W)�)O[�R����;OH���.��ѕB��T12_@�]�J\��������M��UA��'!?*#�u�:C3��w����i<~t�&����Xu��Q����� ���o��-p��|~!��(�
V'2(\J,�i0(b����n��qD����ur���+IG�
'.�+�3{�-���Z#8�M?���|�AUf�I����M�~N�b�j�OG�A:�\��ݍ��{�\�s��̠��0\Yj���9�_��h�dx5�b�}���1���O���]h�N�^<�|s<rrl�PJ�G�a�������jx�k�e�6�Px&$s�M��7E�{aʕ�I�I]N�O0��������*�쟣���!����31�� vt��D(��Y�����[�h��<�HisԦ9�n8���2�x	��ܑ�Vf�pC�M�J9��(F����M@��Y	�2�r��t펒V60�lSڄ[ϔ	�M��I'�q� ��Z�9�w.[�&K���b�ѕB�w���w��Z���Q)c~�%��͍ca���5Z�*�`�d�16h�+�*a�����^崂��	�ި�&{#�������s!}M�Kf�h{���{���J�"c�sYwc�(V�f�0c�ϴ��͘�AtZ<�'��yx��D-�F0~��W�|�W7���|��O�V���a�.���~�t.�y�"M��K*Gc])��U��H��dI�M ����d6����F�s�TB���C�Ml؝%ٟ�4�o�6�f�ʓy�&�&`��m���	�M�d�F�4�w�Z�%^g@��Fr��<u�\���)Zr�җ��j�{{JF�;���8l�V*�Vu<�6���7\y��K?.멌���y��l4�6���c��s��X�4����eC���.��5[�!�vZ˸��%�?h����^����!�O*1�-|���b�)H�GX�<u(�u���Ub�����u�j+�w��Xy��>�*A\Uq�lu��`K?1�x5��9������{�Q�kna�q�9�0��qǕHB�g�ɵ���Z�@���_R�����e��K��Y�`���[Ɍ�f���.ՋU��S=�aaS�&�:.�M��w�3��`�Z�}����qs�0g ���D�`��Y�خ��~�2�ҳ�� �ge�[0���o�<���?&�����i����o�fi2�DQ�`2�T�9ژ�f�����"�Aߵ�N�SD.L�#n���-P}_͇ç}@�O]��P�ʶ��w�9�����>�#�`�NcsT4��Ȅ	��BvK�������?!j��Uq��a݁l���'m:	.*�E�?�Zl��^g
/i(���6��x8�x��8R'菮�R:��GW��T���9kt���[=�� ;y�F�Ԯ{�)	�J�O3vw��+��"B�z�zgN�ǫ�\/�&wTƙhY�(�l��Ư��Sz&��`4@�Qw��&H���v�*�.�U(�t�M]=�SJ]W��ƠҀ����(FBVőmhH�{�������K�������a���0����5N��ǩA�č�'�@��c���q���*(�c�ļ�!х�m�!�aF�UZ��L4�(��¤�9V	u �t�SR\����zO�8N�#�A}��nJ�!�5�&9܈�.ބ[ԺG����v�K�	�rn���I�Np��la%�1�b��覎Wa�]��z���,-�$�g�_{�g���L�"�c}r>7�m��� q��eP��v���['Wr��.�e������&��,��/���S�'ݾ�Ǿ�C%Ux\���H;]4c�:?��h��
� _��ɲ���3o0��CW�n{��{�(��ʄI6��Z .'����+�z$==O��� �	h���J����ߩ��� *j��5a�ю:u6�ǋv�,�M��
�ar>�"㥡޺Ϊ��;�$_���1��?k���#���zZ�YMo�������eר���߲5�����Ÿ��dgl�i�_Q�����F���a �ۋ2В#"<��J}�¢��2��^�FLD�L��@� z7����8���D$
ɱ��(�SJGqIx�B�u�z��7%�TC�{qq�5�".@�>L���W,Ι�����r׺�.�Ϛ��Sd�P��u+ӄ�MF�P�[��)՟�p	���������G�x¯}��	2��0�g��;"���0����k�!�B[��.�c�Gm���v4&�&r��dU)�U�:�
=�,e��%�Di������]�p";�<_Y�?�v$'�2���}�|�q�� ��h���D��]^�}�H<�.	�!�za,�/�CԐ�v�������d-���=s���=L��	�c&�x*���e����"7Z���XnT�9�քԄͱ�Md����qY���/!0���U�w#^"�sx[&���7�Җ���f�f)F�[���W^�>i�JR��t뒕��p������[��`�F�(���m�q���/�h�ҵ2b���������-~�UƯ.�r)t���No���Qe����_�'�\�&�zk�-�!�If	��*���̓++�^�C������Qe����.���І�?�c�k�+�iJ������>� ���>٤��X߆k�e����3O���u�p��ZD�o;�a)���A��j�mmT�xA��c�a��vC6�<r>��]I��x[*��p�5��?��3��Zb��.�(2~����ЄT6�o�"���ۋ� �=�kj������҂Z�pS�o����q����a-�Н��uӼ�6���N�6���XٗM���[�j���R׋�Wp��X�G0o�Ϗ��I�κGRH��_9�Ƙ,r(6u:",�z{�,ѳ�_���+58Z��,5��;�ʻ�- �'�W�Е3�D۱BG�<�����9ܪAO':��ogL�%�?�o_�{���V��I�����d�#�Ʒ�����f�)�pj|�����ku���QNy��㿖Ź�х��T���KR%�ē��;Nc�7��'���W0���8��x�K��p�Q��ǈ����(V�{ʽ��VGa�#7[4M�$�����(v#�PL��f��j��7n��:�EE��,�� ����,��L�<�����8�K�U�����
9����g��rQYiX(o��a��i�*��v��<�+r�H��=��󪋊
B�
�K���q�z�}�5�Ӑ����|Y�/;L�ΒԶHi=�x�2���;��R^�U(�Y�C��y�)�m�;�̖� ��!0��S�R�Ȅ:����S9�@�:��G�(��T�z���I�(�`�	=$;d[�f�d,uv"�"�Jc.��/9�Oa'���S��B�Z�j��%��`�v�YV����~x�<�0�\�{nը����^߆���m���51#��>�E�w�M���5��|G'��-��6v�Y�_^�)�J���� �GO�Vk���	��մ�t
��o?��Ny�x�M��8ll��	}���]P�u�'E��I��:Z@1���:�n��fJ` �-�2��S0���ߢ��1���}�/ta�tR脝z��Tv���Yl%�;�/V�9AO-�W�#s-���p�w���b��%��խ"�I[8���A�5��+C�Mi��G�����'���V�J+�d��b�Ƞ��ض�\��i����0	�e[�nk-�4�_ �ݎ�J�!J��H�c�#+��Dk���;Y��,����NMP �,��� �7I����[����h豰��e�K��5��8��>D�V&��eF�"�"�ܽ�ᦊ��2�Ps�w|B�g����4��+֯��4��^�*�2x���n����`%��/�#:�oO�����@�"�K'ǌ�a�xo�l9���N!���@r�'6�F�	��~��}��3ҽ�]{�P�D{)xD�P�Cz��#+���\5
�����/i��DW1��R���H�`r�0v�_�M�F��3k]Y���^���3��7
	ź/W���e&�q3�T�I�M� |ٲ�Q�_����
�$��qR�tF��UwI�5�4�m�����E��n��s�<ɍ��=��s*L��#|)��Mw��^2��s�����r/9�vj�h����uF��&w1���$��#�M�!+P�LKLe��y����L�[ޫ��?�Ɖ�,!��A��;��-���A����\���ޣX�9U�w�>%�lU"�u��cӖpY�����.�� ��
�'n��oe��O��V!�&q�kN�0���؅+f�ʩ`-�2�{��K�B�!�h�,��Y^��e�%����Fb�"!����F�
�Q&҈�:~��nW��#���1��O��w��3+ A{�Y4�%1v�	3��\���G.��\-��Dӟ�P����ɾ��_ŏ�AGŉ�M�-~W|�!2�^J�M��̩���?�I�0�AX����� ��t�s���j|El�,�T�|z�����A�C_IB�橰����y(��H4�f��z�ʹy��hD�[�{�vy�
a1ɜ������]�g(��6U��Qa�8�xu��C<r���h���ܞ��*Tbb??أl��SWA�Mh�U�n����I}���j.|��4��ۛ�Q�Y.�/&M+���+���b$� 0^[���*�@���BbR��S�\�xp�5c�x4׫�@�+/�=1�ষ��եzťovw�\f���� ��a��"�)��ޅ^&��9R~�|�p��u#�Y,�G#I�ŷ.�6���i,񷖾�zĦ2m�~���#T�y���?Q
�kec�b��ʑ�ړ�x%&�[������������e���?�&�\�@���Q��9�w,��i�����Q��>� �P�*	u��0y)���\b��x�OqS�^g�ID�ct���7���}o�7vc�nl5���6&Ic�1۶���m��;���?�K��s�^{��9s|��3�eft�MRñ���~9������uf֫�z\� �����t~���D�o�-����Oo��J�r�=��hr_�ФUC�=R�%�kV�R���uAkcl�y^�����݀��9���6������`�I�6I��Ҍ8��9b��~\�l��$]�;�8=�Pd׎(�1IFx�VV��)`�Ϲ̱�!��9��.z��r�й�x�"�2Zć+u+,�@:���o�vF�O~� ��zs%tq:�<^����>�A�a�p}�F�i�,��e[��]�@�sDO:�
�l3������)Y�]Mwy�yn3�R�e��a��7�i|���0���32|�>I������XB�}�俠3(.1~�}����(���`I���礤^Ca1$��>�g"=��E��חZ�Ϡ���f��<�=݅e���Ĺ&��V���M�C��f_�����K��e�h����w5}��US���S-�V��9Դ'͏�_I�A}恼?a��6��y䉷��d#���i�2�X���Ǔ0��ƭ��r8�k[O�Q��p��@/

�Fr��}+c�Q��@84��H/�{xHь>t0��v��⮳�<*������T��6�C��̪Lm�����MN������E�܉0V���݉��u.`�a��O����v�	�R�SD�R1P��xL�*�Ӏ��ZA^'S��!o���{�1�(�7�'��af���ȬH���
���^��.���m�����3&��.�+ ����Iէ�S|����0AF����ͪǬK��z�LS0E�8<�K.�@6�V~XQ��2X�Թ���ĦA�E�7�>'��������Q�߃���ɒ����u�v�^}>� ]��+����`�8Ek3�h�䭓+��G3��!=t��tL�fv�/�o�OV�'c�����L=7�4�N�ԇ0�z���}�������ᔻ�N.Y�V�K��BA��J{�V���Nq��wu����!%��pmM2a�0��܊ܰC�0��9�qE�1���h�J.�\8��Z9ݙ����h9�#�ݫ�W`����?K�'�r��=#�nr����V�/8���/�+�xQ?������I�PJ�����g��}�����k�ʚ�W�	;7��>�4ᵴz�E�ݯ��h0�K�hD���t#W�q��QL�߂�^�k�<�J��mǠ�������o^�(��7 �C󫢋�6GmN���������4�YqL��Op=��tٿ�I7�<���
�� }��ת(������6G�	v�@^��nۯ�{u:lx�xg:�^��d=���a��]��oщ���7G�-@�.|Xl���K5P�d�3�bhT]����
4�loxW��+�L�Dsb��fI�����.8�t���sc�ݣ�L���*��Kk�B����ga?�>Lё���s����	���֦4�AX" �ɛ��C�Z�����*��_ĭ��1�d٘�r~�#�]�/"�^��A�]���E�K�G�V��C��D����S��=g�V�Q*��?�	�|	
�	�Ѳ�����˩�$ ;�V�q�6��~{��v¯+�'3�$1��Cj�L$���U<~ZTS��#l���yekxy��0ο��0�x�a�P��[�qyR�~�ڐ���ӻ3y��K&���=.յ��_��tГ�)��o��<%o�C\[��#I��s�1��v�y�T�/K�����W_��4���b�q��'ogk����7-ee��Ir���B\V���;C�SFrD6�Q(��,ǚ�#�Ƭ���A�������+�د����so5j��bH\(��-�df��=�z��5K��87��`�B˃F-U>0M��C5/���8>B�I@�^G�\�U�s��m��}(�,,�p�(�Υ�^��SZ�/�sa�v����Om�xQ87���c�����Y3̗h�����\mH�:vsb���|����TF5B/����-��jc�tϢZ�l����!צi9�U?Q�M�R�)q��
vEk��%��|�'�8�3h��J��R1���	�j,�}���;�:5Q��?���uVQ����OA��+{�32�y�Ξ�d�N������AHw,X��u������RmM�����[9{���V8�q'�B��أ���D�H��D��s�1��kBm����O�ev�@B���>8$0�H���"H��5ք�����>�|nE\�\;������.]*j��n�V�}{��Dkc�"�c����H�J?��{8��M��L���y藡#";��8���U���J�==�Ѫ��v=����g!�:<���b�u�uuN���*|�`/����zR��K퐰]H]�@?����g�׿�Ii�����Č�n<�q��#.j8�=�z��щ÷Sg�����+'�}p�!'���o���u[v�*#������N�x�&�7/f��b��ORV+��������c^��"</�kj��v���t�fӝ�2������ļ(��̤�l�Y-��F;Y����h!cߔ�L�&�?�0~U�{[��$f:S��M�C��L9��V���	 ��,�/Z6�������ݱ�Y0���.�4���)���"{�<�~�x�@�{�@9�ٿ`�cJ1�w�4[̙7����i��Bw�z��3��qCG�X��b�O-o[�j�u���?ː�~��u�3��Y�V��R�y~�*S����/�h�?������C*M
5�zv�jl��ܽ�����/�dĚS)3γS�|hz��R��xfc3u���h^�0���e�w�U���p;"�4A̈l?��"�j��g>�������!bW�"��U�?�hQ7z{����I|F%���r�ȋ�X��x��vA�f ��YٳT����H�*�BP˚��D�!k+�C U��!Ǖ���61TY`B ���}P�Y�[�y���pc�4屭�w��Ǳ���O6����O�Nk#JU_��$��5���Iw��(��ʼ�:;zgY�Ai��(��ZW/�{��6�R��D^fbo௼M�g>KP��G_���ྫྷLA�G�O���׈s�cZEb���c�a���I_�hj�j6nttL^ �2����=��^t��yd�:6���_xLq�nz׻�l�,�d�6�h���]fF/oa�7Ȕ��7p��M?��������^�J��zh�:f)�ى�lOa�߿�i��W�	I���.�� �,���x���z��{���-�)��>�-�D�>���˭4L��m�^���%W#՘!�2�s�>AIҜ�ǣ>�XE������?��S���S<��9��B���	:���r;���k�a�t)*tQ�[]������>�bf�$�tKw���l���J�X�R��nM�Hlq!D-�d��x& �$5�?"�R+��o]A2��̴3�}���^z��M�$�PV�<��h$�+��(7XO�XRu�p�_�j$�?;�|�-[�7p��uv�c��:���#�2��y3gnq���[��hd{���|���?a�IZJq%�刕��91>z��f���-K#�s�>o/W�-X�b���u�/�?0��Kf�g�b��������)�-�4X�9yo�ى���r
��Aw7<z[�F.[��| �up�b��=�Ca�eela���x� $,:(B�^���Ac�d�Ѣ_Do��n���j+�,��ޮ
�a�ރ�=°9E�*0<�P�gat��=���+���K-1	�jy���	�d�D�?��f���-d:��k1��8�����u�*�}�@���0����l����,q�����P��<R�d:�j�[*�_�!8"/����J�(U����U\�	�m.���������0�Mk�Ya�yՋ�9�� Y8������6v��ש^v^�����Eiii��O ���/���$�fO䛇�i�4�8�&Ƀ�1r٦�!3;�i>˫�Kx�>� c���o�Ќ�r������%һ�0�5E� �W�tl��_��Q��|�D4N�*vjQ7�dV���#�_���řcP�;>ZJPr�֬=轻��3O9�����_�_]�i�v��@���E�0nC�ا�&"�ҽ�Ķ�|���1o�]Q�;4��ƕ�r��ǔ6˳+��!�<b�i;7d�ib����(<��]�����=�FY�M����Ma��,�M�+#�=����L����"|Ѩ��Me���w�m����k�+wgs/�U>��`���ױ�.�y2��F�Y�&����Փ7������>8�m�H$�Z+���M��?�������*f�Aσ$,�QZX�᥽~�����rm$�ͪZ���/~f�$bC}�����b�w+�(Mf�0r��'���zw��>������	=�0�[�,���i@j��[y��a9�f�z����?������@�q��c<��Ŷ�|����DS�TX���ksDվ7�f'�T+�[��s��~|@�jw���e�h�>�a�b��oUpn	�YÜ��4)=5���4<􅟢��.�?��ޙ��,��y���f\�II?� ~���e;7)_���)f��K:r���3휺�I� �5%OӬ�]��ez��>��axuN�W��͞&W%�B�I,��ƍ��d��Oz��'��^/W<�R�X
�}?�H���=H��Z�m�Xcy��ƴ�Ϝ�q������Y���~R�}�;nu�p{�x���Gع��I�?Y%6�3ve`�
���3��|�@�������}�b�
1���,��<"E�,�{���r���X�ӑnf��C#貤\�nEn�MJ�?�ƺL޿�rN�&1ۅQ��Gv�	4)���E����;����ջ�yaj4P~�Ïw�@5r>'06�l�pRK=��s{�߾q���\���i*�a�0�ڲ���f`!� �pò���ޠ�嶦�`	��M�b&KF�+�5*�T��"�����"k�l�� ��
-�N����Z0�Y��S6<���KCA����>����Gl7q;�v�9r#�B=�j�D��=t�\�2�x-p�"�S�lߜ�%ޱ�H���/�x[i�g�z���`30m<c���t 8ۙ���e�(��]��! �E�F|D�jE��h��1��}�*�>���N�I���U��]�kC�[>�Z��ʻOW�쉌Z��C�j�+�#K��n�B�o5�@_���^	�?D0^�IgzX�ʔ�&P�OZy�~x�Y+�~�ɿ�o�( ����ZD��R#ꉞ\3���F���.m��Vʉ\�t
{�Pmǚ��,T�ŊEϭ�����F����e���_���/;RPw���QC=Ot�oݦR!.�V2nu�T§�t`�3�� �Q���c�י�V5�{[z|5�����|�p�;�W��D�N6)�5���?͈��hI�bs	��J3�nn��x-��w�W P	JꉵY�x	��Q��m�P�Y�tv؅��<�2S�҆�9���!�\yaC��.w�Yi;�;7�"P
��f�"�����~~�ԁNk!<sn'�1�Y5)�����|y�%�� =*�]8�C���#b�����Jz���lI�Ex+���>���=�W0.xka	�-�V;��3F�2v&��bat1��`����;��h�:��j�l$¢��1�q��T/��ި3� ��P�%&B�:f��l.����q���e�st�"��aj�`�\���0c�p�Y��@���qN�\2@-��}��s�!��z@a,����m�NA9�$���؎��˒����ê�9��$,���Aߡ����N�p>�J�H���������7�J1n��d${��	X��PJ�W%6/��ȆvN`xǭՅ�}l��(F�b=������~��4�L�a~�����1S�D�>�BE��1|«��Q�2���h�'q��A s1���ѮRMԑ.��Y
3�?�,�GXu [Y�kԖ ���I@��t��0&���Y����(�<&�=���v��O��u�m�3��9M��2\��#mu�ǵ4�O/����6���U�S�fGm����[m�X�w1�s�כ��֗6�:��\Y]I��a�O`��s�KH`!�8/�Us�ѯ��K����<��n����8�s�C�ۘ���'.��r�^S�����U)��9x=C'�WW����p�G�9��'9jL�N���l[E���KH��Ie��q�+��]_`��o���N���Z�&��Aɓԙ���ͭ�c�h�k�qsw��=�����M�'2���4d�b	\VZ�[��ls]}B��}����O��P�c������C}m|-S@5	+x���~x�Ω��F�ZD�%��'�!�4�j�x�E��VI#tRsu�}?�B� �H���M��_;���k�=��]5/�{�kh
��W[x�6�f���Eee�(�Ĩr��x��l��JV���|Y���L�2���v% 鈈a���f�عy[5ڜ[��WW��;�W{��k��@��gBS�a��I4P��7]���<��1�bA���*�jZ*���)X�������P�3״u
le)zхq�/�q��_S$�9E%NV�k�F�S�(��������b*w�6"w����B��U�(��7sS�����o˾�� �:��,�!E>QME�ץ���Q��FHr,�B3`	�V棍%5'�U�k�g���F���kf|�z��袕�*糽qS��4q���5/u���$��z��_��?�o�c�w���l^��mf@Tv1�_=��5A�����ǰ�g�ou�I#�����y@����!룭Q�k:������� ���L~H�(#u������ 3�SZ��|���Y�Hk�Z�lk��kdrJ<�p4W<c����#�7�G��R�+g�;�)'��N��g��w.+��j��ɠg�TH�Q��2V��o���_���!�Ӄ�i�3m/}��
oC�`%х�����B>V�����8�fɔ�����Du�Q�4Q3�ߙ;5 ��wW!�+�2��R$���j��(Л��<xq��1C�;Vষ��Һ�ޅ�n�D�_�[f��qЎ�S�|�܆��g݂}����~Q�}�'�|5�j��������O�D�{~Z%
p$kA��NB�tE��9��$�i*/��)s�=������;�vjn[3�S�x׫zFSr�.��O�),�g�����ޏI��݅k�����>�X=�E'�B"c�k�v��缡!���w-�㨕���u�韷�f��u�U�� ��cm���W�G��&(��%v��A�>*��Ac-���av�V@��ؔF1n���#�/�����^�Tf�kZV��';
oN�}�l�2˗͞�-�I�(�j���D�b���d4~���Mh���:m��.Q �4�+�b�|���]S�N;��Qi�lvA����vy�
f[����� @�6hU�'�ҪOt�a,��0�@w!j�p����(*Ʌ��|1߰�6�]��Ιkv��������OH`n��5�S���`�)K\*�v��3�{��m��v	ſj�8�w&��L�K��
i�~��"�t�_�+��,�>��2��F��l�i�`��ɜ:�.��)ulΠ�Wi��¦}�Ǉf��!�V,���W�Z7{�F0�.�6n��a�Q-a���HS������R���Y� �BB��,������C�z���ڵZ}Tgy��E�(�F	<��pG�x<W�g��6�5���l�r�w��|��s�!lt��1^�N s����̭D\�c2�R0^>�v��9���63,�2���>���kJ|j���+06�ܩ��/��Ƿr�x��b�F��:X0�^�Ux{��湄�&T8V�+P�����!�L����}�|J�������J��뾏� �i`9^.\]}�2F��F�iا����&@�����b/�6�����}:������h��ߣLth��g5��BBxω ���23���lU�����B���?l��2�ɦ���|#�&��8�]��*F}����(y����7^^G���<F���?oi��7߷�"GjY��pV$]]v�|NzN�H��.y�D��`a����p��е��NoqTN���?m�0�fѮ����ny���7NW�˗��<��?!�?Ɓ����pH��Iz�cM��%����n�	��`�+�����[�[�v�� ����]�f�
��5wǠ��&x�ù����WW�0������,�s��tp�.����c�#������7_N����y��fA��x�T��m1^! {�T������=���>�4a���ՙhe�짾�trk��D*��
{�o����~0�Ԭc�����:�Kc���80t}�ح �!F"�T����n4�uJ����Q�Ǭ8]'�AR���i�y8Ѩ�Y�dreB�'���ȪQ��KH�S��	M}ee4�A8��]+=�&�$��8�){�0,
�+Cƻ��rnU���I�8�zǳD��Z {F�%v������q���le�7T����h"���*u���#\��h�@)?���^ܔA����CV����H�U|s��j4�Z]��[�������U�c/uAڠ�@n�/G8`:�������\mϵ����5�+H
R��"�Y���p�ո�L�s�oo+�F���aw���T�eI�OL�3洲Е%0���TAt�{�H�@��}������Bz:�#�}c�%\��;��^�KP�\��R	c�":�M���(��{iEl����H�A��^�HU�
�{��k����E��q��4��ɻ�'׼�U�D�����������GH�=Y�D�m��!"qLN��J��?>$�J�D�P�������Z���VD�/i�W�E�<�_���`���6�v���]���@�ϳ�Z|��9]�[�����%�lⷸz	76����u�~��x�L��7�Txqy87?��+�i�^��g��%G��^���xXD��if��s�j��Xw��c��{Z˙�A��@�K�7������c�wR$��h�7kߥ@ն��1���T|�9ҟ�h�L^
S����IC�)-ts��?������;����^��'xxޚm�J�O��zk��)gՂ�sv�WR����/xxb?�ނ�<�tO�� cc�7U~����\oX	�B��v<��j�~�qC�'��^��xn
R5�ʑl����챓z��@��B�`ݥ���[�eXx_���f��7�,Zr�f"��d�hˢ|6}cNb"��.6�1�j]r0��Ho
���=н ��\S����b�=�Bh?}_ �����:K�7�?�5@���fU`>��)��́�?;2"L���B��P���/"�Xb�6Qh\>��Gp9��Pe�9�8�J����%�|4�R�*��p�C��9��/�t�(&����e��_��i!���鮬rQS��� 8k,��ڒ�g�K�XM��`�B+�y!��wtֻ��v�\������UX�t�56`���N<؜��_x��N1�P�][�8��8��_]�}�eU���ÿ@Ҕ�b�Wb��P���f�
i��̣'��~ϲ��K?�r��4?;{h5.k���-�B I����G���f�[�e�\�/|��Vȟ�	��l�Q�T���/T�&=^j�4X�jj����̅�,�^�����ʄ0BSH�8{ڹA�w�
�����Fh� �^��8�ɩ.�7'���]D0_����\)Ɯ�~�9ڣ���
��vpǞr��dg�Ր��{0�%:��Q�xQn�(&��M��=�-Q��|�����~���`�mO���7.'��лo^&��|�e�c_�>kٞY�}ۛ�NV��RU!��HbaBD��eio�g�B	#w�(����}��n�qF4������8�x�rk�Yߩ�w�ls�G��/����Є��`�g���R���� 86�����-��o%`�R�eb$"R��_
������X¿Ͷ
�n��F�Z�I�9۴j�"���ٽ����1(�o���ud2Ja��6��=�ɜ�H+��҅���U�"#�,�!�|X0��fp*|�t(l�񃈑�	z�a��O~���5@a%@�9�(f0�$Q�\D��	�@��ܪdu�d�jo�  ,�y���C��j�|\��<���E����E����� ���3?��[�!�7��Q��1�L�gf�;CRQ0��Fg:t1���_ǃ�(¨>���NxL������q\i���Uԉ��`��+�y
���m�3�j���wZ���q�Vװ��G�iJ(���S�nH����tt):����=Z�2�zM(���Tt��8�u$����4��H�H�D�EM?$_�-�dBa�Ĵ�']�e�ܢ�~ f�VkE�2iM�o���aZӛ��{�Ō�+�">�[Mڃ$-��V�k���,θr�v\	�-?�Ei��5EhY8ZX�RX�#B/SޟOb�ν_WF�t�Ξ}�҅��tV��o�h�#�5�vt���5*�W}�}��@���D ̐���`�aj�ߜv``P����)tX �W~��vr{�F����w�C�	�K$A{g�+v�߳8�ۤL��X�r�@��j�
��	ii)��	��~�Z��]_�u.�fW�}z{�Ú֪w�6������$�3Z�Xm��R\��������gxɟK�� |��٫��1�@����.����e���Z�%���h��U?x�x�����V�&��K.��c��{:tS����H�Jx>����E��x��49|F]���: Y<�i�3x�H���sY�n�48�a��6��On�ʿO*ٯ���B|�+���-��Ȉ��M��o��|����?)��l�o��{,͝:в�]�*,��	�-�����*��t�."�s"�����}h�Lr�]��5L4� ݛ-�㇜��݂�/�c����n�8J��=(��&�{��9r�M�3���E�_y�k���a��|�L²��R9�Dià��� bGM*
s�F��w+�t�opn�n�KT�~��n�/��e��`�Z/�Z(vvT��JA'0��T��J1
�Xz����V�Z�@��gc�l;8OS���X3�o2�hW��|"��_l	&��]���˽<�Y��.��3���hy���tb�Q+7�)�y�p���\N(Moܭ:�8m.ۜ@^ ��5��<�ԅ�}���0Ai�f��#ՒO��,��@���&�nM2��8i�v[�z%����ѕQѕ�������,P!�p�^�͌�}�q{�N���Ծ3&'na���b�$�Q[0��5���O�;�US���Z~�xӲ_$�Ч޼RA�ppr��榽g��PI.3��+�� ^�<�
wHv�Rd�j`ÅM�e�>��7�I�F��U�ov��V���U�����FR���o)����+��wY��Á}j�g�Ny7��#;�va3�� �ж'���`|�~m���m�5��ڭ\���U�r�_C�Mի%dy����P��=�[�j-�{�h,g�����8��&�s��w�+��j�Q�G�ܴ4 (`�!���\��Oȫ>���mj��w���e��x�&&>^<!*ۤ:��X6�0�����>[T�P�e��������K�O
�L��J5GϨ��Sh8p�H�-갟�S3�P� ^圬|����p���$�HS��b�18V";x�� �\���jW�&̸�2�DI�P�EQǠ~H�Ui�iu����_�K�Ԗϻ���a+��<Gf�Sћ��5�y�1N����ڛI~d�	N,�:�W�3���
��vC��X�a��ɍ���(�G�B$T<Иf	�Kv~[w���Xz['�.�d{����bpk�2�q=�0� ����Eu��0�bo&
i(ux"7_\�X�	ߖ<�y�
5@N��Y
�ܚS����5ZSk��*ƒ��EE4�o@�=��A�/7gg�F���@%rWP�)�R��xl,�C-Vz�]ڿk���gd���⸆���|�����6��9-���Wn���+i��C�+mA���
qj~qp'�-Y�@O}�]�i��\o�^�4�m�[@5H�IF�P����X��9Bm�����okyE�C�=��6�H�-��@0����\��>��I��F�����k-	'����M`>^Dn+pZ��(��U�n3��<�eS,bd%A}�dJ��%��d��G���?��+�`��|��Z.,�,�,&�MBS��l�>���Б;����S�TUD?�,#K߃Mk��f9��
ZN⁷  >�Jd*[? �/{21	5�0<}�+_�ߣ���ԅ#��Ļ-N�����'4�;�IH<-Z�|�����PQI������;�D��H�%���c���sE�k��|k�j��hW5�����h����u�;Դ��ڊ��4��H=�}I~�?X�����]�|��ty���
:
.����1ʮ��� ^��޵�zF^oT����2�r���{���c��>�1+�y>8E�}1s�t��m�7
-�@B�����B2����Ob=~0��\L6&��Jx;���������d����g��u�;9MnaHA&Lz@Q��>�;�m[Oj��`�Ch�v��*�W�A�[筼��U!�+
�$�n��{=��J���ylpG������mY܄U:���4��!���o�C�c�C[�	eb!�,�9%R�]KԂe(�t��%@���㸦��)�1r���Ag��RE�X�η���Ӣ��f}�j!5���h���^���oWث���5pĢjy�f;ym�;'���+̥�P5�Пtob�F�	��@g�B 	��.�vq>����鿀5m;�8��jh���i$�$0�/T�G�����RL�]�A���dG�f�[�-}WO��J�4{HJ°GIc��6���1�;�ȱle!�2���	lvѴs��� !1�
����
��C'�أ7�M�u��N�pKߨY�A�X`Ջ��/���!S��q�a�*+bq&CI��-�Ȳܩ�@��Lvc�F|[^�O�偗(���5��Î�2���8��$�\B��+>u 9y#8��=�0�$�_����y|��(�96�O������-�YVO��Q��	,xG�r-#_����������Ӥ����$a����\և��Zً�3�K'E�W�H��O�0���=���|[~r�]C+47�\=�`�-�tbm%�+ 9�Ӄ<eV<��3,�
�P�|ݓ.�6��s�_>����LG[n�@�F���~d�<T��Ew�c��;�
EU�6��t)Րg��9��?N�� ��}���^�e�=ȫ�_����:
q�'žZ�	�@ga������*�#9�dN�uJ��j���S�4����@��W;$M� ���C��c���w;P�����4Z5:dTs����O���=��,~��2��`�ҕ+1z��u,�m��L�l:9�F�|�=]�_������rט �XY��5(�s1otǠ�ա/Ԉ(E��1��O�,��y(�����h"bN�X�)s�$�/����kҒO�A��W;e�%����$;1�
��pfu������/@}��V���,�,V����(˯\��Ǥ�Yj���:��t`�:�V,�-�m]��cI����l�3+�
��җܵ��r��˱(��7tDë��2�N_7uA1�P.�F�OTگ[NE�j��"��(�}~���8�d�e����T��`�3�$E��� �2Aw���r�`�	J/��f@�8ⰉA\R�7�l����{�j���B���}ka�n��>-
}�=M��鯄}�1؟�(��R&�� ��6�X�(�x4cB;�ȼ�L��t�sB�Z}�rܯ�hq�Q_��mÔ9�?���{oÝ|��Xi/.%�ƍt 6�i���Nؓ�u2s�3��
ŗ�O�ΆKGa�-�n���U`�&j��y��!'�v���l��'1������-�H\_�oM�����S"�r�Lg5{��p^uW��~p-݌�Q(%��]��Щ^��h<�ax�}:%
:	�
�~�h�?����~�V���s�J�8�����'Ai8�L�����KZ-e��Z32�4 �~�cg�!�_{~SA�1t�]`����*PF�l�u���\(%���d����;��"���E��ƃb��ӽdP�YtnJ�k�;�>�@�Q�";_���ƣ=���K�G���'m�&�ɽl>�]M��#�j:��ܑ]�$>gg���U�0z�߳ �ֿ@~�c�o1�̇�
fbAE>�4(c�r;�Gd�S��4���:��B���\9� �pagr4�7h�I��T�	:1
[���wF�3��|g����˅�X�v�V��ق�>�i5��[:�x�����45)`�cm���@aa��&�Y��&�X<��/{�b���O-��>�ѥ~�����l��Y��:-��w�r}jH�$�F��0�ѐ ��ϳ�b$Z��.h�ǹ|��@TL-���0S�#=�Y����>R�y�5A��8Ҥn�`b��>�b���3�>О�gO���N�vi%��&�X���l��BˣKJj�[�ˋX#��>c.z�¯��¹�tMq6X��~�f� ��+�ٗȲ���"���E_ԙR�p}f��}��f��1��7�@W��}/TY.<��\�H���Muy�0��'�ϧ[W�TݥE��I��>��?�<�� �6�2�b��.>�������Y8�x\8z,�U4�ݧ<o����;/�ʕ������0!rt��4ú4�0�M��?�F�`����PvL�vW���ԟ�[@�+���x��S�m�}~�yō/��k���M��^f	"��h"�����t��4�=�=���&���5����,�G/a��V{8�{��T����]��e�����������\U�7�O��o�@��+Z1w�D�'<��N�%S��R zzW�ڣMc5�� ��WA��_�QY@.U�C��rG�������d�b`U���.M�E���NfH�|զ������*���b��	�I�w�	��s?��l�T��e��[�d�J�	�2����`Ff��.��ˑ`���'_��e$yc�w����	�?ޯI�DI��K�Ǐ"L�:+.�;��I6
��ACȲ<2�eg��'ӷ�j��}83c^���rR!���(N1��83����i0+�z
�R��Q;70-�	�C��t�g�~呩k#�HBD�7l���VX��_`e2���\tI�[�t7�����HǍ� >�-ں*9+��v@�J[�f��@/|4wW�Q���ة��ȡ��Ҁ#��*�bʧ9y唹7����Ho��E�a������,8�f��v��vn�'^�5`p�B�ۻ��0�rjT[��Y���Ls��p?z��2h��et��+�Q��D��%�݂��z��S h��ҫ�'@)
��.4Dt����ޤ�_��2I�?�e+r�w�nC���Ԍ�k���c�g��vx�,�����7�]�r7_�T�y.#�T��Ѡs��|8���7��[��%*l���`�v�ڮf_\?_��:?�q�z�N
|_Y(�E�k��j�=I)h�+<�{I=�����F h� jv�ʽ>�5h
��?����O��������M��G��դ`��ih���/@��/l4�L�
�2U���"��Q�1H%�\uۿ��\���<Q��8��fv �۶�&�Y�U������j���N��n�luir�C� ��>�c��E�eh�)����n3���l+�7<�6�E$���0CV5�=3Q�C{`oY�oc�WQ�Rݏ����U��Ϳ�u����d�{�[�V���op>RTy��FN��,
j�'�ۦ��������3)��"���Iʓ �4��p^p����K����6�����x�R�=�/4o� 8��z���t2�Å���ԍ`��S�����]�`�ª�i��z5%M��҄��rXڇO�@g�I����q;sC���2�@��n�E�ˁ����3��������KT���J�c�V�~���x�A0���Ǖ�\J�,�Heۅ�J��ZOݑ#C�EȏP�v"	�㮇�{F(���14Rc��=�oY�ݨ���u��9:w*m�G��肤6�[}��x�0�����
��۳m�|:N[#��xR:��5�ns�.t�֬�7k:z��ݗ�{f�C������	2�Q��
�"�P������%	���1�(�����OX��iw�0�y�;%'���o�ay���!�esa�Jem�Z�z�{���ŝ��J��4�C��	�3z.��\R�kU|�H�.o���MH�8-�r�Bm$��c�U<��Ss
$?<0�]�rֲ�<���B�L���%�x��bp}F���xv}igB%Mț�QC�	l��v@(��j� +�����X˘��<4f�*�P�� ��l�cjU�+Wm|�$,J39- �����X�|=��+�}0�P���;qƴs�pymG�K54�`�.����N ��ʒ_�*��K����-؇Dj�ǁS�!��^������s��tN��v��\�����Ú�c�!5�-�Ŕ���Zo^�v��}���͠�{K��vce���L�������K	}����t��x�y���jdXW#�ۄI��f0Jj1M�5ງ�!&��_������p�qQ}_�F�$�K���!�[�����n��n���sh���a:���{���s朵׺�u��מ�|�m��+�|�K֟�1�+�����<r��>9B��.d����*��"�}�w���Ks��PHW+M=��ԝjs'4C�i1�'z�M�V�'3����NtM���~w�y[<b�5?�39��'6^],b��]�p]����o�i�P����7v'�N��Dz�:B5�c��Ǵ%;��[���U&C@���j!�o>��m<��ԫ���/6g(#�Ä��O�g���]\���9��b��Z�U�r:v�t���� K���l��'?�������Ɖ�0uK�j���e����Od����8m1�`���HH��ދ<��=0�f�EqE�P"T�֤��/o�-��[#��/�lE��:��󼑮{neمa���D9>1�7�	)&���JR�S ���d����'��3?����B�c8+��<)��xO��m]�䅞8��^�顢������ڀ�h����I�ǉ����������O+���X&�Q���Y?�8n&L�P��9P��p�f�嵫�-��I����b�eNK:��cW-�F�t5�o�>�5��O�1s8Z�˛�Sy��Θ&�.����������<j!������A�$4��p�S��Q�M����z[<+"Ξ(3���r]v(eT�R{\�v.��<봫��$�O�M����������j�U+�\7�f�B�s�B���ri}S�D��c(�1��?GW���+��=NѾݷ�s�c���bX�^��2}>�m��l��ͻ������-6L��s헫�Y?j�Y`{�l�h;�L��\�<�w�(���%Q����E|�5�01]lIT�n�+|n�/�,�y�Qk��'��~��3��W����h��ԡn4鯪�X��~��r1juO�a��S��N�j��Uۂ1:T�����'������ǖ<8�y�0a�`CL�o[��$����j�a�Ͷ�gW�͗i����\�w^>�� ʬ��B�������Î�zW���!/L��ҭ6U�3ƾj�DU�����v}~_�5�Qx���g�x�"bC�]�M�t?�v���
R������*m>T����9�ϖjg~|$Q��*$cQ�#"�����Q�uh.x��Ϊ��rd8R�	��6j�x��X���	�SL� L���T}�}T�a�y�H��� g�翙:��7��GS��~[�OV��9�����a�C��X4d��5�d���.�����d�0��~�i���-#������s�j���n�y�y���i1���RKnu\>fF��z��K�{��ssb�1>��ћֻ� U,(��~qj�c�?)l����DUYua���+9��k諦��cH�\+��cg�K�#��[ɏ������}��L�-������9-�/GF:q`�A���J�>�&�r�gf+�2��*���W�Zyw|8�s��0QP���w���uv2�d8��d�`(j�Zju�y�T猸���f�|������	��Ό��$V�]+6ǆɝ=o�Ɏ�qό�ߌxi�Xt�1�������	�c�Am"#�]�F"G^��-��$r���<����\�hz�R�qрJ�[r=��pD��98:�g#��.]��{o�I�*�C�^!�2��j�|�bQ�V? v��#���+�?ʅ%���l����g���������$�w��C��&�y���lo���\���c���)In��v�>7�<h�;Q��'g��mb>	��a�9_�v���v�X��ӹ\Kϸ��M��L<|R��,�3��ܶ��@w,��ۯ�q��{���~�6��Fծ�1 ��)������{�8UOȴ.}�H�ٽ�!h� ���e�n���>P��XP��Wz.,&>G�ə'�"ɷ�����I*�w�� 7��H�\��E-�/����ĖZ��ndɝ�g�9�v�N��ml�2B����X�(�}X��Ո�"|S��ڠ
t�h�Ax�RU���+��6����V��uC�ٙ����O�!�uz'���ir�@5kA�+��9�,p������
���4<u*��~���
3[ww�N�;f�]���L��Ilf�fa�(�����~Qxm�d,� .��u	jё���U�Y�-;�6=Z�gS���0���[<]��>�^r�ETl>���9Gӹv��\��&&@����U]~��W����e%��FU�>����vՂg�rr:Ie��nTFY]�;��~{.�7��p\�L��!�u�R�2HE��`�6��'����l�.��L�ȽuП^���	�����{���O�iv�Bd���	�;X��a��cݥQ�"� �����eW2����S�b)����2o(`��,9�y �Ǧ�K\�-|�u����u'g�����}���ËG��2ƒ���LdR��;g�.�v��V�z�BV����y�C����)(���{���	��?�]w���*���.na�3�TZ]��$Z�G~���������\5� y�������S��{�R��J�NRL@�؛~�pu�^���1e���C�=�UH��x��6VW���H�&>��>.���o��j���T��f� َٓÅ��:��f��\
�Q3���� {�k��N0��]w�.v��`������R?�*6z��k���O>}�i[W����s���&��;� ���"��Ei5]�	�(U����3
{1f1���v�_'��:
���֑�������OjS"�)��M�i(�@���p*��_/�2�r~'��\�D�"2$��|��.�m�+%)m�v������~�<��1�_�]�ίK�-tHhȵO�6��{t�Ҋ�A>67����"v_����j�5�?�u�=��n�&Al`���z�#�~h�����+"�y�US�GZ����Ӈ�؜0Kf��{��9F����T�\,�N�Q�6��������kBh�ЙfQ���Π�&��5�?Zz����w�E�[	�=Tβ�?����+t�j��4&��'�cw۾2�u�#�nK�9�����.r�Kw��!޳�p�d��f@<�Vw��i��k�~:�2���2ᇡ�����צ-��%��x�����y���ܺⅤ�:�6J�,�.
�uA�\�.^�"t��`5�`�q1Ҏ2���ܷ��,�_|讆�~�#��@�mWz$:a��C����*�E���Ye�O����zj�#������C)����4�>�7c���Y�PuD��݇?��]�� ںD��>�|b�V#5'�h��E%q� ��,�w`���4�7 ��E�h��������=�kY�+�?��"1[�}�� ܙ�n�V-���*���Ǹ�p�{�Z|�X�W}�,i�#�֙�������<���]����fJ�&��|13Y�s)6�޳��<%�8+Wc����[i���^#���珻GT"���ɡ@rƝ��&+d^�
��������in��m��J�\�����O��~�=�D���#�`v�Z,G�y��|���%oЕ���VwTㅗA{eKO��Ft��.t�����J��}ϕ�
S�b�Ш�@2X���?�)����μ�����Rj��������:�����<��16 �yC=#��K]�wSb7N{���w��o�C�P����ڣ�=��B�C��m��1���E��#W�~U$�̏e�m�P��y�Oq/�?o�ª�ֿg9L�B�X;aw[S����S�F�腰Ob��~������&�M�2@��L|n2��&�;������6����`���t\6������b]k�sQ��QŰJB���c�y�]�s+_ 4V?��	�5S\'*\#��zS���������%\������L�h��i�HXN��P�=��'-�;���4�ì�>Y~��}EWVN%�J��s������\?�z�֊c�j����B�#��c?���)j_]-ȥ�"�:?���]Rȓ$��Yܧ� �1�M�4j!�w�E�.6x-W��\,PF����f���7x
L���k)/� `���5�Rfu�yuJ��q�̗i>п�.8��	A�?�;�D8�D���f�����,j�W�ěq	��n��c��I��c��gN�ǽ�W�.a&O����c��5Y	A�s>����@ΈmP�h(�����|��;��E�ɧb0����g'���������;a*�	~�=�d3��K��%$�=���;hݼ��x3rvt$o�1��9��iC�1 �d4�J�I��T�-����{TQӫ�������ϓ_�����|m�"�?�}:��,D��@��<,�j��u�z�+��
���{���|�MQ��5$�z��jB��?�����]N��MK���M����85��++stM�l+	�Dr���$��m"��-�1��-���bX$lr���X����3��i"�ܽ�@�m�1��6��~��u`�l�N����f�aÔ�P2A�����Qg�����Ý!b��[�{^oM�T�?oA���
��p"lI�ƌ���V�.}��x�mIrmA8GI�N���\˃M����0�tGH���cۃG]FqAI�z�(�F\E����˞��:
�	ˈ���Dpj���y�Jc��Cm�*PR9����u����ق�d���G�t	B�F�O�>�`������� ���0��	��N頌Y~}�-��3�,r+�R�)C�B+�c���=����v�d[�e�c-;�4m�-eMP���Z����o��E��}Pk�*�Wa��2Q�p��x��_��/[���9�ݗ��"�<���!��)��X	N6b���ɛ����O޳+���q�Ӫ�~C��ѕr��[X����
�ȑ���5���v��_��Xg�L����o7;�/ɘw7t�s�����ZIfsC�#�^�5.'Y�p��W4�YFc��e��W�Z�LG~R�KQ�8�Dw�> =�z5�-��2�kT���f�����?Ю�/n���q���k�ֽ.T׫�K#���� 0i�O#�-7o�g��r/,vG��
�<���O�[��������U��j���+��P��,�rR�{���m�C7@4د�L��fWz+�U��I%Q�C�޿�����ٻ�����k1���� ��P\���v��m��ɨ�1L�5�[~Qw�y������hUB7�E��Q��3��$�wf}�`٦= P0�ؗ���k��`��o|���ڦ׃�����O%1�_rt�c 4sV���n���[Tr]{����(�K�[�S)��v��lZ���m�Қ����]��<���3�i4]����mi������O����Y��B��X*��-~���]�Ϫ�}a7�:�ԶQS��Jt��.GZ]U��b'd��W�c��q�cC��5���d~JGǹ���E�o�+��k�c
NZ��[|)Xp���*���H��������#�\���]нƏ�[�y'ݢ=/J��=���z��,�;b�^Q��a�kk�C����w_b0�(c�	N@<�!�G��$;�h��M�
���ru'9�Ml.I�m�o}ޕ��x�We !b:�9^W�+�;R�l������}���eO��c�]���V�K��`���{�y�ڑNT��b����U����ۙh�cLy$rm��n.��j�+G6�]7��s9'1�������{��?�i���=X>]�`�I�,����y63�sd?~�U>vx�p�?�;=v_<���1���Z;�I# ��j�l�y&�Dz��],!2zg��R:?qj�E��!+�=��xP$�k��W��`K���I�W��7��8���������P��G�ׁ5��?Nҡ�ȩg��u;t�>�=
)�'>�����d�޿{�x'z;�����c�{��^�q�����x��ջ�h���+OD��6�g��'�e"C3E��`����>t��QL��m�_�KO��y��@�~#K}�\��/,�D��� iJ#y�/�4x]��Gm�.�ԡg�8�J�L�鐹˥����V�BnܛT�&�
Y���ÇwYn�X��'rB@i|_�8������M;���D�\��N�$�;;����kw��hhǗ��>�6���c�S~�Ps�{�%��+����Yx���å��85B,����b�TA���wN�_�bz ]&w�����ܡRDd�ks�LLQLnbٷ�]��!����J��ѸJ / �{����hN%�դ��+�w�&Z���
�\w�ҡm�Е�Y��C�����M���n��ӱ�k����K3��cD�CP�Iϥ�����Vv��lB噸�����z�[�L���Č���K���/T�v��+hyQi�.��ꥥ���
?땑i��P��H��ϯ���s4l�a�3��&d�Cd�����B����Zbp��{����ͱ�����`����]V�ƮӚ�ޯ<��Jbd������wݫ�]5O�4m���64������o9�����X�G #��o����9����d���5+���:3cz2u^�;���H~h��$z^)W�	O7��b���kk�{��Ik���e;��#��������˕��fB��f�I��nj���gOHn�-l`	�̴-Ai )�����'$�@�I���,~��B�ϫ��E��G�����oRd^[>IT;��N�� �Jl��7����~����Woj;�l]\� >Fz���=�-2�00h~ҝ�G�+]h��E)��0b*����� Vb���F��ה��Cf�t3�S���B7����\��I����p �_�M%�"���᯹����a�q]��~�����y�ߣ̽e�`�h49��6਎�dm�}v���N��J49Ե�U�^p�Z��:*ҶZh� %2��aTg��K �(�1��N��?���̡�z@�`�'��R�a-I ?)p�u^�^�uWޞ`� ����r>4����-��'6+�]�ҝ۔�������ܚq�{���SA|��J KG��_�I
�J��8�#���uf����Y��x<l�*wW���8*=��̬��ڵ/�L'�=�+IV��-M?Z���p��-��+D�xl>��W�~����5�N�6Q�gU�𓕗z���������5��U�¨�#r�����J�T{���L�|���ܘsO�ƍñ5�1��m���h���+T���L�^�9~d���5k��)N��b%Ew$s%�p~}<؀?����xm��#n8��z
�Y�#�qu�-�/SGLt�oVi䗪�5�_�EV�)�M��%��̔�j�44�ߴ8�[z��#െL�����q=Et���<�4�����������51 V��H�/g!�[�\9��ɖ�}�mH��ێ���|S
{Qlⵀ��HO������"��3֓�y����Oc�N���)������4K9�:ɀ������Zr٬L3��r���b���0���F8��k_�/��pU�	��3��� �4�L�4�Tk�Uۣ�	 UB�Z���N�?�|4����P�[���r~�-q�q�����)�S����~L�w#\<���֕�If��ՇBm{"�A6d��՝�1�m!͓��DV�n'��a�+~�(�H#�S�՞���!��v5���=�Ckj�HI�Z�Tǧ�wF�9�p����\Mh�g���v�'"���E�4�u�����ksܼ�CJ;�7���;�q�D�
|��Z���)	�SN���߬V�-p�/��ߪ"�-^,����GS=v-/�$�/�!�9K)|���M���{�Qn�myk�6�>+��d�e!�QC=������ %���'w�"��Jx�)�3+"T���d�8q��f���=�|d�z����
��퀚QzՋ*��[�w�q�c�\��#��B�e���{��b&j~�,�<_�D�3|�� ú���b���8�0?e�*a�X��!mY�t��@�.=xDu���ڡŸ: ���ww�����QU�a�ͲY�����K����;��Ż��ٖnPq��R��E��OgZ�+��S��г�f.����˽z���G:z���b��b�]9v,a�}r�2�S%�!Ԋ��Bp���Xp�|b�z��x=í���%{�X|w���N9Yf�P[~��c�@�U�g��A�S���p�I�����M~G�{n��_W]��?�|t���;�u�D�m*V����s7y��) z6m;��V��|�oP�b$7���ڜ��k���h���
�o�wS��7�Q�,R�%�+"P7"�ή��T�,IT���k���BH�&ߦ:И=~�M?���+q�q�����C��9���#79ǒ,��w�(�h������j]��h�gVCVp�� B�h,�(�O�z4r$Aoy�����@��l�h�,;����~<�=?��V�0��������aI>�	�_DNX�{<�
�����4>���N-/%Gr�As�^�t<���� ��&m�Z{�C2������9*�+�:��L<s�׍�#�e1�d��O����S1��1on�������p���¹;{�?x�}�ԇo �H"ҭ����������I�­2$\<S%�J�'����,�[5�Q����O��_]m0���.�>���+/�RҮ.R������-��R9��6�{�p�y���gr� �OO"5kz��+�f8��
ŢT��o����6��	��S5~��+���)��B��<�r�U�=F�Ͱ�6җ�S2���A4���<>�#W	__��x�	�U���U+q�tb��}8���^��*5'x�N�
�-]����Y�T\�.Dz���Y�fN��>��ɯD����!���6v�R��l*�8*�N��Y=��j��0v�0Ir����픖��������_Ȭ��ʝ�G�	���pdF+_6�VJX�$��j+�w��K�l���N$��y5��ci_�٬u�mr��� ��ʌ�ʠ�����s����_҂��EC(;�����I �E�$Ћh��yɢM4�a��&�|HR|TN���M�U�i~p+��K>,"���/r%��l�rZ�	��*���_�A�B�r;,���{�i��[��wK7��q��"�"g}�顉�����6O�����@�������,!z?��4�[ѹ���������jN�q���5e�	��0*O�v�I6	��hgˣ����f�Y�
}�Y �������٫�GDO���L򸙳�O"�V s��ʬ.9{�W�6�;��t_�_��˙�cۣW��D�A\E���LB�{n=�H�nx� "��9x���,g�A��0r�A���8�0z{ҥ�yō���ȓ�w���n��#����CZ�')��x�	hn��b���Ժ*�7��lcJ�O�=V �p�_���?���7+�(�)0|��u+�Iܴѯ�u8?2��?� ��ӿ���`^�Zt+`H���_��sEפ��C�
*�]_5_`���pd�_��ꋏ�����O��Jԁ<�.;�~�'̛0N��=���'�n�@�Z��(����?��|N�u�)�~M����N�����Y�/Uv,τ�wy�Vm��5\��8����~����"tq��I�AGo~�-<��h��#}0�{jp�/���7������n�Df Ԡ�D��Ht�V��?N= �Hx�e�=%�^f�.X�D
�Q׺�"l]�cx���2���V��hXe�D: A%픧�w��X����a=�Im���+~%�ª)���~`XnB�T�^;��\��J[�vΝ֒�>~�^��w�U���։��������UP�QP�a���M� �Q�E�z����$W6����
��C�wߎ��7�:�����%P��U�^��\�%�Z������ܲ�l����4�n��6���཰K� �M���}�ސm�׃���c�z��E1��X�y���ݨ��{�q[(�j{�ӊ��A"Gi�G�1\c�z�^�_�no�U߅�3�}z���@P	�70���"ZT+)Q�b��7�����.0L��1��ѵS��s�2�O�m�SY������:M�G~%F�{e�M���u���ؾ^7��gK)+������ku[Ej�px�i��h����T�X�����CFQ��[տ��/݂�������>)�c���jȚ3��p�1΅(�I�d17�p��e�׎NF^ �5H\���Z1z��O*�������!#�BL���Y��B_Cl�����q����Gv,~��/�G)c��Wi7�0���TDD�:f]��oV�m��E��7���KM�D� ������Q�'�c�Z�6}�;ǡ��D;�.+fq���u�����!��/) ��Z^�_���k	 z�:/c3����i9����|#x�s�p7�Bq
���������2�H���ɬMR,�9���'�D@�x�]v��R�ʨ+�*r!>��=�����K Z��I����.c���YV�U��6w�v~+OBx8��>��H*�u�|��UTZi�ؽ�5-���8�VBG%@С/�^��� ̞���N��AA�c���Ć4mp��P�#�r6�$�S[}_���׍N���gY�>��q~2Jsm7m��t�� cy�� MUs��lGϿ��A�^p����R���Ψ������3��C����_9
�A���,���͓U�D�N��vQ�m^_XQ�fء�d)d��9��]�Y^>�J��l�s�y}g�E}������E�_Y�5��C�v�}�/B����HF��LպH����֙Թ��[�mډ��u�R\�?>wR�@'g������F�*?Q����p2A��:Kd�7K��]�(���a`���8���i�Ba~1%�5��me�{��	ZW'��6��U]���Q7���#�~\�f^1~6��A�o7��Pi:��չ4�a �0�u�wD�X��4�S�|Qf�����g)�WN��>��N��Lُ^�70n��w��@�Ƥ��EW��4�Q��~�լ�j��q�7x"z�.'�����&��q��ɿ-��T	��	��6w�:K��z����#ۊ�G���2G� '��=B2�i���M��5e�E]� �a+�u��gai=���k�dVw0$� �cuqp���a�4�J&�����`���P��.��%](F��qn���s²K��؆D��6�ʺ(�%�����<8��DBu5?�N�����7����oݝ��)�e�g
D���`Tt�~���Ea�4O�Xc����Ҁ�"��O�ߥ�d�$l��˿�l�Wd��6.\?s5�uJ���1N,
#Z:�����Y��_��y�� ��k�cB�5�X��.F�L�vK����r4V����/Da&o}}�����_㯹���T>T��;���+�����Ʃ���PmUC�:�<���rJE�����_@ժ'o�؍�sz���qXa�0��r,!�����dɎ�U��L�J?�E�7~Ok����	������ �K�Q]&Ẉ v�,��}9�;�[ZW~HN�O6G��CX�/0�ž�����1k��ɋ������c������mǨ������|E
8��O��p����=[��V�e��w�|u�'�Q\�a�pnH8�I�W�3��ֵ�s�U����y�qZ\\.W����E�yI�?2�l}��jI�,��a8��&cnj�[��Us�Yx��d��Bپ~�0п���}Y���6@����P���/��k+$�y��i+|���Kd���'db�6T�u�ŒK���O���BTd��0Ops�Θ'�a��yHA�Е4�a�(�nk^%�7��֝�J�a�:U�&3>}�:�e�n,YmTr�)���9��_�'���OU�@��V�ٮ���1f������9tG��o�IӪR�+ؐM�����[-X�X��!ߍ	��l��V���b��.��T��z{!�ꃃ�q@:|��.�����K~�C6��E����Ч���=)	�^���;�x�	��d$&7�<;4�*����`˷O,�/�V����R���m��i��xGTA�¶&����IV�X!A��(��g1�p�
9Tdy�n�	��1�h!Z���+�c��֗���_��1`SQ��^Tq�^[\�!�>�5ڴ�����xyP0��*�&U���I�� 3{8�|���ӷy]-�LP �QȨ<fr��K͸�ƮXx�`f��I�#�d�15X�Yn�c"E!��:�Ró�!D?� ���ț�tx/�a�SJ�{�������A>vgZK%��|U��K�H4���b͸b)k�ԋd��v�h�kO���ݗ68m�h��C��]�l�Z��uoSg@��Y��zd�-��x��;�7���n�"���z0����ްѮKW>�Y���,����ئd+�T�&�|
3�WIX�a�mCg�g}�qz+53�$/�ί����^Ŋ��Z�Ul~QNY7�g��v;X/��uH��9�/!E�����u��|������zX�F����� =� �Sx�u+��0O���ړ��J\r���h���O|�|�Kum�cp�������"sA�|f��^�M�-�_�"l�x�/A���4��uZ˞h[v�H��qR�ku���:�n�l^G%XK;���4��}�3A�4?+ZW�!%z��E��8�/U'/�6��v�$�^��#4'E3�a�`"��c~��#�2e(_
�� ���'�� 6��B5�[�3��{.��~܅C����W�R_�L�1�)�M뷂��ӫ�1�[ճ����4bS��V˥����9��VW���-s�� rS&6�VĨ�<<�[�r����ܣ�ISo�k�N>�t�k�h2R��P\<�i�{��a���V��z�Wf,���b&�Fĵ�;��.H��2���'9D�����d,���ő�kC��n��H,�"#]g9&_7/.f[���9\�s��0i�/��X�%�������:?�H���*-��_�;y���IC��-�o���B�sm;�]�x�߅��,.d�x���*m�W࿢�ؓ��Ky�M�iM�Y��e�X�� =\����vOvNl6ί�M[����>8�����Z��,;�v�^J�(n���gG`�"J�|�"��h����k  �F�\��*u����%m��rF�6*�cA�u����N�{�p4D����7$}�
�$�w��eR��F_�c{2>%#�q���6��ڔF/�->�_Y2��N��F��3� �ދ%��{��&ꁌY���z�k���T��O��e�"�,��# o��D���'�G&s�O�þ��4Tr��`=�|l��N��d�ϻ�\Y�j�uj7�x<���~I\�CbI���ԳX�iS�X�W�>*;(�IkE��qE�b�X��ӵz���B���=�����r��z�*ֱ��o��'ݾ�qL��!�Y�
���غ�w��W\����E��/6���h?x:d(v�iS�q��k�,ҫ�ِ|=>ce�Y	�7�U`� 2Z�0���A���]��AJ�2
`�.%�UK/��CԼNi��C��s'���yᆈ�룂�X�����U�z����g!z�N��iQ�K�7�\����rpX�C��Q+�I˃���`�&H��Q�_��Ճ�G��v�e�\���7?J��BQ<�3�Ƕu��ZJw��)�ib
w酼���;T������w��&~Z���E�1b��3iz��7���?D�4�d�zC#��oid0h�Lq���.x�����"��E41�o��fP ��w ��=���!�l,3�P���\@�����*a?�(A��Ĥ�BT��_�`��}�VY��1d����)���aHF�j�/HK�u����8q7����wC買E$�$�*P�tuFQ�܀�y���]�]l���Bd��f9�͊����ݢ5<u*�,����뗘׹ *j��$+A1����ݢ���K�-$}�د�=K��!/x��[��p��Z�]G@<��Sd�ʕ����f̋m�)x��<D{m�Nz����.�l�����Zۡ��l*�2�N�N3�!N�"�<%��T�3�י�[}Ң�������Nn�D�/%
��r"��� �����6D�^ �h.z��U!�))�N�+o�?�;�E�b�S�m�6H���{oJ]b�JH���,��[F��v�aK��o1��X����'�5	5n��ߥpx_ܹ�-�PS��z���������3ޮ�B�� �a��A����4@�Y���ag�[F��3��j*��8��J�.{�U%�}�B&���У�lj�݀2����V�$B�q��I��'+��o���9"20�;z�׃,�����j_�_V�3���� g��7���?m����X��2�&BP.����m�~0�|�oF�òQ71���C������&�8��KY�U�ו�>��8����+"��ӳu�OM����݃HaTu���5��%,��/iy�����^�Q�^��w �GZ<�Vhy
�	��cWCk-m��9���-�h��$i`�~�ة<C/��a!��XQ{�9�I%�v��{�j�Af��w�Me���W�ߋ5��N�i�w�8����D�_@��UѤ�5��o�l��L��Z0�u��Dsj�4ß�4*�vs�(��+�r���k��!�Aᗱr;�lS&����6���w��YE$��QH�-v$�&mxg��k`
`1�\�~E�u*ơ�N��0O�����Oh��=`����	���5~����o�ckZ���V�RnѠe`���Yc�O7�!�	��l7��	(�	v�8�b��g ���,�/���4�ͽ�����U5�@n��{je��8�/)��q�m&��ҕT%��e�A�:4DYDUr(*���8<�┮��#�f�0{�����=�t�߸��6)�� ���L���E^���5!dc `\�vs�=A�AZ��Ɂ�E�_�`xHS�I6~d�p-��c3Qe�a{qVi0�O�_�'��i��XD|�T�O_Li�"}����R#�]��I�&��:y��y���]qxF��H�Vm��K��j�Z�n7��ۍ#2�������ڡ��-��/��I���=0�)���S���~��9*7��9�ט�t�2T�7"h ��n���>���������^�%����!��w�K��W7e?���^~�z���<�2o�9Ih5���3Q<�4�N�^YsH��{x�>���u��ZbB�}�VY1�1���ԇ�B�u'.i��xx���	�����¸W�g}��6�V������ˤ���0�K�1�?,qn��r�`~_�r,۟�YXH�ə�V	�I33�=D;h��*|;I��*3r+���YQ�g����� �����9Q��[f�^́�@:��1�jdy�e�Ŀ�%-���F�1�c���}�: qϸ��MsKn��)��xM���� ·,���o��L���6�ѻ6��� 1#8wSR@v$�uE����d�B+
kXm���y� e�(G��m���8�_m��e�r�hN�6_M�K��j�&��O_�QG<���j����.�5p�+���v5	gy `��}ן����D���?��aN�e&��L"��{W�����O�ҿSڜs�U_�����֐�m�p�l��+^�x'иkTf`���i}U/����Y���n��h^uO| �O1\?�a�vU�;g�b�4�����0
��0��_���A�T��M���ҹ�	C&�l��Y2� ��C��\[�;���ȗ-��4P0����g2fjX�7��?i�mK7����H+��(�Ӊ�����Ui���V������:��m�?����:N����C�:�kM�_�.���K.��~�!����w�A�%E��'k����m����S3�ܭj��V��oD6�[5��dvY�CI�ڋ�Hco5@XN�\2SuxڗM�>�?��!�
�/z�hr��d�5ot9����m&�WF@@t�B�uU��X���/a��>����XD��d�-�r��g��9�{rd2�!]i��B�q���dq�`Σ$�gÈX*���S���>-�>�@c��&�""�ة�V�]�*���hn��^b�a�;�/��m��)|}SA
��!�������*1��V
�T���>���ovq[�� B;�=���eB��<�,Zq��y"
�M}Dݙ��&�k�s4�p���ϣYXq�� 4���*�[�
\v����$N3�D��^�A���/_#�kY�g�m^6G��c��9_�x�%w@
�N��B�._,�&{�w�����h`o@������[��f�mJ�7���)�Wn�	ٲ�e~����&�	�KDl��lS��y���L��Bn�*􂓇;�Y�c�t�,��^�����'dt����r�u����C�a��ʒ(��Y��?c�:'�d��%Ռ�`�;��\g�SR�:sYln&��3�S�K�.'vP�Pޙ�/ի�??�r���Lr���j&��~F�-�wz�&�hQ	 a�^�$±��O�W��H'�����_[	��U�E���8hg=O�K8F�{�A��ˏ�Z�\=|��K�mZA��)('�����¶CQ��H]�۫|��"o]����hd����0�8
�U��Ӓ>��?),Ġ!���K���FNg	o��O������m�˵e�U[�m�vkٶm��-�kY˾O�}��=չ^z�:�9Gs0D�E1��@�g�+4.W�~r�sZ����>Ն�d��g84��(*]᫉������;<�����Dj�n�ƛ�&N(�*�X�+�z����ƥ�\>�{�_�bF-*��\c��fCȄ�'��FXY���1��s��[C���~�Z&�Y^f�̷��{��?$�A�����L@�)iY�}O�63ZUX���̌m�Ew�`/Ik��.F
ՉEo>�&�^�E�f��S�����çG5����DnA-eU�%���-�v���ݏ�)4��?ٷ+���ߗe~W��!�/x�zP��}���u,��~8aBC8�L��
g�5�+~��H��_X����G�`_=n<Ul��m�H�����P��g��-\�
�<�\���x��Z<���fcp����"�4�|�祿Z+a���gA���Z3�zzZxW��]�J6��Ǭf���S/���-2O�|L^�p�b�?Y�:��"�._0�_9m�9���>�L%�<I�?m� %�6Myi���i��Ԁi�|-�}����,��Y]����_�Χ��ո����-�^��[��U��K�-Y�����-��-ְ��yL�,�6�x�P�MͻFb�ot�).����G\ 0hR����;�����!��
����S�Yl��Ud�X�'o69+0
�ۻ��?߰��������O}_
�U1m�r햔Oa^׀�]�*O@��-�TF'������*���7�AY��;p��\�7�e��i]g%�G�(n�l�$�䍈�;u6���oN{h[ybca���U���%陳P�G�h+��HS$�B��l6��a�~�����3e	��z���)`]��!��}Ux�0^�q�E�\�k�:4ʻ"����KV� w|0�z��΁��m�?��*�Mk��Zm���\�c�w�,QgH��^O���ɚ��aJ���V���Ub���eQW4��S+������59���p�jl���E���|gZ`{��E�����GY�A
�H6����?�]h1���>��?ܸ=�ݢ��E0�۷�iR�X�-[�>�%�E!4��b�B����n�a����u���],�&�k�^�E:0̚�%�Oj�H3����S�1Ҹ����B����p'�`y�ϧ�������pw�K�y�(��"5�I���>��=AX��;��o��̤�M�i)�8T<��{Ж���u�)��`���юrB��N�p�ݺ���e����p����=J�ix�'�{۫v	�V7��&�7�ٲ��ʿ�٩���H\�0�Q%�SP���f�)��ĂG.�|�ف߂B���&��=�<2�ao�o�O������dM�O�a�^^=v��4~����Lu��T���1vE�\�[ӓ�˽+{�m�t!��Ҭ`��-`����/����#s���%�o��z,O��p6}�O���]$ݟ��n�B�W�T�~M�����0PYdj�Q���LSz\�<.8�*nՆ"��qUd�f�%�%s��5ͷ�ލ�J��x�a{z���݈�ݞ�Tm=g�r+1ߘ���%�ٿ.��%�՟���ӡy=�j��Iu\쾨�'�LW���AE.��`��n�	�S	�NFWq��2Ԅ;���`���T��r���3��L"v;e�Z����:S�mM���,Q�VF�i�u��Q� �;�R5%�e���8��m*L̩�~4��j�y��=�^�Պe�_I��O�?��6�a�f¤�����"8
���GA�է�C��uAu���x/�u�$$~#��6|���e�������b&��A	KxQd4(����'���j�3�b��`��)]�0R(�����_�Rq�*��sn��|~h]o����}���=u�-�b)��w��;)��c^R2�kv��3��0:���]@r/���ˀ�e�Ĳ&nEWnyDf�!�4żZ`�CYk`! @����3/��퓦��Z<Mވ�Y� N�=��5�M�f�Z-c��O�7n�n��P8���I���Bl�~�zG/�d�+q���y�r�{��v���e���
J���F߮ұؾr^JVL��h��;�-��ҟc��ҁ�
�%��$���,�=>b�f���nY���t�`��l8/����O��w	#� %����Иa��Y�VS)u�������U�3,A�ʵ�	��B�>�b_'�'�A�Xx��_��Q��.��Z�$�-�|Q_�X�ތv��r�~��&��.� �������QƼ��e!Էxz��f�[�0�9�[.,`j�B��1
���v�l���z��h���hٔ����꫚�t�^�s��&���'oK��#z�^[篴�|�;��$�&��=��g�*�Ztu�QBU��bM���lI�� m���Q��}So�6!��_�����v�N�Y'�6�(�E�B&W�Z�ya�Ju$��e�
�H��1�D'�+v
_�3^��Z����r�u}�J�r�>�v31y+8�pA��Y�1���}�A��B� [�~*��⿁����Q�j�#����U��ϳ���2����)})��Zѣ	������	��Ż�4媛��l�h�<4ҕ��Ȫ[�����q�5��,ק�Xr��٥������go���:����mE���,5�>X�{��l���������� ةn�q��Y��9�X=R�o��y�y>\r�)�C�H���d�w��N�.�[�<�0�����t�0c��}��ke�ݗ8n�f�(�.�|(ȢӞ��^K�0���u�J"�}��pR�m�#�l�5���~Y��`�k7�d�mǠ�r�^��hC�p)!�e�}q�a~?��_�T�↘�ɍCK�L(��l0�hc�YF��I�Cz�v4FM���"�]�K�Bɟ{2�!XP��9�Ӛ^�x�a~���&Z�����^0��.����<b~[EQo@VBsn�h����*�l`���i��Ĵ`8<�i��Y��x��SĚ$�n��fA�RRW���<ha����/�J#l��]�F�Լ������7�F�\���[��*�Y7��_:T�nX謡�c!�z<Ol��D�S���N�a��o���x�jV| ���c�:��A7���Ô��/�j�Ę�	$�G�O�;��,�ɻ�3�g�ˋn�U�I�?��u:�n�Ѻ����v�}}{Ȑ�͉���S:�`�[�h@�>�q�P��8b><O~Gnj��M}���N���n��m�mzA�I8��,�,�[/`�:jH��~,��X3#k�v�z�q���*\�X>aȴ�3�n���ފ& �#:���,��zt�&�0Ѩ���.���֌.H��od�^5�fŔVz?�G|�v�,P��4M+�W��㭹��8;�b#x?Ƽ�h������py�.�V���S!�[W��,�J���7�Zo�n�<0[�6�����L%`E��	�&�={�������������H�����g�J�Z����������#�o�����u �r��"^w�5k֐{>w��}h#_Q8W~9t���1FK[^��Z�e���Q3��[��A?�#�"���%ڝ&r��SoM*�� ���`x����8��-���ti���W�806�5t=��i���V��y�'��J���u��"ʿ�W��3z�r
C�I]!���9���=uK�b#��i#�N��G��H�\�4���.����<����a��Z��[@.A��M��n�脄��|~����vm	
ZG�,yI$��X3lH��b�-qo��g�%��v�}�Sw���pgꞒ���o��}�,�wh�}���.�ʐལY
F��&��w"��馒%t-C�>ӊ��$EV��#���\�Jy�5�T0Q��Ҕ�w����mʨ����_����b��$���9-���``}�q�����oF����=g��*?�"O�����[,�g��L!�z�6r�'"��rO�x����˚��o���ׅ�>��f�cmL�����UC��z���}�Y�k�j��(v������IM�I���x�?ڼ[�*2%�Q�vGx�m�U�Ԥ�ۈO�\�G�:�U���F�x���V��	&|bJVWձq�\�z1���bЪ�c��N"1]��jH�a�'����gl_�!F���C�^K���+j7>�Ē��3��ve��8I��g��+=(b\rGv�nձ��aS+�ex�f��z{@U�_��(��E�g���'(\��-��(k�Vy�D4Dc��Y�W�c%���/Oݙ��sqɨ���&���� 	N�=pB�ޚ���%7���[���U�����e�<���j&f���0/�|5�F.H}Rf��Z����Y�r.b�g)�P�Q�Q��|K?�P⍭B�eT&�kBHRg�+��6��Q�>�������,�Q��`d`���!p���%{F���z����K��)3J����O3R��5��˵]Ī����j�� ����Ҫa�<�E�v���f�%��AKKa��J;��cg %=��`X�#X�����l�IzK�T�S�ҊY�P����%	���Q��3y��(�LOIʭ�T��V2H�}w��V͘�*\S�>m?�X��
^�6c����Z�[cH�3E唥܂9��r�J��&H��Iu+�
>��yj6B���6���}.Jf�j���T��_�?�1'q��_i}�?�QfYU;���
4/<e�9����+�aۊ���q��
/i|)G]e)�C+�^خZ�"��SS`}�䕉�������U�2y=�y�.�xmx0�x��8�c5[��Ț ��'��i~�������BvS���6�ي}�`�bA�6�"
�F�5��ms�H-k�/��99�d�ܔ)UO����]�ؤ88�痼����3�� ��^'��>�`h:��Y g=��l�F�b��G�}V�=�䅸��<��uD�pYP`��bo�J-��;I+����������]�%y dMv�^���o��K��o*�)���j2&G�4�"��3H"h8�fT-���B<:�����^N_״�Xe{X�׭�]����xb�WL��>��;*iux/<k��c�BF/���Ē���&.�Y1tm/R�*;[T�_��
tA@�ZjYrcU+�]��!%�89�(���d�r�^a���	$5:�S���g>��p����N� �Zg�����Ji���hD����m;O2���6�K�U0(:�a�47`�El)��K��v���ex@X3FE_σ�g������PA˸'�9`�&�?>�S��L{�\�<k��?=�1/G`�Й\��N�N�S΃��I�Ove5���02-�9%�am�U��I7���[�\1��?��!�9� �,������vQ[�H	c�w?7�{�!���� i��������[��?��ȓ��[q)�����B��9oc{Sw$2Z(��'�kG͂���H���嬣���>��
�_�j0���t>VQ�j��{�3�i����
~��e�i~��г�iR��_ΒF��CN$��К��)k�F@j3[rK��s���ڧvA#|'�ϫ�/V��y����*p9$�u��Ή���v�<���0�1�TF�sCP*P9�	���&���&g��P�O�gZmɏ8��P��\���e`[���)_D�iK��B�j�?�~ͷ{�ƍ#�ao��o�;��o�����n���(�HAIy�vJ��RGФ#��^Y�)�S� ��J��&���M����6�O�|���y�i��Z]����d�%�]��6C�H5���!����0C��Ϡ��F�1�G!ۤֆ@S�]A�9M�JĿT�?ܴ��Դ�yR&+�e��G��C�߻VatІ[R���'X��}����*4�|k� �y���glp�>F�(xp��s[/"�����3<��5W��k�����0�y���H�5VJd^��ҙ���h���f�>�����H���ٹ��AI��z�H�����]�5��X	��	�TOEImV�� ^
�h������k���Z,3�J�d�L��z�[����N������_�����@�<�ͱK��Iۍ�L�%��Zs	��њg�8�׶d�&`q���K�I"y���.�;q�M�<l���T��S��IZ�S�i�� aW��u��ߘ�7[�:��)�.���3DmZK���0M衶SB턹�L�g�/�̐Z�*ư"w�ta\2Ch3iW��nWv�Q�L������"f5O?N�������q��� �`a�V.Ă����@4����?�FQı�4N��3��t��՜��[�hED�����0�k��ֳ��n�m��"E���_ey�q-�0�sC Q���:�"��o�h9%4��C<�����/�G��(�I��-�����{����BM�=y�]��`a������j`�b���0�
o�ÊK-ƳJF���f�M�c7�ˮgT+}ۤ.<^?T�Oz.-)�P�n�R$�U$�:��1������=Ex��M7��Y��7gQ�*��#5W��X�x��u�9�вV����h�tNR��f�(Ko¾��ަ����t��ҋ��
ҏ�	���Ui�6m��GB���ܽa�O��=`Ug�zow�[|�x��ț3D����.>dt���c�%rWr��z�'��:Q��E��%/~�Hy�jIZu��^
vqc���P�>� �tQ~�� ��3�5Ī�m(���D4YII958a�ڍ�W��^���k��%9�Gɇ�����CWܗ�+!$0�,�w5a�E�/��hÙ��b�sg2�~k�B����~���m_md�oL��xM���y3`�|S�����&�����W���dV��k
��߹~3�����@g�{���F�j��V8뽾-�5���WƂ�B�j��{��"�>ܥ���;�����g0Y�y�l��ݦ�D���ߔ�n#�����:���V�
#�p�56��y	�֭G��z�'��8���*y���!����Z���0TjPNh�-�e1в���/@%UX�?� =�hB�ë��)��h�V��mC��>�i�fd�X��K/�Ii�-M�+�����O}���ZV�]�\�p������n��1�����@�h�D���l]82'J��wԲ;;S�iS�}��x��܆/Y�~H`m���Z��V�?-PD%��Jz¨��\���?me.�������J��P���h1�0Ļ(��IL�vJE�x}Wi>L���NW����P����"��K�����w~[���nQK�ĭ��؀�u���Vdl���X~��ic^��q���U���*�&r��*��i]Qp�)����2���#o�Ҵn#����Þ�G^@J�bF�BUz7N1�v����$��B�'P� G(���%�貸�aW��Ìv�-�8�bΔ�E����D4���x����$sZ�' mjD������]d,GH$�X}���J����Z`dR�(9�Ղ�|�Şk;DY��-p�����ќ���b��s�Ĉ/u=�IH��7�����G��:f�!ePr�9ժ�}Z��WK�v{C��M]Q����t}SO�'����_v��3�;@�lI|�dUO@�կ��XO�\����)w\��_��)R+0���w^X���}:8�-fbr7��wE<�7n���<+.�ul�#�^��C'ۺζ�8b���1�A���9��~o�>��}�^�w��F.�q��[d�*�7|��� B�~��5��"�;Z2��@J�ĊyAt��e�zOZa�
�3�:�Y���\BB9��]I�V$�/�D3~	ms�?Ȯ������6�<}���;��!C@D`�ޢ��;Dd�U���J��aF�����W��w̱�q��i�Yү����jy�l& ON��2+�9$��V;[�����$���y��X��B&��-}tA=�cy�&4��<RE��!��@.��nsG�6��}�����Zn3|��U=��=�]�A�sd���)[���	��7ػu�Xu��d�9���s�{���qF�N�l�d�ҢL��W ���߆���D�:xP��-���u�s��i���s�������%��h�>��>o���*����_k㛐���G$�[s��Ew<.�0�i��=�'��<�N�k�u��#}�@�.��ʪ˗��NUҋ�'��je�ᷬ=d��Z�����y��a��fL@K+�x"x`���,#����Zi����g��RÎ��IX�{�|�[���5�$��(,��27�ob���/}Nҿ�	�����32ɫc�U�A ��d��!���}�K{��od���䇛4*��0��������[��)�0�ؤ���ue��L��x�m��?'g�4��m�����E�A0)�]��v�,2�`��V#d����}�����YgB��ħs��0��r�ҫW/^�[���Ũ����'[9Bn�Ӄ)h�΁��O�i��~sމ%�bǡ��g-S,8}{vv˨��q��&��_G ��$���o1+�K���\L�+eX܆b�<E	���6�}���9I��h8�FiJ��ie�oiW��:R��⧋��u����ݦ��3uI=j���]��ΙI)���(2���8��\n���>�\��粝��R�8�83�qr�)��m�E���±�R�N$���_p������x��r]��r���nS��p�MR�#�<�&�b�����J����l�u���^؇I�WĦ�+K�c���]��u�!��?��a/�OLA=]k�k-�\�D�d�X���U�����r(V\	a	r��ݷ����&��Akݟ(O�%��o����7ˬ��9v�^Dgn�3�D>�s~���|��G�k~���]G,���*�k��_����?��ݧ�0�0x��䱱UI��rڿ��y���yݺ����)�B1��_���}���xra��'V�J���/QohYv�N��	O�F0��]b
���EZ�]b_V
�^S��Bj�kx��^�p���/��\�ܯ�p��1��h7���j�͂a��������U-�f�����%��,\u��z�u�N:j�Wz�\�y"�P]O� b�p;��q�`�#�:Ss��
=��Z��~ѱ�2��`,in�hYo��*�nĐGNC�>��/N��d8�q�$Q$�;�6�w�������j6�
V7�O�\=+�8_�����W
�F�;��< ��2X��	�ר)�L=�R�;��F���(~�W5��.Qb]]\a�۷&�����+V��L^�u�Ak|�֟G�H�.d?�\R�
�M�'N�
�o.�b,UY5zN�����&Ş�	Y�H�lb����#��:�b�/\�G& �!w-z&�e�u�q�?+��p0�Tu��
���vd*�@���.�W�N
u����b����F�K�7���'�e�q����g{���k�@�~�ފ��R=���1@�~M��@����{�U�%8�=:8<8�J���[�OP�ߖ92dd�^�-N$h���j��
�l.��ٕd-oh�l0����K�kj�uk��^���/>�]���7���Zx�!#��
��;B�x>���.	�*�}17�{���\����ۋ]?�Q�iJ>�A
idpg���'cF
�.����k����Py��M>&����^�HU��g��_�1q�K�s�h}) B��k��f�U��T�<�b`}5����͞T|Ĳ�f�%Ef��J S*��`�n�@����t�������W}B4���U��ҷ��k�N��S������`!^�(9%������Z_;^,??~��vF�#;3V���j�FS�uzVT)���I`M%�]��#���u���m9_1+��\.说��lN<v+���s�b�TB�����MSxV��^��J�����.�t�n��Hˬ	!�ĕ�+tڭ�� ���CV�h�b�����ÞJK���[�a/1��0:����֟�_R,�#k;��s+�V�����>��e��/�'~���B�}�8j��#���v���V�f^(=gM�[H��0u��}�P��z��v6:�iL��lm�� �.^H�/��玻hB��0����H�K�У��<�ѱ�z�B���wEb�n�~����)0 ��IY�Z1�]������6fȸJ�Lţ������xP(�T�H�{^�ȥ�ӧ�C6D���򥟕��R{�Y<��p:M�j����#u_>a;�-�oKj��r�Z�������r��λ�g�JRbM��l��];&,��#.{S�}Q�;"?�s� 5}s�<EGC�_O9��!MN��L��!S��/S��e˞[�s_oMp�4�WEAwב�Y�t�t��h�w��,Bu��Є�H6����w��CܞF�qe�?|����_3�Qw�Jku��,�;3TkiF	[vF�i�f[<>��zm��(Av|���I�F��g�P��@�ƾ;���D
�r����k�}	./]^�L��c7#��&/�"�$#?���rWę���	h���&E�鰱弟p��<��D���:L���@-3��������}'�`�FŔ�ͰP�﹂�=o�)�o�R��z<Z�Y$����px+Mvl�o���}R��bS�$t���ON?�8�{#ۓ�r��s�](5��O�.��)؊����[3�����C�G,'����L��~ɶ_z�U%�x���#"_�V�f�8�	�rl]V�_\��/��8TH!X�D���y4��أd�#/멺�W�{�g�����ܷS�_1�L����Vhh6��� 7D����%����fI��RI�t𕯟>{`(I\�@w���q�bI�U�\�n�㍔f��( ����S����.G�m`�Z�ki�����X�=G29q�.��jgM=zj4xEV�y�
��%_��}��T��������©��f��q�����ޤ`���<��DcJ����S��π�����)+�9A�d[4J�đ�O��X�3О�j�Ź��Ms�j�j�׋�/�<��ƤY`��6��XZ��T��;�G�^s3ԧ,�	��8pdAq]b��� ���&�o�ql�_(�ٍz%�K��;v]����1 �~$-X��[�႖��#KgOW-���z�Q�`���
b��V�Zd`b���gj��I�_c��ۧ�|�B������R��U[+P�d�Ã�h!_<��B����+�����p���"�,��~������
��E����<��g��	��՟Ļ�0& �ic����1w@�ܗ����҄9�;��d����=�G�|��LM�u�8g^?����u0B�����2�xn�.�������ggk�P`W��~�Ǵ;��"܊?޽ةa*=F+C��y������Om#�A�E,�-��p��ĸ��4�R(���`�F �o73��P�v�`Đ�����VU'��L�i`q!:,�E��w�o~����c��u�?���q�|Mݵ�HL�A��@T7H�N��p��#U�H��}C 	2�a����zc����8T_��P/�q�����þ7��+b�`Xg�Zx8�}�V<1�o_�$�AG-QP~?9�-��ѐ�!v� &���$-&J��?�mq8�+{D���_BO���W�h�AJ@s�}s6YWtI�h$3;5j6�����̌��^�~�s�S�7n���Y��A��ՌDA�U�Ɵ���C��%��`�ʏIk���� �?*����T~2%H.]�ˋpO�VH	P$V��O�8y#��P��5�:�NH�Q^�B&���ޙ��_�fC���EY�f�B�-�Z^&0��2��!�^�DJ	H�f8�s,K���J����v�#z���-�2�6�˾R^���Ho_?�C0%MD$pR����
�^�W��ݝ�u\��dR��!�����߳�0��<�*,�8���^���u�d]�Ǐݑ�Db��Tfj-#��V�/y�H9�m�]ī-��f��!�W�׵9�>n�$�������_Ţp�t3��%�y�Ϯ�~6�~(�
����Q�4W�v�H.�v�<��Z��&&Oe���e�
�=�p7^��&*e!'C�8&ְ���A�k��
ў��۱��$8�;G��7/FHMϾCAX�*���
�J��7��J �m���TU��:k�Oi2�DbC�<߯��o�z�ԫ���v�?`�"$�t�_�ִ�j��o�^��/�ŀ~h"��3u��`f���~��>*a��r��zN��6�^�u??g�2�)O��ӂE]����zP��6Y��R���<}��B��]F��\b�W�I��7��s�%|�&ܶ��7�|˺7������K`��\t��#�3g�VLr��Ϗ
QE���i$��V%���$��"��5�&ۓɢz��Ӈ�~����We$���.�}%�F�T����y::���ѩ�E� ���7����Ɵ�FI�/R��rBB����?�=��m8�J�MƤ�7D�����p�R��l)����ϫ����4F�����X� �������N9D3~��Z��p�H�+}^�
i���DZ1�͕D���3�n�qmv5���<JʠQ�NB\9쎆\�)�/TF�x�G�SꓣV��oʝN��*g�.#Т���p}��ة������;0�aW��rc$�����Ӓ��ǩo>�<�M��H��wv6�]e����8����r�
�FFn��)�ޘ�@3xh[WZ�YQ"X؝Y{s}�[���|�Yj)[�ys�Q&��+֕��MV_��j�`	�#�`V��؈v��������Y *�
��fT��>*�E��`��V�)�Vc�Ė֯Bi�d=~�Ѷ��y.j#�H���qЬu�9�*�� }�g���<�"
:!Ǔ��$�P�W5�w��A�8Ip�ZD>���F�-�(�����綢��`���R�
U�L:1���)��V�b�=���j{�9l�ak\�#����i2Ԗޡ#V���������T}��-(`���x������pUNlñZ�C��j�X�)��aT��J�`(D-/��Ò�1����D��t��Zj�:
 R�c�vP���l�o�v7��E�gу� W�w\oh������Ŝ�b���z�aP�d�ؠ����W5��R0":�?���[#+S��zem%�#��;)W�����Ux��V�DId���1~���KSP��p��՚P�
2�*����`Y��^��]��a�fw�dN��cu�)�6@cڑ��Qyux<��9�'����;u{kf�jl���<GDh���P��p��-�[��E�#u�+ڨƭp8h69]q%��2�?7�F��b�Iu?����J��������F���L������������	{�n��#v�Q���������oЁ����ἶ#z{�)����QaF>�ZͶ���k��S?��q�hId�_�27�z�DalM��vf��ͦ�sN�ې��x������{���>h���b��X�{�<��b;�t+��8�-��q"� �s�T���
���uF�{/S���5����X�Zb��~#���"FUo&�*���C�B��`ъK7���_�~�|>2�.�|�]w��?�� �ӥ��b���rV����dY��������6�����nO��V1�����.})��\�����!L��ó-#��b���+��"������@�hv�K�EIN���EYl��7w���}0�c��b~�h<�˧	_=Dz��$�����g����%c0�i��c�ju��fѬ 4 ��C#"�_ ��&�����ܦY�W�L�����������-�����g��P���%C��$Y`s�"�����} ZVK���!g�D�2o7�8�B�W��&
~>����L�ȀN���%�<�c��bQ痪�D?Ӑ��A�zb`ݩ/ZU�*A��>uT���s����Ш���g�6�M§�dD���-���8�gW�T?T�����^��h�?(η������2�T�i�a�ֿ�ڷuO�c��+U������:���+�NT6�:�pP!���95m�0W�RS�֛�R���,d�0�$>�5�������9fL	�b�qi,Et���K@%,{g��!QҲ�1��{�Q� 붢«/�l�79�I�"�atžA*8J$qն��B��(4�rC*�J�����
�����O3�jqsdZ����)k.Ĉ��zr�;����N9z�t'.�1�
�nA�d@$�x���m�|�.=��祿| Q~a/���	J1�N6�?)� [����P�u�c����d�c)gjk��-0���ke�52Q?{:�g�b�B�.3j�m���T�/Fαީ��r��@f=���{!q�g>�r9�8ǝ��v����3h.-O��W!��
�!Ұ�5��;��3V1O�X6�WA*�G��/.:Z��*g̈́#W��\D�-(t�Pi�2f�� ��dB �%�&Oѻ'Zx�7��V��!<ML��O&t�ҥ�ˬ��/ ��"������N՛�;�0��TvN��V������j�,p�������&� B���\�g��kF6VN9���QV�8���,�&\Y�g��	KzC���K���oq�4�V�s�'�E�@ן 
�3֏���٩�V�&���I����a��6���[����(oҞ���Z�5p�����̏���� �ޜI�����|�T����@hu�	����<��Ʈp��.һ=}Κ?P��>�����F�/��P����M<9uDt��=�Q1r�:�R� ��޵yD !��Z*��ٖG;�Ǣu���&�e���Yu@Όy�V�v�Zg.�^�F�Γ��>�o_�ö�+�9�W���(vWľ>i2d�h�&����Ǣ_����q��&�k�g��P���C�ɀp�%l�w��~v[c������2;��N���U��x��ٽ�`z|C���;�����I��n�Hy2�Ө����{Ɍ���,��#���\���A�|o��~�N�ɢ:hF�U���rZ��l4��:F�/�a���6��N�`����V�yK�`��9��	O��N}�_ZT���c����O��)ح�ȟ�k�`��Z�*�H��
�'�,�&%B���c[e������w�aaqNu�_�9�{!��y�h�q��W�P�xw����l�����
�K�����v��q��=I �)����(PIȍ�c�R�U:��|W�AM|�*:8� ���;�.e�>��Jh_�[�5`N��W(�=o�jw�Tcw{Wt��Q����(�?H5���@#���h�b˳h7c�'d�#j�ݫ������Q�!��Q㷹���6�٩Wʭ�n��˥ �f���	(�ɒ�m!F�
q�OP�O�dّxϵ@��D�]��r{i�o�H�Z���y���r���c�#��|C-�Y�<1�D$aŽ�}ظ�5/��ʹ��q��W���p7�*O����
���Ϙ����&i-��������$�����8yd.��p0���o�"�D~���RXc����|���P�Żm�,�Жg��E#�?��Y��+|��?��Q� wZ~�5�4.��ā0qc-a!߳�a�"��B9w�������8S�
W�N�+�Xx���>98x/;���Y�M��Q���V��/*�IP_���,�%��n����`����3E���Wdq��'P��O���&ԷUEi��anL;����ۻ���ˬ6���]E�>Z���HK�u�G���?������Y��bW�;S�b�bV�G�f����13���+C~- ���´�1HY7Toml���r�2���䪉A18��6̞g��I�"�N-GN�?M�Ny�
��wt$�j�8��x�8T��%�R��_����c'5XEo�8_������k���a�f0���ر��S�H��JZ��H�#���0�<�<k��i�`/G�THB��4�9�NګZ�U�fr*w������sڴ�u*������`N�H���Պ��i����|([+��1ALEĈgH���F��wVX.�^r� ׌� -/HL4l��ȵ!����i��O�-�7|�ҥ[�[ b�����D^�rR"�U*ﵶ��6�����ҁF�F��`�$�r�I�^k&��	I�O����[V�f*~�/�Ce{uD����p�G��u�}"�N�Ϟs���!i�N}1�5���+�o	�����n`�v�"r���(�0�߹'d|�T�y|".��|�%�q�������N�B�QKF@���Pݵ��O䴨�(�k�ʡ
�Vy2�뎀���p@���5��6�h�F3�]�T��!�/5�ؓ�����NGh��h�c� /�{�P��o� �kh?�-f_�"F��]��������Y���E�������TH\Kc�6A%m�Q�g�ç���Q�C�7���O)F�QR�*��d���,8sJ'��3�ɉ,�C%?U̔�	�&����`k��DI���U���~0���;�aat���`LʱJ�f�*t"�;� z�	��B,�@���b=�3�ѩ�2�j4nb��@�	��/���sN9ʆ"�C���������{߀�$�f@@��F@Z@P����;	a �F�����A:�n�3|�����>�<.ed8{�{�q��u�Mu8�J��F�hlK8T�?&�{���bYԻ���� .�(\ԣ���|�A$���Z[>��/�6VF��H��`w1��-D�S���)��3mV�⵸8�v3�O�Y�}���ԅ��#w|��[Fܣ�_� �T����p�	�&�/��W���	 b�ٳ�Tek�"���Ziܣ3!G��ɉ� B]��z)3Zm3&�/dɻ��d�������ӋRt��(c�SX�8���R��0�]o��  LaSV��+C�j{WԐ�(�s��0�z��m��N�a�+\Y)"|Xr1�)`��1��u�������B!GX��t?��z�]��(���z����hisBF�:?b��R���|�^AI5�u,���dv5l����ư)����ҫ6�޾�1�c�W=UJ����%�i�c�
�L�X�����x��#�7�H]�DCf~nF�/]�8�m"�'�q2;@�����MAI��AM���%n������C�{�K�)������cp�ۓ>MtO/�o���c$�#���U+��jIS�H���>�yŹ�C}*
��T��]9m�� �5��|��[qm���P�+>�2����_/+�$ �*o)�Bp��Z�K	���=��������J~H��C�5�%��VCj��}�	%��H��pE� o/�2)6�q�H��Z����7���XF�JJQ��jb��o@��ӻ!��1ý]��N�B?�rv��ϗ����W�Ʊ�R�� 2��i��tph�8�e|�ZH���zԨ����᤺�n*�R��`��4��^L����������PYp� �B����W��s���^.�����#i6��ىRU��j��n�}�3��_X���Pβj8Т�V�C?�z"L��ߓ����SO�%�|�"vt� �%@�{}�6����� ���Z�bR��w�'V����/K��D�9��t���zK9�*Ȍ��,���>���$�^/���栖�0A49�i��:�!ˈp���P�z
2��7�uBhU�Ȉ N�d�y�1m}�s��ޒ\@��e�ph/$��	�"(N	8����k�)K�b�������Mė���4K�r�p)��}�?�|D��VF;�ЦdϘe��H�Cn�*U�)�ta�*�Г��3�z�+E�� O���_+���~b����X��6���W.	@�'w��i�:�9���]rQ�_���#4�c6v�,k��O���>Ġ�S�U��#��{<so����v2��G�A2S��<)N����5-ɘu��=b�{���0��Y'|���˃e��p��ח,]�
탁�>�hM�� ��;�b�#)5h���\�2\x����x�kq�"%ǎ[�����[̆a�y���1��s��FJ��:_A��;���Yw�N�R�5!�rq�XƑN.m��J�c��}6�v�*J�M�����q��y��^ݯ�v]B:����:�-S�j����еD_bY�N�4���QQ-|k�Nb�����~�����U����9��\\��#���%4����ߪ��-���b�Vp�,Rh���*縦Y\}��o���y%�G��:��{̞�Եq� �[����������˜���m�DAG}�9�~���t�E]�ք|XF�� ף%�8h�#�Rhx�N�x97)gsu��p��':�o?U��k�x�քݑ����Gӛ$��
*�T'��{�D띾O�|.Қc�\����vI�m�����v���"�M4,��שE��gw<�3��Ԙ��:�Y�M/�`_�V>6��=�#�P%�\�8��GX��/�Q6YhӋ�[�+ �z(p)x�~gB�-��$��G�k��!�8���X�z�u�|~��t�Nt@���>���yL�S�h',���#�~�)�^�?�6���a�!5�l%:'�V������	\/I�ֻ�[8]�h�f���y��D�ז��(@u1�~x��G�=�`f��ą����9!��ge�j�S��x�h����B��D�����qU�SF�o��\N�t���6��m%0S�~!�uU;O+vm֐x�X5�l3�d�|�B��]�0�Uo�wB�d|�χL�d���ټ�_��'��A6`<B�k(T�u�&T<ϳ~$Sū-F����ȇ\{=�X�e�s�T�j2Z�^ ��^���;^o�
�uNVܘ�fA��E����eo#|��7��P��x(�n�`�)� FR�*Sej���Ѽ$mȓ�*������ ϫ�GQ���A珹tʊ��rsT"}�6+4��~�+8#�ƵW{�J��!��H쑈�ǸӧC:���F�s+��xslç�T=�ɞ�71v�9�5�#G1�c8��6g�Z��Չ9�<�V�F��ݓ�ǗT�GM��sA�[%�[�,�&�Y����B�"�l}m�ѡex��mW�j�g�(���;���d�(�0��WfF�H�JO�\�l��.�y���2M�ȟ���w�~�ȥ>->C��H�������^ak���_/@��1����P�g~*��"uP��<�u`B�%������` ��`�ʻpK}�B#4���f>�����x�?��f��t���r�]%ڟ�w?'.�ÉINۏ��~�{]��`rN�6��L3�{�8��5=y6�|sDi��g�ݓ����Oߠ�Y.}l��c�l��=!�r- 8:|ʟEz�F�������@���`	��J����F���?���Z|�k��"2AvuОrݣ��@$1/k���'����hX�*�,� t�x�^������75TM�3B�	\?�<�FN��\�(&�s�2L`;[v�.+_�u�gw�o�dޭ48K�����y��d�7da�l��|��S�3��ʟ���#j=T��6��� Ox)*�+�$�N_�2����U�g�4]��X�S�ۖ0�P��.��rq�A'�4���\���L�#��L0
]͈����ap_f%��%R���o��u��c��2Pp�Շ`�,�e���
�&4��1&Cա�3�!Ma =�px%��)�47��f�&6��V�:%����7��t|�Q�_~F�E���Y'���
a��<�h��Ы!80{���:Gcr*����s�9*~��F�I��7���ոl��r�ƚ��ӳ���_V��-���$�ϲN;h�lr�V�EE����}��B'����������(4P��`�Y!k�8�
,�2��{�ЇV����q�IN�(�SիL� nR@FdQ~��D��Jȉ��䃰yw�zk��'��uBܶ.e�Ē���9��&��d�"�R ��;wf8�j.��M�E�:�S6�&?�t��od���ф��b{�	��X�gU�?��.���4;�	��#����X�Ƅ>{�t� X�/;p:϶.'��J:Ԥ��l��
��ć]-PϥS��n�c�����	��n����ѩ�����7�V�W:)W6YȲ~�i$t|wFN0��J�pרq��/J�O�l-�:�A�H��[m��Kp����
q?u��pP�O(�WP���N�� ��qZ�^��X:b!�����o���]$�~�����=[�+v����{�hg`Ct~Q��ݕ2;��b@���^{*�>��F��m5?��̥�g�����(+ֿ��f� >���b7��去a��8���DjDJ	 b6�ǜ�_.�?��"���y�H\m�����q��7�Д>9�������n�]@���D:�g�nF���^K�0�<�-X�����f;�=��WȰ7�G�B�Ų`ۖcc9,S�"�)�CғA�����h�Б��}��'D�u��U�T4�lH*�<aN��Z�̸�\�lI��S�C�� 6\W]5T@�<,�CL����s�S���1= Ռ}��S��_&���.���dj��v��"��h�I�5s��H�s������%+L���	�󕨬`�s���ߎ�u�zl����|�9g~>����"�}�1L��|��;�T��$��x��ex'#�� -Lq�b����i�;�pV����c>h�O��mo{om���%:H+��*H]#�@�u{<V�����U}���h~�n~�����Z[D*�|�����t�e v�j���}RHlк��Ժ�E���X�>���
)/��:�027���YU�0�IXWA���,��jt���Z�y+�l}u���(������9ԥT-���S;�rV$���t�!�ޖ_�=����f^��S(`�y���MR|R�,+Ӑ�j����p��o�͑RB����bv��������ߝ
pm?��oI��	ܭz���L?��M&�`��<����IĨK�H+���Y�G�6�=�X������+�mN1y���B��v�����S]��}/;ј�q-���#�	v��<e��	�
�פ]�XR9Oz�o~Z���uH�iPlwDx�㛳vn���ۥ�ꗅ3l>UQ5*�X ysֳ�� ����#���[�)Ert.BꩯB�����ח�=�_Q&���|�n��B���g��A�zv�y��2����)A�]��ژ�`m1{�����D6�3�yJ'���K�D����jO��l@>�Vձ)_�T�?O>ڐ�V�/;f4!gn边h)���j�F�OB.g�v��+�E�^I�{�+�����[ҲU�Ç���6�Br�R��]�PQ�����Rv�u�����'�^�����'��&W!)B|�s]1OBF�Y�B��v��Lnc6˾����"v�B*��5�����ܓ�޸��>�5��P_��Z��~[�oW��>fs��kT? ~���Pi3�jO������M�g'S��e��~�7��~E��o	�6NQ�����mH�V{5�d�0���>��׋�ť���� �8+��P�fT��|*��<���M"�H$n[�,�l���Ų�	ڐHOH��)>�]/�#��y#o�63WLL?i��jj�ڙ�v��ޕ��"���^n)�;��-��]fX��ޓ�m��2�6;>W�����鋪9uԣtav�E��%S�>�
N�C|M�h��������s��g�V/_���gv��_�w��̘|F$U��T��U��������^�,�{.�Eɴ�x���'�q1�p*[Z>�҇�������_\��o̼�o�։�4�E0ֽ�a�F���E¸�ag-�E�!3;%<,�
������T}B|1.�\���Vskק�G�F�b/�v^s既����r�|�(�:��r������!�?��+&c�UYz�ey��q=���-Z��W�������������S���On����( ��cGˮ���������>_"�#�a��)M�X��7��u��l�s/��9W7�Ͳ~�/%w�]���e!�I�6���=Րi�jr��<ܑ����}��]�'�O�}��Qi*�bð�E�IS{D�*;��\b���.ff�x딉��F�ے�jL{�+U+�I��i��) �Z=�+�fO��E��U���md��L��W@�8\���􅝲@���kN�iM8��/f�Ԕ�f���Ē�_蘣5X�щ`������үLT�5����]��Rv��S��1>7;����7ȷ6�̧xR8��x3��h'�M�D��ȭ|H���}iٝz�a U}4L:�D��H��?d��x����t��*�;�0�����k�C鵭�k���6�]�JџeX�<�{�w�m�`��/1L�B�5��K�\ �����t����V��+�'���qf=��8�#S�����f5n�GL���O5.Ht'0����|�.IY�1]�X�c�>�7q�e;y�bf"�����Z��7~󎽿���)��kB�����������]�д�������
vT��}��
�Y3�9�S�$/Bp�9��IM�C~Z�[T���))��q��go��<bb��;�l�d����"������qm�Ӎj����^�ơ:����Ɓ.���l��B�X�9憎��F�4��N/����'���<��� H`�b�d3&�1�d�°�F�b�<yPѳ��Vur�������?�6ì�d��u�����?ߏ譆'%�:'�Ǽ�%e_KE2���Aq��T���D�����.�~�Jz�'�v���,}����Y�u"�5�č�?�l@v\X{h��p�B.�2�`�䝍��{l !�}�����2��%��1$Vt�ЊZ.�ѿ�`�8eO:惺�T�bBǾ�>��PP�:��%.2��(C��j=���-n��a���Y@�Z��$E�߁�Z�:�O0̏��^�lg�W9T9<6nKi�8"��b.�h-������V� �9�@c�	R�YO�3�(��l#�\o	?[�OI)z	q�|P���1��XKd@P�M���y����o�T�mhE��~r1ID�8�q2��t��M�}�,���B���ڔ�.eE�F��FG�#o�ɠ��ɺ�AD4�ƼIV�Z�M%����<HN���)�J�7Ele@X.��V+�ʺ�x�`�R/�� ٷ�X�6��z|[�#z�w�G����p�)�d�Q@^�יc-1,Rǩ�������k��ȋ���mߨ�a�߿�����5zSs5mȩ�vS�|#�6�1��2u?$^���O�Ĉ���:��R}K�!�Ja�>%fz[T�4z`뱩����G����A�:����#�q��
}j� ^�:�`޸�$���/�y�˹̾|�w�vYv�5���ƀ�jr1a�E�pfs�#{�i���8�%�j��e��{ZJi�R�ޏ��ƽ���!��Q:�𩇱�#�I��gpC��|V�r���ʰ��\/������7�6�*�P)�63��Q�.��Ns��J$\יuVEy��-%6(��.@�޺[Q�p8��N�YBS�>��Br�ӥ�X��%�D{�.u� p��2f�6r6���m���H�-'G�:9=O�F�6�$ ੽��%U��M��@2�\{}/�d�RV�xo6�W�	�|�Ed@lh����1�xrS�C�S�Ǒ�������Wʘ1�D�ź���tO�:��E*����
�ʵ&�E��b��	@���6�Ej4��Kr�E�b��t�/��H�Gհ�h}�$.џfXM����!R��c/n�G�u���@��?h �a>a|�u�������J�;֒�i�!-�c7
�bME�g:�]���Y[��(�\t�����w%;uלEۜ9������3��OM�$���J܁ ����9!m�\�����ҫ�q�o�i`_����#���P�S	7%�R��s�3�k����'is���ےH?ySZ_�ѵ������S����q��������#c�]/�6��oE}�d/��s����B��c�,҉����G��wIF>���e2��~|�\\-�{�8�0s�w�����3䖑�(����%@z���j6�Y^���EAs�r�|���QJ~���]i�<�
�����|�9���7�C�����}>�[��Z�5�`��h�\�Z��C���E�s�?/,�
D�b�e�̚�P-�v�h묧B%]��D��u��K<@>͟��\�r)ӆ��;`�ݫ�f���n8��R�-Y�r:���)	��j�'@z�E}(�2��1	LkK���4*Z/���k�����63T�U@���8.'�.���+���u#�w��-֧6�Ɗ�)�R�*�A4+],Ŏ��.�W�/h��^��JƷi�B�I{�C}���VQې>Dx��s�I�ض������&I�Os��#w.Qgs��4sy�����n� �{�/�;2 ��y��uZ�T$�-��6���J��/c�Iޠ��֩���_�)	�-7����[��Ee�C� ����cy����O����kq���ֆg_؆��F�B�m�Rog�0k���O�HJ��E��[p"��J�-D Ul8�U?����0N�;7|�u|���6�]{���^���fMDs�*�)l��E� іj��| f�6�GMT���!ħ�]���wï8�5gF,�9H�b�O�$B޽o�!ͺm�u��,5�9Y�Lu�Lh�t_U�o�]���?��s^n��5�3~9����4@"J��B��/�)���O�b�z�c^�#q���L>��Gȍ^���־L3����i9�]�rq�Խ)[Ք�UU��e\�`H�105�#ac��v%�k�HA��?SB�r���k�P��I���#~��	��~�<֔�m���(1�a��Eؐ��!�/م>�W[r���f)"�?����Kq�h��x����N����M��X�.����)�qFWYRZ�|XE�/K�|�+�Q�}i���!�n��㇣�N]�M��`Z�*��<,�cM����Oݳl{�<�gK���F�4^�D#?=�S��s�c,]e��W0�D[�o[y�� �)�S_��Lmy�/Bc��%�S�D���SP�R��L1��&{�r1�{��y|]@��<���;Q�hD�������icWTV�_�WS:^~b��ameZVj�V6��I�y�=���'G{6麌$[3#O;�}9�4=��'��l�޶���8�.|Q��.�e��_Xmu+O��C����'X?EZ�#���Ӥ%1z��oo�Z3�=��Rh�<�چ�L���h8�L���pc6���:˲]4��ܪ�QC{��*����iV��l�OV��F�)�B���]\6?l��E~�C"| �/�.�-V�*�%S�1#K�����:D��M����]��2n>i�#x�!bܱ�b�җ�/mlZAf�:��u��;��GA���H���Zd�Pupe����[��� @��-fFB<�����(wL�r;i$>u�2������f0�1�̈�i��gS�p����?��pO'�M��vT�@ Z�Q���O�E�Fd�`W�~ǯ�d{Z:�Р��n�B��l'|��xy���Ql�'�K$�w���"m��7R���5}j��U�~e�q��ZEη����O%�ߋ�_���p6�?
���*�Jd���>ݼ cy�,�"�Z$����rט��~[K§?O9tϳ��&.�s 7L\#>щ៥�?_^��2*�4Ӎ��uzI�+�h��Y2�A�8Y��K��b�;�7�S�X��i1s�J+��+NW�|B��ޠ/�Cl�:w5�t�(,��.��ɮ�X�8�`�je��ߦ��ݧS�Ѵ��Q;�y�SMi#����:*��-�ޕ��]��΄���ۿF��$$ /���N��]��e�u��Gw�g7�=�U	��[-r�/"���nt��Z@Xx���_r��=EɀI ��y��2ͅ�����rc�/���v��Dj�,�x����Uz9�������� ����j;8d�U����hi.�l�J��X�;
��o]m���ugs�6��:*~��@�^���m?k�C�XTon`l�8q,�ɮA)L���ֆ��d�'�|F��vDO��]�&D�R�qhű�	��) �^�.E��2����k���[�ci����f�ۑ�,�Q�����ڈ���j����G?�Wvx�4��u�L����ߔ:�<k��e�h8��wL�N7����J��a�*F)��|�1�,)"nr7�"�	{����C;'����o�H�Y�o/�����E��B�˶m"ż��M�4�w�4'�HYa��6����3?D9����Xä��^;�/�U���ė��%ǫ�ƀ����_�ex^1�:�[�j�1ޭ�ۈy��{��hn�ʽ�_��e�yY0���~<n�oc���fQN)e�+�a4�c���2Spv���ĕ��!��jnB���lz�Q.}�Y�˝�TJ�P�?�������힟���5��y��'M������6���C�h�x4�X�8���t�M~{c!��!��CE�>��s�l�{g�-\�9��I�[,ܶ�/�?߽���f�����Yr��z��Q�]:������a�\����'�9�w�=:˵ouqd���Y|8���ο�9�М$�{�1=�~:��7:���*o�ibZ<��7�I�ԭ�����������W݄ܵs1��]n|�E⽿�.��_ͯD�4���]�HF)%��^����DA�[�&����W��o��~���Б;q��^�s��0�����՝�t�����CL--
n��Ƣ��=����/���u};���c�׹bW�7��Y8��씝W�������h%�R���Dڈf����u���ፅ�\����֧�U�����0Bz�Z���J�ų��{��^PҜ��EJ�Z1�z
D��<	������������jћ��Ճ�CGyb�;܈��Iϡ!ů��G�6�R.e�}h���7٣�>��?��|,����x��8b���{�QBHo�N���dC>��`EM���-V8���J�+�˚�ϪBvSy���F�mO�A�����/�[;D��ֻ��p���(�Yʩ%!�����/��f���OGEl���kܪ�gv5�5K&.����2/��g6����o�m�û��9�4���$������9�v����.��z;��D�����IB��F�8)Ǜ��m��>�t8H���/�fw}#w�WL�����6I������D
:�����D[ �D�ع�%�b��l�?LJg����<.K�I+#�}�ʎ�(��8�-�x��~)��n��p��Sm�\�@�7ׇ%7���K���j��ծφ[W5�N
>���,�?�9�Y�z�<�/�W���d��~{'է���5� W�BJǆ��hl���pk/��Z��eK|�sw3�tJ�<b�+����N6oa�gY/Q>S�XV�.%e{���ϣ͎�H�<a���Ǖ�U� /_x4�������V�˾ o6bZ����S"�X�����<�"��W?J�w:�����V��˵q*��h��(� ���d�@$Vp0�����T���̧τa����o��D�F��MI����f���A�mfv;��]'MƔh�C5�`�g��Nz��cY�=�nm��7��ZٺXÿyu�d�z3���y�i��ϰgk�us���W��Aj�ܢ�����r��[��mo� `�<P��Ar�u��*�"i��-��F��}m:2��p�d�k���ܬX|����XD&z����g������B����Tir�����~={q)y�9v@t��к�堕�z&�}���9ux��a��T�X�K[=����L�( �ź|߭���=������n/�5�;N�����}�|O���޻��$�E�
��«m'���ꦓ�)(iE�u��q��9�᠍q�����p��W����&�2��{�ǋG�/L �����y�Q����.�ۛ���dY���n������6yT��\d�6ړG'�݇z�VD�L'*�z�-z��ܼ�?X�ە�1���|��~k���X�!Zc��X0���X��h_�9��Bx���d��Q���Q���^f\mm`ֿ�Air�h�6��!�)��2Q��D�s���K�l=��n+���q<wi��g�P��B��q�w,}�	k�3yׂh�.:��O@Ͽ��SGmt����)�@�aP�vEAs'��hx��C̨^3�����J���Y�C�sXa�����˾��}Z3ɕ�N��HD�Cd�����C�Dʫ�Յ�N���9�~���q�[���B#Qo�&��m|蒿�N���so����~T��!`m���*+m�S����ҟWԹ��ầl��y�� ��n��O���<%3�ou�ԡN+�G q�OS:v�z�,�uq��_kNc�;�	�։�sQA���ŋ }�w?�8;7��x��)�O��q���mf�\�r�|-�O�*/k3�D�J7c��.�3���DG�����8���wW��jL�N;��:yH9|&�G����G�	nʏg��2W��Fϡ�'��>���;�D
|��|g�J�>}��4{3X�r���3�T��R���.�����-�_����s��o���/2.��Ny ���,��ݟ{J�z�6�Ғ��E��(�b��B(�`� V�E��mY��L� }��n@�aÄ5�g-%��ۓ+*�芮�n3�_%A�3W���Τu�S![$�7<d��Ȧ������,�;%��f�g�L�%�����
0�֗�,������顎���S�	ѵqo˾���ŉ�zN#=i{f���Ey�m��� �Fx�1�l�	�V��V��D�������+b0b����������Çݙ-��C�6"�Y��1��/��ū_��ܿo3_m/6ye�i�Cc��`�MzE�E��p�Ep�ѺE1���_�t{"��^�
�͊N�M�g�X�aꥩM������m����]l2�=��X�`(��m)(h� ����R�d�*�T��2!�M&��`�TU��Y�l54M���͉MP�BvP,���Q@�5fv��f��&�0��C�JI�9h:�NEd�dW	l��6[t�WSmBO:+��gNW�}����v
��ݜo���S���`q�+r�=�xATP�E���m�<�ԁn� 4��|�h��X� (	���~�D9��d|7��� �i�3��{��D�z�{���>�H���W���y�r�K�6Է��o1#�	f%���s�
=�
�k�?B�"%�7E#��z9�E�X�����>܍i����tt���dL�����Ӑ�7����n�����`���!U�%Y��b/�=�2���e�����L�~S�dAمRuČP6�ߵ�qP��|8St��w1�&s;HOW��Ļ���y]�7��k����E��Mu#��_�E��g�4v2q�9,y[l2�)B�	,0e��4~p���|Y>Q��7���J�Ln&u�1����Q��Ź �0�� u)�� 6�w�g�*q�,kp�FQ��F�T}XJ��w�$�i��,�~��얽�i�z1��wdꁢ���,|��Lyjn3EڷMSд��;ݣ�������/����"<ON�k,ϔ�a�'�<=?m3�xA�]f�گ�{3y�D��'G��+�����.5-80����r��G(-ݝ\�E
e�kNJ� U�,� �ct.�L%0f F�ҕ Ky1/W=[�>�_�6Zk�뛠�B�Ϊ�G&�Ǯ�7A��^(p1�p�����SRh#�0�,P:�����nJv�4N���,8;Ϸ�( �.�tu�=�������wk�Lk ؖ������
��Џ��;�%�lϵ����
LP/-yKܘ^�0iR����N�>$ظ|}ZD�;���@��S-��v2^r��R�q����u�FU��j̋F�"�y��u��pߞ��ß� 4��4�����آ�b\�� |�ч+4ٷw�!�߽1����_*|nq�ۧ܍	h�0�h�vЭ���s|>K��������|�NJ��9��z0���&�0�g_��nl7���0)���gx����F����Q����J /����xz�[_1S���|� ] �� �����������r��MZ�&nRO\�=lh K*��{Ý*+��¥g1���(�L�a��W��ƃ'��n��D�_����|�������>7��/-��M�@�h�����E�����BT�I
�P~�$�� T@X1�ӳ�z����\�q��O�y!�����a��?n1�Bw�]ulgkYf�k�z������ 4��f_�D3\4�" ���_��z������pV��̦�����<�_� P@I8���'�
�6|��S�Z:�_|�u>x�RT���kf����Q����ߓR�;f̊% �iQ���J,*f�G�[�g4d��
^�c���N�4t'�"���a��&UX#��_FP~ �,����}Ta�@K�r]s������pN���������x��_������*�f+������
�S�?��7"��1"\��t� =�d��2�o`b|�6� ���t0dy�� �ۚ��{��Y>B~�h��8Aj��0�@� Q:�`Fq��j����,�ǐ����X�^���l=�FI�6�Ct���̴l�X�~�\��/y�D��_���21��)�H�@�=��N�B�H��ӿx�d�N���b\�W;C�����.�襫��}/#�^������^Y=~�\
�U6��Ǔ�uu*3�����>B��������! ?���(�Tv�r���;��t�C^��~���$�����elG�ǹ��f1C��p���Z�P����� ��$RQ�΀���F2@�� ����)����Z��ͬ���
���(���?0��'Ih|o�/QAZ��nO�{����S���#��!��˿ ��n����7��9湖 �6����U������X�uՂy���v�\����ʍz�؀�s1#�q��e�����(�O�������$e���_������x���П-�9�KD䴴�w�8��7�O\ݙ��ǁ������^�k�8�r��׋����,���n�r1�~,װ8pg��H���zG����kƳ�Bw'Y>t����2�}�2��̅�;��Bp>���d�Q�@u魩���m��A'�����Q�� �:�Xꦿ�Xm<��]��se��Yюo�]�W�
��ǈur�J��M��r����`��" ��"�I�-\O�������&��<���ݬ�u��Z��~l�v'(��F��D:C�@ý�Zx.�;�?��="���ͨ[�O_n�U_feKd
� �UH#�W�}��휓b<nϢ��ΞZ��ܙ�n����+>)�~\�
� QL3[��:<�\�uگ�'.��j�F��WJ`y��UGZ=o�M8��2����*�0���x��Wo���at�����m��`$q?B���D-�W�
3��N�/�n�h2 �P��E�W�)�Aİ��xI�G��8ɋ��o�(��yw�ٮ��S���g	3�����W+��^���l2����!��i�.��t��.Y> E�.4^]]��hv�.��EvRR�Wr���|��z�5�7���	��L$�*L�j"L�Sn���^=�\�������]Z�٠�� p�=�f)���F�K]]^��2I&�����𭭭������)t��9������s�0��e]�7�׋�-�NX?��������|U��Z���!7L�bcc���.-#����E��`~VV`%�b"""�buU���ʕ���q'j�C:����a�6%yy�K<PW�����+J�� ���,AY5+;;0dsk+b``��87gjH�׎ML����:Uo.I^\\LII	S!��ɒ��gg)���:9�B�L��}33m�(EDD�fffbω~�r#'������#111�hCU"C�x�����D� ��c����&0�����p���R\L�1�릧�����@
w"9HQuCC����Cx5�0K�����Xf�{�W���$6�8�Xmm��N�ٹ9K˟�@�X��k���P2�%2�e��,����2Ŕ�����/��^nF%�jNN@P@���ب�q� �8%%���R�K� �Q� Ϊ6����%a��ܬ[�UM'((�*�2�@��_�{&Y���SS��׊M^��  Lxww����F2t!� zYZY=,þ1U�����(�'�� /���J����� d(3�0s�ktQ��ΐ��)7pp.W���ZXX�5t���]�	2�GzYƆ�]���EL��--����>>���<Ȓ�H ��p"	��'$��z����G�Y3�۞��^�ズ2��ʼ0�a�!�+��W��UaE�@$no���<�_u��Od�~���|\^^>67�.��ϐ+s�p~qP�ّ
PH}5fCH�����dH��oP3�U�(Gq�Ww77�dnɽ���aTPWكE��C
���JJ�qdl���/ܒ o�R|�����슊�2N�g~b�����B=�������8W|���wi�x&�ާ^�d�[1���![,���I���^�@�G�AU�-���8+g��o���Ly��/��As�XXXDA �u��Zo��^}2��*R�nۛo29�:ε�����X ���5 �<n.��si� �rs${���?�Rj��I-Y�m�_�@ʍ�� ����:��:�R�<T�]"��e��B�tm���h�.���{�M6^�YW7>*��Z���s�>[�Vq1�|� �q��0,M-ZL^Ӓ�Kn}�����L�qCke��/K�D\Ymn�,y]ؿe����Ȓ�t%���I}�!��¦���覃h��he�Ty�{V�������D ��	(��?�.P��~�#��#����񮮮����e�����\�h뙭�G�T�Π͘�����Ckt٣�@_���شv���F�d�=�1���(
H�YF��/C)�=p˼�#�I�ؠ�oȴ����� ���)�W�  t�~���
r|��$%���n�[M��4�@m,?*R�̐1S�ӏW*��"�FI�x?�����TeJ�N�gh�@x2 �v��y]@�O��7�3k*���	��O���Oo ��MZ�,��ȋG+ژ� ba�
8�����0C3N���xg��|_��!���s�^�f�1;�^x����9I^���y���A����v&}�z)��v�PCt��EԀ�� �O�ʏ��eղ��p ��8n8eڱ!���:.#��t�p�Ls�e�v7\&���~wz�L��	�7j��rG!���5~��B.����g��5M'ekū�;������X��o��ɩ��줱���_���+B��3��}������ҫ2���h_9�-�XZ�2��wtp�_KV��)�5�d�>FtO��?0��#�sƤaS�9@�ݢܒ�#��/ǹ�H���H��]�o�e��U�D�4�zm���' �����bz^���vd��Xn����ҏ˝��Mb������h�{^�����˛,���XriǏA]?��ӧ��MI"�f�*���.�Э��"9((H�El%(�H�$H,�J��BDr	�sPB�d�9�H��5���y3o�7o�o��^��j��瞳������K��j�j�_�Jۋ���
z��)V���Oy=� ��-�vŏ1�?S��5�����ӆ�`͗Wi��U;�2�|�C�^� ��S���v��0*�|.`胩_���5���3d�ε���W�Y`�������I𳰞���.4y Us�Z�A\������CL&�Eu�����Y�	,��{�hs}���V���C zk���>0Rb�F�@�S������A�nb�$׀���)���C�ueh�Y�r�^=7�y�/!0{�#+��jH'�a���̙5�������T�}��\VV������-8M���Kr�{'Yu�R1&�ɑ6>$t���c��{}��-�h���*o���YI�w�%Vs��ce533c�]�'�����b�s���
�$����:��/�0]\�)1%�<��<0��π��~�^L:��Ͷb0菨ޞ���{���!�S	p(�E�������]��7�x�����+#���N��~f>��:^��v��ZW���}����Xa
qA&s�O�${�))�j-	�ZuF(�vp�0���=wW$R�=����gX,.2�j}m��bj�������G��S�%7��S�W�&���Z��Y�k�<��2*�+~s���O��K�4��E�-��|�Os>�/n�6~��w].*G�K ����Cg'EFR捁���^_��y�[ev��w�/O`}�Y2b|�;ޗ/ܱ�����?ܛ��X��dsn%Oy�89�c��K�+�#�B�}��,W�,���UhK� �r�c�>}���8������G��끏����_������k}	�����=iK��¥ nYo���j���O�3>\��������Y:ff`�O��h��!��?+X��ؼa�T�ǧ�Kl�3,��I�ҊMr����Ķf�)'c��9��a�~�0�$�։�ǛUv�;ҋ���5�`��@	�1[�YX��G�	���Y�J�app?��`q��:���(eKf���E�$�������������F�&�k��oj	f�������jjj
�Ȥ 3�]��
<�;BbX��nv�:����<�xD�e�wĶ1��b�#�aa*��a�Z\�a� �}�`Xٰ4�%�7�rW|ko$�#Y�f��"��C�����|�$!� ��m��I�\���������ʷ�5�ZI40؂ݣ5uѨ`�!�������Sߗ�&$��O&�_���Ԭ�tF�}�u��9�$=ֱ0�<=���iSp�긻�ǀ�I�D�֭�c�yWW\�Z�3ۈ����lidE`��<���}'��?~\�1�#lL���	 � Nҭ�;V��Ť�]�*�ݭ�ꃆo�W��.,-�t��f;*�D���{�toR5C��xk{�n�Vr�`���p�"Zht��9��@�s_ӝ7�G"��m��C��o�U}�\�&���~d,&�"c�n�+�j��6��E��H�<�[i5�~o!_u5ef:�<gV�PxH�������T�o^F���g�rrcR��N@����i�� -�Y�,?#yQ��E�Y�Bu\'1y���f���� ���z�9�O�w:�d'����x����s�$���y�f�Q,�FY�5��}�R����ei����u�pb�*�g- �NOO�X��u����,$`�
�vW<��
xypG@�h'��Ġ��ss�/���ze��(����g��`R���?���X,`���v66\�1wڼ�o�,2�i+��D���n�MD��kbl2�Re��[�#W'�n�M�R˱B�a�Ǖ��CSBq�S�����O�L��@�h��a�  �9G�_�F�uU�TW��P�!~�e��N� w�(��/��g�׈��%����?��P2%����&��n��?~\��L����,0�***J �29F=�A&��NǢ�ٖ��)�+��NJ�%GL&�/�i�/��|���v��:Ji�! �Z`u̽���<aK�� �����R�Me��	�J��)=�������ު�20t��S]�*r����E(�#�����O���6~���#dd@����f&F��/��
�� ��+��<�"�W?�4x2f��3αs�h�#����������X�$Uvrی��M�dʙ�T�"�k}Q�ߟ���8 ��!Oݟ,�\~���B�!�R�!jyy�_ݟ�>��AdJ��0M��D6W_�
�OtPe�|Z� 9��&_��JW��-v�7g�0����'+����(���l���t�Ce�Ƨ��57���^<O���s2L�XW12�����)��#%!�^��Td>Ƅf�¯wD
k�B�1�ĝ�Mr"�.ClT�S��j�bj�mƶm�־�}�g^��,J������j2���3`���ν�}�4�
�8�5�֘��l����&�l�e�]�����J�?$�7�������Q��\	�Dl�J°@��9.�nP�m������V+%�X5� }@�pt�Տ���c�kQ�rm=ۣ�5�	�`�(��f��i���n���yj�߸?2��pd�`��B@O)���iJ�ԛ~�_ř��S�T��>��	?���aE���9�TFH{�LW��(�1�]���T���X��i��	k� a���9]��{��gǓ�*��>�߄���f�#�1�|��x��+�Y���=��p<�����`N����lD����~��~��,�=�(x՘k�
e�.�C�O��'�+�>�>��a�W&J.9O'O�/V�����!�C=?:.Z�*�[:�v�z/4����u�*�#
�C���*e8�KP�4.����Vμ� ��鲐�Y�0�7&�sc�ҋ�H����R�ߧ��7�1t��{��P��Jsכ���7�lԗZ-�s��n�r�����)�#`fAr=H�B*,���N��O�G�%Ta���O0+�ih(׌ 	�t�vJ.���ׂ �T
d�>jqY���{��"D���s�Are���H�Y�pg����A+B���u�X��9H�v
$��!��i-I�nÿ	J�v�k��>|�������1����0	� ?�9ّ�������j��P�PJ�_��4�j�$e/�k����φ~�@7OO��� ���rU���!Z�1���x����#��r{����T�����F�Ѥ�����q��A�P��PzJ��$� Ҧԁ��a�(nVUUm��ӑt��i�=�"��Ez�L��`� ���R\v �D6 �JO�?�[���1�9)S�Н�6�=���A������ϢdP��1$�7@�r~'L�X����c?�P��?ˁ@cޝ"���w����u��@0� �d�;)�Eu�K2#up����X���n@�������(����K'(AԀ��`b1�P���ES��6|�d)B�АLN#x`�)9�+C����ѱ�Nw��`;;����$7�l�;̼#8���o�<w�G-8i���M��c	��J���:���z*�i�v� vQ�լ�������
Z����ʓRY�ֶ�� �X?W��W.��
IIafEq �Oxn�t�����:�1�T�9��5H��y;���hCb&�f��e�ף�e��X�n��B���CZ����8J�HR��~�#5�Ĳ�'w�G j~;ZY�@�6U�%8�w���ħC��Ф_�~2�� �q9��T�����W��ȡYh�LC�M�h�9A�z}�[�\�k������
.M"�+UoP����s��"�ed�z�V��#��mVh4D�a����Q�d81��I�I�	��+��C龞��.[)����BQ��.>�˥J=ʘr���B������;d�BLF���YQ�~�;�xQ����8=�Ǥ�o��"Vb��9�&�����Gs������N�5ұ�����N1��P�4`��c,cTbܓdiY��_4~>��eK�+}_�me0bg=�O^Th�@���T0��us��,2W��R�
�k�}�Z�3lhs2��(u�����Ed
Mu��UDy���G����`���yƑ�"
g�<"$�$[�crt�>ӯKKOv�C��"(l撢f	ƞf8Z�|r��r���_z\'{ef�[�h�%���ͺ���q��纉�6]Us-aH-�\�X^^M�+d�VV6�����y�\m�)�4��\ 3���g"�MT`Eb�gE�sy�O>�k`r.��m�U�.hl����&���5��]�v��(&1#q��O�ݲ	�\zF�5��j���pOT�J�}� �Af9��+[)Ѩ�!/���o��vc6k	B��-�7arB��t/b���]��ٯ:�*f�j�$	�`�+6T�<@ǭ��4�*�O(>I� ���ZS�	�(�!c�(9>�ll�.���r���q���G&S@/�UF3�L^�jn�L��.�yd����q�_�bi��rt&<J(�~ƥ���r�=� ���z����K&t7��N�*���b̕�8�3ӿ�!���|�x�a�wSN�N��wC⑊Q�b�_�ȳi/��w#�J�9�e9�X�p'җ[�� �M�Ϡ�������?����<t��㨆�*��=��K��;��?_&�3i�ʏ#��;�B4�o�U�I}6�A���6m}c7B�����&�nq�CAt�0�h(�x厷�ո�DlF��'CWW�P�'�8����\��s֌������!רar�U�/���i��]�^�lB��Խ�=��gs��l�B�x��m��)M�ca0g󂀒��{��^ }��>̂�q�_�G�W�߹b���eh�P��������X}]�)Z6�UԷ�6��&NG�C�?6��|����{��H����f�Z��d�9�S�݄�IMW��w6"����qޘ,�`HJ�l��v�8[f�F���n�Y������r��#�_=���؂~ʜH���"d�[�F�
[U�R��v��O k|�	�H61�r�l�߈�ؘ(��5�21�2��&���Qf��gn�(!-�4�pf��L�Zخ7J����]��F_\��	���ZN�af讽s21_(9+:4)D�wR֩4nI�R�5~��_~���۞��ǈ��B+��ly[���`ina������A��X8���{�^ґ�:��Qޫ����\��&7%^6R�^��<��C Bc걔���~L��e���ӧ�2�e���d�;Z�R����-I��)gzn_����*cK�8����4�������*S0�PѲ���KG�u��ږ5���0��i4^Z��T����[I>�z�<�:��q���x3�U����
���A�� 5F>�������\%�+	���a�Q$1V?���&��I"(�m�2�O��Ig���Hs��"�\�~:o�Z#�bR�=�Y��V���\�]��n?�>��s����Y?��v���GC�n͎�LMЁ�����5֒�-􄡔~�Q���0��T�3�q��	���� 3�=ZC��NMziB0�k"�`���o���wxH\[�?�3�lSSo'�:�B�3�%�'�ih�������)f�G��i�+��]GY<
���CP��P�j��&�?��#���p9���`h�^�T�1Nr��p�\k���=���ˍ34�}13�Y�^�y��/B�LVj�D~ jk#w�mLx�Ñ�a/?�R=En��w��b�/�_�_�x�gAw��黨�woμ���4��Y����vm�7�c��'kvߜ�h��E4�i]P����u�C��y�;�d�����ȣ�Ĕ�T�ά3�'���L��1fƓq��{6����R�f����W��:�+�ʊ�bQONv�L��d����]m��ՒJ6?���^��ix2'߽�e�G�Q�0!��ϴ}G@7� �q��_3[]���>!�����Ѹ$(8el��2&���	k�xƩ;��e���X?c2�-oX�������C/W�P�C��L����]!]����P,��C�.�q�@6jL�@;Ӫ8d���ˍd	3,�4&�&�n�`���}D�h��ds&�#��\�<9^�f�I�>����g�Vz`��5�+7�e'')�<2^��##SCAA��������,��8"zX��Ws����K�?"�wy<\�t�4�b�*2�]O�$e���N�,�p����&3�+M��U3��P�kO�Y��!͆ok���W?�*z1��g�0R��4��{�]qI�"~���d�S$�dd�ڠ�6�xrX.�h��F;yR�F&���q�I�֏%�T��yϣ��)���V�{�X����T]��<"��D�sؐ��U�V29����	�� r��ٲ'/F���Z�f���c<�B�%�\���;����,����\|��I:�|�٢��qs�X3q/�_�����WV�R?�,j�8G�_�2J/ڳ��]#�t��T��z7i������lԈ�-�1�1�t��z��F"���G���/��WZ���ަ)����Gߨn�	��3\nbf��gĶ��5q��w�F�u�Ũ6��[�G2�g��zG"C�5'BA>~�r+ͺ8Հ[�-��g��m�#�������vA+|��%:���A����-��ղ/�z.����'�t���v.�`.�������AiQ�=��?+���"��S�n<��}�=�]�W�Ճ#w�!�!���-f\�z�J!�P�M���E\f�=�ڭ��� �C6Tw��O��BPP�&�#����� B�u����U���2�G�tGk�h��f����j-�4έ����w�ޱ��A�2,U�|��1�<���p;���e������c�'1`���d�a��L ��lnK�[e�6�����\���8��`����Q-0������Zx�#<?� �����
�����utu)f��O.?�j�N�흚�Z��=������Ϟ;g�+�l��>�B��U���g�B�T�Z2�/_�\�؈���Y��&���뇷�����n�P�M|���J`N�M �+�a����_��{��9��OKO���"�i�"A����?�y�\eHq�b˷oA��Y�ԡE6�K�����`�	�`��`ｽ�K���L��nƶ����I ��6��6tuum��MJ�|�	�{����C��G�$���(0�< ��ܺ\c
jj$u>�=ML7�Fw�(��P\���@���bۡ\0̾��o��UTy���O�	+�X����|_���f`�D"I}c ��ᖄ����͛N�������D�MH@�����u4 c2�YB�`�ϡ��i������u��}�a�R/�>\��EZoN6
��҉+�P��M����ZZYQa"׳�޴�&<`"3Շ�=O����m�P�yc-ťK�HXL�H<>�1�K�V' &?�Xl��\(�:W�ŕ�Q^8�Z)��Ko�E�ϓz�(�*�h���I����s͏ĉ{��}3���*�4ESfpA���ϙK=f�5���e� j���V��czs[���P�cBB�A~4��F���d��:Y�i�gMy� �ns�O�;K��?��(��� � ?�uG������n�@.D���i��^KE"+F�x�|||d����g�G�#}z���gi%�έg�	 VE��A�eV��)�9Sn 	��駼.4�ԅ ��_����҉���~jy`}T/��m%�C����{���O*!��%%%r�kJKK	E��ڳǶ+��}�Ã<3(w�a���C��ED<x�}7f�:�Z^�z����!���{���y�%Np��M�2�y@����{�#q����m�$+!$��tR��n��Pw��a�*>��Z2E����d��E�E��n6d��$��T�IP�O3����'��;&���0��)���m��^��P���!�i]!�n���p
�s*CL/x���W�m���X�7�U�u�sM����\#��Mf`�ԫx��m�/ڀ۞�>?\����~�y�b�N��2:~Xh]��,�!���L(����#�z���4�l9F�,�jʅBP^XX1I���&�9���i>��x4K���H��`P��|�׫�X�b�U5���ڠ>��z���e 'j �gw4�B�@@'h��{�|gK����Ӕ�GX\.~��L��H+j-��!K�9d�F��Py �{,��R��J9��~�:(��$��ǌ�~�(��m,���)٨7�U-�8_�ʮ�v4@���,G+�*�l���7ÀS�LC�����%i���r1����O�f�5`i�YH�i�'�J���O���i�h�� ��=���Bk��<�ÏA����;���`)��p9n��t���Qp�@�ka�o�!c/�q�j�Y���k�#͹'�n6e���Ҟ��C���Ò�.I�L��ȣ�������Cqqy��W�������<�!�=����#�-)3I1�`�u�s;���WֿC��]���Q��6���G����F����)+��M�N�MNS�1�������<-.0��-�H��%w�2�%8(��K�	�z�o��/�M�#�%�����v�=�GC�^ߑ�L���(�@�M��!PcJ���m�L����RC	P��/^�,p��|.L���MF�[PH�*�w�oͫ��� ,򅈡i�0}x\J�#&rA�h�2�\JBJ
J1��o��N�)}�cU�3�hkk�0��HUU���h�߲��>@�6�-A�ke��@F���VFS�_H'_���9��"6��q�=�G�(E��e�|�KLhrX㾷���%E�"����8�v�LA������Y�J�g��B��ן�*�V ���T4+�y2��ZZ]
B"�?<�yg��23���l�4A��7Ԃ���y:�!ޓ�.?7�Q&�#�ϫ��]]�Zn����H�#�R��'y}�)¯�ͦ:�d�q�Dɇ��8�6��)�9W�;M�qE+�����3�`*r`�u3L�wE{�WQ�����]� ���>�$������Q�A8!)�,lz����B���M������eU�}����W���*��#ƅC�Jd0��)�� o	HU�@Pt=������0ƅ��{�q��� l���V+SC��I�����)Ѥ�������ͦ�/����3��/8����&��W�߈�^O��Ww�UD�~u���(&Ij��s�J�.!11��H ����t�W�C&�K���j*N`��a�ɬ����}����t�@w�j��-�4�D����8��S@�F�{�)�Ҿ̔��z> ��(�+����>U�(_'��j����j=�1�����V���� �|1��z�����x�+m�|�6Ǎ��w�V��Q��\e�X�UV���*C��.�<ܠʔ�ͽ{�z��#.���O�
�J1�ٌ�E��L��f�@�G5)w'�o*?*A����Ŧ���=%���[�XL����0ח	d3*��lMx�~�����
HJ2���@E2rr�ޑ�x�{�/� �&�*�P�Z��:;:;[��܅�?� ��;�Ѐ&������ }�Z{�A%#kM�����\��ޓ�O/ 牋���/rQ��yI]`?���R�/y�mJ.-�P��T�#���15@@Oip(�6e9:yP��z��5�I8S`��͝岤^����������O�k���45���<NJ��=()���z؄�:tWz�����(�[2(*�����)��O�M��5`�1�좱ղ!c�������
	w3�L�)o��F1;��il��	��}z���
1�ne���C�f�z��mT>���{�w@]��m�H�W-�EV�>s�}�Oǈ)�E���\���/�M�;��)�����c�}"c��#Ѷ�n�#��J��K3����:��&i�&ݱ.��WR�k�}�x}ȁ����sZX)'_1?�U+	��/s_ɫ��;6�P2[\�ߡ=���qq�{}�V1~�y�6�;w�=MX�j�	v�M �9[�	f~#��#��,�Q�d�$�\|j��h���<�*@�
��_�4��'�TQ�r�(�bՉ�":���+��>k�l�Y�(KgFk���hZp?�"(�Z��S����� o]�Sf��9��(:��j�;�وw�6M5;ӳ����#�+���w&�EL�ycq��s�y�A������ā]��d0�G����K�5���I���H�[E^�L�Ϳۗ`�=�ⵀ�29�CWMXV�` C}#[#�;OQ�E�◡�8=�w���k�D���%��]�H�ys�٦ԉ�f-����|#S�m��W�b��=�v�=��R)4yHsY���{
��~�pwh���d������PW��I��v�Q��K�48�3��+�-)heik��{��dt�i$@����d�`uX���f}�Z�&SJ��=|��ew�ea�°-����z�֬���Y��*�T�|0��3n�lZ X�^+�"V��j^YP�0��;S��n�_�ο���񒁮J�0��T���%h1�,���}�$}
:A)�+��k��";T� a}�~>��ݒY���S��S��5޵�-o��� �j�b8����|�\x�F�� u��.v��W��H�v�nk� P�.����j��3��-{]'�c4���C���Q�O=a^��&�C��q��AG�H��SlҠ��~�=�������,�_/u�]��F�_�iʙ�;#~�
�����е��"�j.�ўT(�,w�/:05A�8��<���:jo�߈��w\n���ér�j�t��!�+���H=W0j9M�מ5��)b)�3�y��;B/V�J��\<�vV�\������՗�G3�WH�=4*�K����
��
��Hn�����5��T��&��h��-�^���|zS�����1���d��ܙ�.RN��e�J��BY��;��Z�Q�T���T�;����t�l2|.�(HT�׶���P�96������6�:n�>�8�V���D�e�-��G�2>`
;�6Ѵ<��~@(Ӡ#ƶW�0������NjڂmY ��0Z�D�N��I�����z��U �nN픜k-����L����mڤu3͆T�x��G�aDK��tq��rW��h��JQ�m6 꿤���Q�y��haн;���P|�2��b����`7�!Hz�ؔ�ino�0�����ns�2�y��^ ;nt)���]=(sjj�(�02	ۦac5�)��`N潜�� �8FHxֹ�U0��t�܁��/������������JX1ߣ��ky����+��Vw&��G�&�k�,�v9X���=nӇ+\��Y�Z�����M_R����ׄ4�����t-��W���2�mH�o�D�m�߂t��v��,'r��t�"�ٌ9�h�Fh��A�쫝c�<�ED����'2�?�1/��X�8ffD�ɫ4w����G5 �Z��,bp��oK8\�a}��p����oE���8a���Ȕ^s�1&���u67�2�#�|-d��; k��R�q�vo��� �iס�f��%<�\�J�o[R���U:Fc�ʣ�^�J.�xf���5/3k�$�/�p��,~�$�b�kyhp�^���ʽ�C
��cj�����#�qڀ&[�K�N���J�D�3?Vm���N�D8�i�����O0���~�Ε6{�F0��Bo����~u�?S��
�ߓ�VJx�jP��]Zc���Ӥ��G��0^�����O@u�uL�]Z���2��_}z���]���x����[@oe�T�<n�]��&~Y1��|��J�fǵ�]���ۭ��A��:?q���4�z���L�k?�Wc���=>�43'Z _e#]��`fg�R��Q��ȁ0��Cq6b������` w���>�,��������?(�ـ� ��e�z�s$�b��Y��R/�I��]>Q���{�����lI��w�J��^Tm��<�﫶_4�Z}�̜�A�]^S/L=��o�8�(�����&\wƛ�64S�D3��;�Tn1l���=w�&R�^8�?]}��Ry��zeGK��fEb��2����p��e���(|̉���e����[�s��Y�{���k�2�%[#���"3���w`�iW(/�0Y)N<��m+Ə����>\�MW0�Z�V�d�:���o{O^�3܀|��a����Z���_�2�����I�P�~�p%4}���5>�fUF��B֝��y(R\��Ӌ�L��0��>ڶ+T��������]��9VB�%d`J��b��D�n�Z��;4���vY��C��U�
��k�؉BI��2E��+3{kj2W�k�o�L���1���ե�5�rx�V��2�����Ch�d:���������N�Z)�	iƬ�n�@��q�9��@�"���b����*J���|ΙW���Q_�"�!	�s3qh�%�r����C�T?�*����r�g���%#K;C�I�K�ۯ^�q�F�]�����Z,[�k+�\��Q2!�wu���|�J�d�A�w�h�����˂��$��J�<�bjਲ਼fsʥZf��T���0"ܳ�z���j���嵐�JE����Of5
ƶϛO��jb�;>I�hJf��5]0�j�5�5~jT���92\1q�|�Ҫ�	C������J.Q�j�V̥V���B�(Q#uT4{����J����xv�K���c>�ʹk��1�.f�����K���|�ٴ0�c��'��S^ׄ��^g50i-I%�
N�U�@>[��]���{ߣ�T����"�=���\��j��xRv�E�i=��9��ԍ �B>s����:��0����*|�p2޹�&W$O�ȩM9~�])V�~�dK1��̐��|^�h�Ƌ��+3��Jn�L��'�qn1������I]�P�u��&��\�� ����I¼z��Z��\Q z��!y-��(�#"�c�������׏�`�G�RĤa�2�S��0EMJ�3�st�!⠪��
i��2���`�CJ�<�b�.�[���r�v�zO+W���r�`�jo���`�M=�o<=�s�_81�����r;�JcJ�b���1�����0ߜA�B}��nr�&��_at���U>}�Я��U��(�z�"�������T1��N�r[[�Q��_W�R�J�j���N�_:8��S�~�S��x�}{f��[܂��pl$.19(j�F9�Y�_���s���?���D1�_�r��t)����p��wl�q�P�s%P�;��j<�R	���U�W����X�3R��{��i�oټp\�����D;�����!&<ី�=���uN=�����1	���$���;OP�(2�@P|���n#iɯώ�j ���7/��mB:LX� �z�5;��i��J�	�B��X�# �NՈ�z�:������5/�T��Uc;����:��;`]I\�W���;�4Љhdt�E��L�������f�s���O���3����Ӕ.���7�q�����i*�Z�Bw���#`�5�!6e�I�+��u�Z6WڕGv�R�D���,-����x��6U#�s����TEL�G\$`L7�u�k�1šڪl�=w)��k+*���� �q@�y���	HKSc9v�2z�q�$9�S��pc]�U��L�a��f�wԋ
�4�}�wr�'�Z؀�:\�������e��S�{��ˬ������_Wii�S�}����*,b�o���B�g%��*�bj����[�hx��I!���0���ƒ�Jj���x�3!�n	�(I����� <�d�RQ�䅳%�f��^4��i�%�O{���rA��N;7��}��$��/o������3�����a���+�P1�LP���S�`Q\蚔#���,�T�i4���Wk��W/��:���D�����٧,r{�埻qA�>&]�w|1����(��	ѱ����C�i>P ������w�Og����8���[�>R��Y�M��x���	yX�jd��������L)!]�_�Q\�)�� �f��'X���1�p���sRϿg�C����J�]geޔ���g�JY��t���|��,�fFC)��!U 
���4�2��k��Cݻ���kA�mآ�w���K������z�$�|q���Z���9��r��[s����si���l0�ɩI8�f�W��﷩�Xcm�߰In�W
��k��\���xڅZ8�����Z�Mp�[�l�x�<��p���tf|�,�ҥ��xtQV����"��c��������^~��`R�@�`av��і~�2��8�2Y�-%�2�>섏;⨥�{1e��2u�e		ݶJX>��s/�X�l�@���P}w��9I��zD�V�$�����H�����b��P[U�P�������8��L�#ܺ+�߽��]�:�:�eQ�`��2AP���f�Fb�a%�iGe�9�U���e�U|Oy!�b�[���R��&s`���y��%u0c�V�R�ͯ����[/c&*��-��^��\�D��AKyS�K��8"(Z�`!�+���/0$�H<	GM���1��璂A tZ���\4�9�װ\�,�q%$�`�&���N:dh��BH��h���ƒ�j8h�3�~O�`23��ߐ�V'˷.�����Tќqy����+��e���z���*���n���X�~�G����E#��n�i�w��z�������D͈��8����b+ѐ@;Ύ�U��1.�0o���BVʨ�B��oD9ҿ�ް6<��NUK��<\l��^����.�"�h��6�y����a�>�H7_'��یg��T�VsQ8n2gãk���"�f}dd'�[����.fŌ~��J��
ɒbi�Y���k4�gn��%�H{^�(���Qߞ�-�c氩��.���+X%�R��/�?����D��͕,g˙8f��\j�-gFi�M�0	exOGE4�x�@���Z�}8�[k*,��y����Պd�S�To9z�֜�%Kӆ�l��a��\l-<b�T���3$PO�ǵ2O�K�цm�x.@S�.���[yy]+�A���|sz�;12�H|��l��T���F��4��`"�7��~�nX̩�px=֫o�}�(:*Mc땭��n~u�l5��>Sg}��]���ޜ��.<*_vX;��1�؄eg��dFU0Pyy�^���\~ve#�R;B�U/�H�^��!�w��"!\+7�W>���
_�n��-�y���"uEϵՀ��NRPK��j�HfRk`7w.���������w^�exӪ��v�v��㛵��t���`Zz	
yW�<s�'��p����-4��gV��n [1tK���%9>����ş���ĢJ�����r�"����`�����S>^"�ɉ�����']'F�'�R���F��GX�橉Z~7�G���I�$X���I��/�ݶY%�R�O���%B�x3eo<�:zPS	HÚ��j�}�ߥ�"�P7T9����)e��U���1&��y�Y��
Ԭx��+��~�e�E*�.���W�>���_���<ٴ�P�_G�j�Jj���hbu4�fre�`�!��Rf�ݝg�xj=�3�~g��WI�:�K��M��팇b�ʖ\�G8K���Ѻ�� ��U�Я7J5 k����G�P���@,P�nL��o#hH�t���+�0����GQ�~{b�E�g����c�sM'��K��6�e,���wDx�l6\��3�{�тos�^��mQ��%�>S��m�ճ��"75fM!��[��3�$S��t��kN{�[�� ��2��q�J7J֫;���N=B-;x�ɿ����)ǰ�U�f��L�X���E�Bb��Y_�ZW�iNȾC#�|�����|{z��I���|�>�~�ΠǶ����~�
�lw��M�r�d�X_'��cڽ���}h�(Hװ\�d����XA���ˊ-�9\�d!&g��5XװH�Rz鬗����z�,�Z�d�.|s�v�G�(��(�s�M��n��P4���y��kf�?�G$�Q�0�(�`Sd=>1���Ô8Ԋ��4�˷ǵߘI�����6���""l���x��F�A��<-��w������w��z=֣�d�0�����U�(L=�ϔ`�<������Rނ��1���z}bLܞ�X������Y����֙�Iq����99�EJ�[,~S�+��YO��"Z
��������*����������
�O���(��[V�zN���L�V�XDi��;����roD,��xh+��W�p�HD��
�zB(�.S�%��ȫ�y����t�;ZCRF*-��4MR\[�4mdQﰛ�6c�J+�����u���M���P�quiڇ�<��.�A�u�AzG����!^=Q�C^�q��<&�у!a����6ǥ��Ջ�T��INH�'XJ�9��{�������ϸ�s#���澏ojw���ǁ#]ւO�&��]��e'\䟘��Il\)�mC6��o��WP^^��5*ĩ��vG⻠������Lf�ӱ:KhQ.��Rg(N��)th�S��h���3���C���v�1�~��ޱ�J�"��P>����}���
������:~��-�5��B���IT�@:�.<z$��6����yO~�{Ց�5����i��.E��=v��b�>���rR�!Ci)��dZ�(��#���hv7;d-q7;I�8�<�Ԩ��RDɖ2����%�+�~q9~��)�nx��}�+O�i��޿b8���'/?w���j��{޸w��P��F�$�E�ޑ2�~M\��5_ִF�}(1(��[�ͼ�}��˼�/�,�e��3�̾����������9�Ѯ�v���:�+��������_O�������A�^QM��T���HW��G���c�<��M���:��є��|I[���D�n�{��?�߉#N�^�Sn�۟�َ�<�W,������N(#15?:e�Y-)B_�c��8��z@��W�h��[?��<V����IΚ�#���I蕢y�m�z2v��J+�$�E��J�6J��^�x[N��&l����62��.Z�p�,�p�r��0p�UZʜ/X���e�!��{���r.��^>�����o���N�[gUժ����޻Y�� n�:����.�ݙ��K%�÷>u�B?���n^�T}�rϳa�A[PP��i�������NN��݄��U�Ԗ�R��H
���е�����o}6o�2ߓ/(4Ѹ>����R��G�Ś��ߪ��g?i/fQ|^�:MI�}��֗���Nv˴��^�&���$)#�=}#I)��j�8Q�e�W�����>����}��'���K'z�>t1�2[T5�x\R�Z��s���j7xK��;��d�205?�����6W����d1~/n��4!�q3�2������~�ٚ�8Q|V�cޱ���<�jO��[�l�(�]���+xՀ,r���Z�X�O#ꯆ,	�^�/^7��%�&�ck�!���>�C�@^5&��kzf�*v�[�:��oFEӏ�/]]z�9�|�/���$���kje^=�f|�E}�o�A�i'i�F�Q8�Hn�wz���R^�[p.��н��IAUQW��^Z�����������|Z����oޤ�v�ʩ��֍N�<����%S]Oo,Z�z�|z��k���T������l���*Z�FQ�>t#�NA�%�ҭ �҇.��F@��CZ�����ý���c ���j����-٠ù�
V��O#���V!l��W��8\�p�ϔ5��Wʕm;�����@4M�ӠlR��H������D<�xV����0�2ױ�"�T�����Y�W)���m�ӥ��,r�sj!�5�.�.��­`��ܓ�ukR�g���x��n�������1jvP�ZI��6�|�<!�	��#̗Ɩ��RᓞZ|�\�"�Ĉ��8�84��ͭ��t�[�䉿�������ybS��땗'
����{�K�m)�vE���B�=�� �4���+>��K�@��H� ������]����&�xض�*Ƹ?��`\�25�����=�F;�����7C�����a1 ������dz�S�FT.�O�_����"�;Z�#ҳmPI:����\)�)���kc�d,�BD�a�@" 0���YZ����kVk�Gv;����]���u|f�>�~_��v���'=�@�C`FD�4�+,4�!bc�I\�ڹm�B�S��Fp{sS��hq��18��&
;����MG��GG�Iۗ9��Ri�hg���˶�8�'�Е��8(��:�9�X�>���������*���@�
����r5�<�-�in&�ӊC�=�sb`�:�x�qh�W�E�_�@I�������]���pǞdYEK�<{��QSpiKȆh�f��ly�`�1��E��͗ݨ�E���x��7�'�2�7D<��)�_�6L%�3P�2/ش-Qx���9(���*���;�U6He�=�}|����o�������pz����6qp����I���!����PF��/808��4��#�G��#H6y��D�(�0��]o�>���
�����7���^sک��������f�ca�)����4(���+3�|�CMƻUޤ��5pzZc��b���D�)��(Z�T�D*�F9T˚ȧ�;Z�T�7��ZR7m)B`!J���0z=�i� qg��j��AM�o��� ����/�]T r���u��� �LӺ��S����)�_�*P�G(�=c�a�I�u޿h,��h.#WF��z<n����ٌ!՝H%�Û�Ou5f�����D�����2�x� � �h&�g��� h���,�8�����,��1�T�Ȣ����@�雚�Y�U s��Ĥ��V7��Di�W^ո� ���yb2m�V�LSw�\�P�fS4� *����o����?�B��?����*`j.�����ю �����'��0�>��L=
�쀀��"�A�2$`=W�*J�v�-����[3�o��.�'(/�vb��������7\l�-�i�c����o0���V�c�}�����"���/Z]��<4:Q�#n����]^U�Z���z_:1Z��{�6D� bne5��=�j�:�5>]��ó)޴V!��&�c+�~�X�@��ie�$�+$w�(!y�9Y��$�����o���<P%c����<�a������!5��z	�S`dͦQcr��j=��l�g��K����_�c����X���i����z���˥WE�u�;|������O���g�s������lA�\����=<S._�a�b���b���o�`)(�H)��	�^����άR���rT	F�ʑ{��?I���E�
z�S-��
�����gXC�������90���A�I9�~��t#����̵�)�_��&,����e �J�8Á}T޻�
J|���y��,U�JO{����ǂ{k�c�#Jʘww�0h��5i0�%�(�Q��n-9���"EPf<
�?��q��vH=�'�ˋ�Tv��s��+���POf�ϻ��L5�Q>	�MJ�Aͨ~@��X-NdNt�Fg_졒��撌Rx���n�lS͢���_�7����@~y ��Rs;#�~�'g��7g�j�8�xE0�!���� R�^N�����E���/`�2;�[���� �d��4(K����b}�����	�m
�ϣ�}[�*|���q>R^��eSÍ�[��>EE��t��] +y̬*B���]Q�f^��q�)�Og􋨟#*g��:��߉m���r������f�j�2����)�6�[/�l���`�^������r��Fe�ӷ���`�A����x)gIlh		#D���o��@��_���m9N �gR?�G'퐻��g�2r�VOdҫ�veOw�EQ�q�e␍���W�� x���ʏ���	�v][�3�kI�EN������Rǭqrھ���}lPܾ�K(��r�R������;~e��4|*�˾Zk�E�������/�s��r�|z�ޑ�EĤ+�(}w4EYu|+�0���d�ک
ƃ�gÞ����@�ܲ��3��E'-�����������g@"Xbx>�ˆA���H@�9�����U�9�i��n�ً2l�0����$e�Y�NJ��f�W�HH��j=@�AkC,�+F{	ˎ*�f�j�T�OJ2m�p�A�*��4 b�(��IV눼�E��9�YQٖ��g�Q�����ަ�K?S�U�K#�$�٪��I�,��;�@�_D1�k��I�:
 �#%�Q�"�@M����˓���9n�d&����0<�9ߩp��%,r$wl�g�����<�W�1��L��=��Hj����n��p�Uק�����N���Y��߿��l���@I���to$��� ���=F�9���P��.�̂��{�>ԮF�}�jnF��Ƭ' ��)��7|��/(�`g�,�^��ל��I	ںpں��wN�@ů�� 6�ހE���6N���w}�?���38Z�Rm�s�����CIty㥯�a�)�c^܎����B��h$e"�x�,���� �G��l���a�};��X1�-��O���D�Z�a+o]#�U:ٗWv�k&,�|�r�-1�݆��Co<�L�FB�'+�+^W�xހ<���W�*�o���Ϙ>$`�U��9������{E9%Ԯ�Z���ƿ?��=�0߻e��������焾�sF�^P��9�>��(3S{��G>��`��$��̵�3Jx���� �1;,�@ڛ֯]��C�;�!�^2V�w=e�#h����"PP��J����V��ޙ��щ�3"�m��?[�ι���H	C��EzuO���`I&b���̹�z�� ���[�L�o��y&��t.����w!&O)ٱ$C*b�G�qK+ri99լ�ix��Z;�\�u��x�V��-Q�K�U���àz���Lо܍���2���1˩~�G�1cyR�����'��K2��ò�O�'�h9s-^f��q��E4V��+��OWG��a�&|���V���W����)L��/��W	�3��ۗ�R�4�L'�ۡ���0�$l���|���ȅ�8��Ӛ|��kV��F%<�'	ٰGz�r��Ň�9DkJ�Y8���cȡ�T���.��r%�7�!xH*�����@ZH27��}��� ��*X>��51��D�d0p��A�@�4{�h|4�2����3nZ���̪D*��eK���F �ӽ�Z���^7՗/}�1�e��,'1�����!Mr�K�{�?�z����Hؤ;�q}Վzoe�_�4�U�m�(j��Oy5�J廋>:��ժ�e��w}�n��l�?�P��+��o��n��#G�;�þs�����B��
F�L���L8�^@���Eᙼޏ� �&�;�����ܜ�r�0M_g��Ý��>%���e�@����i�|P[,�|j�r�� ���d#��`��{�IG衟Q�/Lt�G8���֧��7�Ĭ:�C'4`����-*�. �x��
�#�"4�6ԩgõ�MaGwf4H��Q����vFtj�[g�M���a���ʧ�Id��KK�_�]�a�E��c�Χ�S,��IH�{����d�,Ը%��0��~�*���a��� ��xp?��}�>��~�h뾉�H
��E����|�`%ת�E��������f�ul�fg.@(�L>��P1	��]�D(�[������_J?#���(��'������s��ݍ�K�>{���.*������i����Jyڌk�\�yD}�����,p����P�p� 9�${r�"��S �.̭�2��P`�C�����|�*�$M�f�("B\�R�Y����T/;�LF�@j�^�$׮}�ROQ���(��`��~�ȳ�x�{������A�G%9�Ҳ
��(:�b�x��[�i�����}��Z��S���1���v"�WF�"���_�Zc{�u���3ny���%� ��%�����6+�K{.K�����*�&Z3��u5:;�+wP�w��-�Bw����s6��w�F���>��'/ς#>/�����<NL`���A0�`,Y��}Ɍ.�{���ĉ�h�uZ(	/��:>f������giD{q\�S�����ş�*�^@�86���s�$3��KS���� /w���a�(G�V�*;�N���ПK<�@�eg\� Hy��Ω�Z���'�#Ҿ�	�xzl���x�q %����(�_ǭ���C9���<&&Ufӡ��I��ՕE�괪�B!���>�QZ��c6g		��yV�I���i�RBշ_�:/q� z� 9%T���9���[�����?���=;���֔��
 R��*L28�ժ��Jk� J�åYb��g\�{8�*�k�y���]�?��_�qA��+��y��k-h�&����E���6��Wۢ����c�'���U��Y�
1�)�=��6�����pV���]�����e�8ٲA#�WA�}6�S}2<O�+�����^�l\�ڲ����kaFl��ˢϭ]�%[�~�X0�O���@���j�"�q�t��Q���Pv��!�i��\�^�d{W����D��l����!�ڮ��q6�|��k����f�?�� �z�0䫨�����U��O�
����i��
�C��LХ��d������M~����W����Yi����M��e�`��
K`��x�������,-z���ڙ�J;
j�tS�B޽ɵ�}z��L�@Fk��M��r�\N7�k����ϻ#���y#B��!U���2��]��׫
���Ɣ7�6�a�}b@�[�^b�]c�`�>��տ
��{w�G�k���l�M��F�a�\5w��ݿ6���5x���ɚ_�=��H�,���%!��ў�瀩S�7$
=���75*|�"5���z�,6��o�JcR�ږ[�����Y7I�����t�{&���I$y��KNH�溡z~G2�R"��ǥs�������;�o�;��xʅ�����щQ�:S9�l�o�k�0v@6��]���^Ca���t���Ц8-��__�ơ��Q�,`�ǡ!^���S+����N�'Э�4��1{V�FLa���IK����B�|�uUI�H��6���oi|��׎r���%�
c4�����s Sn^vR'ӿ&�8~��K@�Hۍj"�O��\����e���#�&N�����������e}<����m�~}�J�Z�K%������7� `#�'d��A�H���!͒��� /�2 О.Z��zF���[ҵNMA�>^q��}E���kTD�yeU��G%�?;Z>&�ȏHqX����>Bo�2o��K0�K]�@�l7�W���[�l{������tv��/�m.ݱ}y�=�u���҆�P�9�����PNſm�㟓ę.	�<֛Ԡ՘Z�N9����\��T&۞T����;�>�0H[T`�I��p���}��˜�=:D#D8+�K� �G���L�^�7I�!��r�ZD����1%���%�^��gK����A�$���<l��4C2�P�7G�\<����	)�_1���%�~8�
�{�t|C�&�7�d�ߗO�� �O�/o&���h�U�M�/��hY:}���N�L��H�"����K�[!�C�t�����pMW2��݇@��H2(km.��8������.���qˍ<� ��]1�t`�}�����:O��n��
*�e�zR:th�_nij������l$���m������x�7C���h��^���M�l)���U��Dp��exѐ[)�^I��t$&Z��������py��ǒ�o�=��k)�Ђ��i�J��)E��z�!�Ԡ������zAO�Ib�
%�9ڑ���� �r3�U��2�nY��SD�2��^S���C�A�%����K��K�p�Q�O��о��^l�3�).ҍ$A�ٜF�RJ�ȵO������hCC�fl���?h�hl��V�<��뎃�4}{*�D۱�f�</�	>��YO��kU���X�7�/����{{��䭤Tԫ���P�P�;6�	�W11�����������tMW����k��2_�<z�2�ys�J�qŞ��C %�Ī336Y��G�2[X����u����;�@?2��
�i��#�h��o�E۫�D.�۾؊}Ie�vT%ocG@�����	�gU���~p��x��'��`c8i�lr�u?���j랏��_O�����I=�0T�a1���}����6�
E�~t�r��J��#�%�:j��%����]V�˳��T[i;<���t���)̑�a^��KuJ��i�C��^��I�=�f+g���{�7�n�-��S������J�����E>+��;d��q�$c�����U�W�@��7,�Q2�uin�����Hj2������qjA�+�ȋ����8F�h����#$]<�@آ9�7�-.
�vߕ=U/�!�f5)�w��e��+E�bD JR~�:��`���2�$a��Oླྀx�>�~M1}߰�!���aЊu�O� lj:�>��0,�J&G��/��N���av(?�A���㌇	PA�a�Wx�if�,����ٲ-Q �/���N�f�4M���}t�Ox$ا/j��YǱ�̊\���]I.^�W�]�)�*y����VC����%@��,��U��I{H��C�[��>���v�ɼ��{��ɓrK�y�<Ln� �F4{XW]K�L^�l��|�Ťؗ�-㨅���*�+����{k*O��K�@�]UM���5t�u�t�P�no0��v��	Bx={�����l)�8|$V����ݧ��1G4�����!r������}��F���獾��N�piL��`P�I�:�v�dQo��&��Q	�Y7�Y��߱5���?�)�����n�C��ݚ�\�(k����y���òJpPA�F��6X���4��i���Մm*�c`�|��--���I��C�m<(Y���!�ɠ����|����}x�K�b51��^y��ozz��Y�R�>� �n�Z�B�1��vlAY4h��a�}����[p��*�#k�*��L���K��j���l�w��/0~`Z����0��@���0�V�r�P�� 
��Wo0:�K)�y��[�}ߠ�ǔ����E����"�;?�,tA[�^aa}K�[iu��T8/����t��b�T���8Rsi%v&p�ˤ�z@7D��B9���6.E�2Qxad�%�V�F Ғk�
dJ{vw2���%��̤�������j~�R>�IwL��ӝx*�U�;i�$x��8�[��d���ޗ&������\��^�ڝ���`����ӅO{&h��O�z��OPy5�J���3�T��Ռ�tʆ�R�(�ua�!oS���U��G�(�5LgT�5}TR|�a�%F�WUu���X`=���C��=*���D$������&�n{RnhJ�| �qig/e+`-E��x\%ј�]������z�t��)I\gUuSضyT)9덗�0����)y��q�2����Q�����1�������hsoW�3N��O�Z�M��F��.�֠%�<���C��w}ѠX?T�w*�����ɤ7�!���-���|����5l(����?y�����'Y���ǦP%�#��oY�m�����~��LJ(��S�RF��A2h%�u�"�S�7�t	~�oh����	�L��d�24����ywL9��
۩%��'���[]�Gû��71����f��qI�s��n�E1��b�ñ)9`Gw����o�W�y��d�_%�~p�yix��:�_�%Q�2s�d�t K������lZ����+��%��oz��(`�?8� @�`vﳆZ�F�U��6�.���lx��C"db�$)S�,
Ѓ��~C��Ɠ�z:�4g2��Z�u� �v7�Li��g'8�-;�P��U�]�mY�P�\�|j��i��3�5H-ͱ�{��86]t�cT��z�p��D��W�^����L^������v�K{�G�Ƥ��֩<N���P��ą��V��(o�^��Nb��mJ�{Ύ�dJ�`9��	�͌�e�ͺ�o�u��������H2Ŧ[߸���K�_Gd�ȼ����;3VVp�=�( ���T��J�ܥ�=Q<$�`���NM%���A2߀�k�P���
X�0pz2ASi��#pr�%7��aw�KН��fg9���|t 2<T� �(0���M)y.�U��%J)<�O�b��U�O�7b	Ä�~��ڷ6t��@F������SE�G�e�����W���M��/�� `5��)��!0UH
�z��m~2��m3�nC�rǒ7���n�*�rG�R�{�P�xm��Y��r35�@5�Dx��e,���3E��3���y�厔~�H�tҀ�A!nz��'�^����h�zc{M��w�{��_�f�m6��[3��w��B ���
H�o�%5l� Ѯ�+2����PA�wWХp�Rb?LDrv1�H�$`NF	|��J�g������ؿ⩘�B�8w��c�5�m2~��s�5��I���&4/�>$d��p�u8��u4���u��i�L�~�B���V�˧\.[��E�R�@����3�W�����V�����1*#��j�ާck�D�0���I�7��1�%�-��GD��j�|}���}m[Ƿxq�Λ��H�8v��\U�w>֡MF��� z{�Zt=�Ei�p��GZE�:�< r���7=&���[���a�߲m�I����ǋ�	(�֛�MWi^QU�u�Q������ۋ@*����
�� �����ˆk��S�u�K��Ƀ����g Toy #�I�<[��d���KM�\��"a��6��7�U&���&�g����S��4����M��Sc������
�g����f+�$�~���c�	�\r�2׼JJ�~�]Ws�=���ɰUp1��[�ܓ��z��jU�������;�[�.���&�I��2^3�J~𐤩�AF�ixn��{�^j�2��dYG�R�8�hߌ1ry�=8�$��	t�6��J죠HN4��ݞ�ho8P�v���q��HܓJŘ�$�!��;QQ���.9��]�NZ����ݞ>�r�x����2�h���
2�ƭ*9цt�rдp5���T�����K�������L�X��p~|��٨4	;΢��.���=�V��
l��?KQ�m�O�o7ea۾�G�o�hq��lԦ�G0���o	��~�R�ל�>���V����J��m���Y��������C^�� W������ 	y �я�d�b(����^DZt�+��S/�ߑie'Rp�[&`�stOϏ��#�Y�X�kXX�*Ok�7�C��k<�*O�<j�����_l͓J�+9�kF�"�׋^6q���:x�C��֕k�ۅ=;p�Ͼχ�
k�k��m�w�Qp?E��z]:��u���24v��M� �;a�'Ռ'_�����c$�Vf���P�~��Q���[���2O/
�Djgtpm% �l�(o��BDb�'3@���ޯ(=p����ĜY� �(���q��5�M�ᡉ��k{�w�z�e��СZ�i�����	8(V
�()�h��]��fq 7����2��lM#؝�)2���)��𴚂9���~�`�E4S�����ߥ��9\�����v�iߘ�ҿ�a\E�f��|i&�_��j�j���.���A�Z��]j������W��������F���#����pq�Z��y�����"�	��mvo��{���}	#6�mL���;��f*?�j����P.D��x�z�L����6(Fl.v�����%4������-bob��j���Gf:7M��Í]Oz����'�4����c,!�_�@]|Uu�P����ǉy�vP�����H��B}cȁ�pC���~
��"{��r���Y���}��� �=�=뮸s��&��`�����8��gyJ�;n�����'��[����4�ieB�L���A4�^���{0�[ЈЌ��Q�&+`����B��i}�8�JҿȮ2�C�F�Jd�ɏ1 OU�Ϙk1N<�d�Ϊ�E���ye�i��aU)��8��0�j���jTM1�������m�w�dU|�N����x�u��r$2�W1:���NA��X��&��c3��J�fi�Z�JJ�Z4�;j�3�����\����iw��y�Y�+c��� �ؙ�S�H�b�pИ��Ya�������ե�ac">�������O�;�w=#�B���-�ю;����ψ�v�T�J��8g���
P�k���}&=8���o1�iXi�#\��ěv��R�8�͢����^bfw;��	v��O����������F�ȡ�`�A�2�%m�RK�Z���C�Y%���j7��=�J�����m%	��8@��9���TZr�1�X�.��ۥy0e;�m��|�|}�U>_���薠Σ�¿�¦��V��L'	`/� ��K�m��4��^�����b�Fٯ�kޒ�U1T ���CK.�53ĝH����ٱ�es�clu�w�����V�G7��c�rC��9�_��+���bM��m.(Φ�<\���Q-.�L����T�����o�w{�o��+�!�qܟ�"��b��(�"
� *Y�����<���s��vX1�������0nA�^O���Ta'���O�/�η�Aq�ρL��Ϝ.g���_�(�?�rT��x$q㒅ln�#D=%�`i�Q��L�s�D_�n8�� Ř�\"���>�pR+r;�.��ѳO�s,}�o`���\��,�Ϊ�����])�e���E��Wl�R��MMach��lQ��R#?�P�����Wu��l���f�5���LN.��1�̈́m7ۯ /�����seF7(����� ��w��g��_W��$lڱ��(�׽��"��xɏ��=�����'Ym|Ѱ�(�6@��=�L�`Oc2�����X�B�]��bP�)�����U���/ft �Q^垺� ����D���mT7g`CQ٦�7ܿu!�s�~q��4gڛ7^�sd�d�i�������b�l��_�@(`#:��je��2Oʚ
�I��Ш�v�I�u�G�o�{a����x"�$���������E+"?u������/�7I�!�w���J=��Vȯ��L4��!���k�E�2�&oD�~��S����n��P�k�Og����^)�4v~s��������a�A�����D0����;; 6�9�#��{ �����j�m��p{}�p��֣���ɇ��M����I'�izH*�Z`(���⤢Ft���~B�)�	j���J�0s�{	^5�	<̪+���A�TC���Q7����^#4M�Ԧ�W�u��t�Y�ߣZ(�@�8����~/�S�=��ۂ3HD��� ���?5�%!���{~��Ǭρu��=�
����ǒ�0��@W��A M��M�	Cܢ� +
�f���	(��^�����WR����93�H��b!�XJ
�RE��������8X�SU�RXG{��=��^��}�W��3���g~s�ޗ�_Mo1�k�j'%��֤e�v2.��߫Hۂ,�wA�v�0=�Rm>���e�����Ă,�D�w���	��h[f>����
�"�]�&6�����MB�F�3����˺�eot�����'.�,�y�viܲ���:?o!��w�W@���[t�W^�<<<P<MD�]̈́���H�����F0�׷�U��֦�5�u��<X���t�[K���C�ξ��3����3Nöӯ���Z�F�N/�a�&s�-%َP]�4�?a=�h��;Y����n(� �����BA�t�!������x%	����#;��^iyiH��-6���t��H*�$����t�$��j&oa�Ap�lX����i)�{�X�p �`0Ƨ�70��Y:Lb��oV�I��G���s'�i�.{JԪ��:�1�&$Y� �vm���> .2�p(TO�8�LW@j��v3YIi��5(Z�#@p6mB:��X�kG�y�jz��X�_I��vjX߹��6
Z�/����l��zާ96M7��O�_���W&B�p�-.`I��:6tP�.����Rr+��:kDp���'gcj��`,w���;��W���K�k��<B��{.je&ƈ��h���?6�\ T���BO&;�{DM�E�>�GT� T#�\&
�=�7��?�	1m�q�nc����+�q��� iL�&�0G�ߌ�P�t	,���)ǕP���=��cC�o� ���4/��CEMZ����x}i��f�z��}��3Tڧ�%'1ؼ� �!D#�g���q�/yM�n}�0�d���Z���W����'a����(��3�=24�d�Z�ޢ���((��z)�Yv��)��3���T��EL����<��� ç\�_�&�;���X�{b�k*u�߁�GmK� �a���N����[�c�+<����8�z���_��~� �m�t37�t�ر�g&@��f>_r�P_/�ʭ�l�wDN�B��=��C�����Jf9�T���'���G9�{�y���c5�A2�@��Uʹ�x������.&���nL�c�����#��-<����i�2��)����2������F�A��ad���_c��M�
Q_�i\�=4��}��9`���J������ͅ�נ���Ɲi!j������n���k*�(��Pzٸ�s]L�7��/������(����6�)�ʶ��?۠|�F+���0��u��^g%��N�70�Jx��1��*V�,�&
`-E?��Ƭ/%r��5:ʁ��v��H^�Z�O�� �=�~S'��%��}�a�y��f\R�r�~K,�w��*�X�����O�tA�4�8f��3�/���b&�0��Ö1������.*���#) 1ɴ빵�We��,�EP�B�'k�B�n<�K���❏\�#"�7l�Ab<��P��'7�}:ߊ�	v7t5�UAA��_�W���d�An�l�7]�l#�l����"��L��.a�4���j:�Ůh�0ڧ#���8m<�+ t��Y��(��3ۡ�'r��I@�����_תg��}1�v����U~N��K����+Đ��]`9��"��������ge�v)�4��<ӑ&�9{5����i�s��ċ��}��<!c9�)�Sc3�>DH�-_�"Lz�X�0�w�uaӨqM}��Q�P%@;����<���7(1�^Z�'�X���h;#e�ܣ�ߛF�9�(�97h�^�uw�ʮd�y��i���'���=n'�˷���򂑫v��{��s.�[iX��s����cR���w��:���QE*�����u��d����^*�:ݾn�|ki����:ЮDoy ����j6�N��4��6�!r90�M��d� �F���ؔ[�h�R����B��,�`Wy��lt�h|����@j_�j/z�ⅲ(3>������������� ��P ������T@E�:��,H�#����P��3������Y t�;9_�h�P�_�\3��?d~�c7��:"#��}�vU2cVZ!6�ј}:��u괽ړ"7x8cYP�lVyZV$$���~���5tu�@t�O/���z�j�+�J~�L���e4P'�='��OVg���`�n��< ʱ��Čc���NH����ߦ�,�{�R��nEXX~4��6%47�m7���O����b�!n���G�#ώaɧ��k��f�8Pq�\ଢ��/^�ݦ�A�@Sw�x��J��0���;g��EwЂ�,~"��t�<=�P�%FJ��R��[:�^^nNM���o� ?4i:C�(�~D��T�H�4�.��(��^�g_�>������t�Pu5�ː��x��F���0�(��]�r�Ư�W��߁���4ހ��!BXpXf+�'�����u�̊�͝'���$�������	�`�3��������~ъ/��p�C���<%N0�cq)>�u���r�ӢZ��|x���Щ袡��V�ȶ�\���%��ź�*��2��8�<X I��ZV ����ֻ���[f9�co�&���_�|��;+�ퟪ+?�"�Cd� �����lGs�o��	Fm�F��_�⮶�6��HLu�Ph1� l�#��'<�0?�Ϋ8�l�sY�8o��?)<��U���]��*����8�_(R�u؀�;(��X	XF��$��I@p�h�[(ݍ�qmz�m[�cIyo%�����1]EG��e��
���3gW���
����Nx�d0Y���2��
�?�]�Sha~SE��{����J	{� Sl�E�ԗ)�W?��؍e�H�� ��TV���BP��U`(؍�kS*�"����iz*8N鞕��S�hu���?�͓� ��,(j�eph�ϝ����xt�](n I[��)�� ��'���	6���4��d���%��z�ha@���Sڒ���zzM�վ�[�3��5�F���z�}�&qȦ��k!�q@U�.�~�y�!8�ӵ��yJ���_x�b"Ɍ(҂E��~*��=L��(��^�ԯV��K�R�S��J���{�O�}����Oé�� �y��&�A�Pr�ˬ�<��'�z۾���f�F&B 􊿟����� �%��&͂_CC��_#���h�����	����Ǿ����׍s����zWM�j���mU�����go%�Im�-��IP������"g�^����N���;J������p-�a��by��hO���8�e�e�}��)Q���������F���9�8��Dܺ��!,�w��c�ȗI�䰭x7�F��Y=����bZ�}|�i<>�)<�Z1T��8K/'7����7�xD�*/��	��� ]p����w�(T����nk�45�v��g+���*�0����y��T�	���4{���$ʩb��z}
���=�/�5�6+!v����^�|�SŐo�7}v��?Vю=Sٚw�C<�u清��R�0ww��M|��Է�4���|�?xc=Q��j?4�i%���'h�'�tw��H�7�A���sy{�Pfi��z��kw�ϡ��8�6{+D��+�9=ȭ�y��h)1S7\��_��z.�M7}R�=W_��{�ŋ��t��Uq�������L�ݧ<��	l#F�#����!���V۔���P�rg5�%}���V���3w_�Gw}��f���3B����|��e&`�\�_t]#G�WwE��/	.��)t̻aIɻ�V���!kr�Aھ�,~�b�R�����A��N���]��GY�F"*N�oXI��#�y��_�O:��:ԕ�V�̛�;��u7�f"~e��8,���4�ߒ�Y7��zLXq�:���� ћ�}8�Ͼ��";v���=���Bw*J���8ܘ���d:˼^�$R���tz36�ʒE���%*��Zd`�T����e.YQ:I�@H�7F�@p�Ǿ����Z�̺WmǄ���-��;a7U����w��d�^�'�L������mS�y��qP���
m���v��8~Њ\�AпE�}νr�\_�+C�h�ֻ-�4j�"S& �e�YT^���9�|��׻����
J���1'�n�����(f�n4]Sk��4ұ�N!X�'��$�W7"�`�o����m�e�k
�~y��|���'����w]�&y���m��we>*���sF]��z��',>�ܿqJ"e<����y���G2�xM�y�[�4�L�D�%dڄ�t�y=3�)�5����~0�d��:1�c��y�HyQ_y}�/���ǾĠc&�����-�_���K�O{�]ܥyD\��	���� O'؏�����f�VoIJs���Yj�b7���,��.�.v��yu4����ȑ��_u6�������z[e��)�X����@�w���s�U]�*���\�)����[�����"���'CGL�N��:ӫw����P���*$�'ӷ�B��@���!U�kB���X��s��!����&����N�BT�E���� 8D���sM��h�_t2I��,�c�~59���L��jB=�~w�>h��D
�C�k�'k0P5�UT��9�� Z�M%�n9VU��3�. ,�,��h
h�OF��udstjb.����O7H<v��!�G�"�e��{�гt>��tgZ>�B�b�6��(+�QE����(κd0��eNO��\b9����G�j���Y)@�
/OL+Ā��S6p	�n���'G�0����p��2�����(!Ï�:"���l[��֬��E��/.%iӜ! ����F\O��;�k���nګ+U��d���ғ	�ѡAz¬��gժ�'�,f����L?\�)g�a_���h�r���!��Y���E�e���?'Q�D�y|�f�(�G��p�\<��s���������a�r��S,&�amٔ���M��w�FV�p�I�T��x&����?C��r^������X��أ�����d��ls��o��C/����菛���7�B�>5����uȝ;��$78��V{���Ԉ���[F�9�\��|. �,�zш�tg) v0%�?콅SQ���;wwwn��Cpww��������w�N�_���om����ULUf�{n�{���L&��Q�z��ԑ�����$gLƴ��TC�=�Cǩ[������ ~0]npA6�����h ��s�ī�c�9�u��|i��e&=Z�����,��݉Oe�l�yo�n>�^�'�)c?I~�쯱x�n�aRk��
��_e>�砸��W�Ƣ`�:,��"$<1ey��h�K��B󦭗�'k��ձ\�{т_&��&3�#�R���E���v�jh�75凿��ő�H�`�>���=�����j���r!U��~c��:aڛݣ��²��VC|6�]�x�j��䠻���U�g��ͮ���*C?3�Qۈ��(�`3�T9���|�]�g���^�s� _��r���˹��A�grnY圄�F�\o�=j-�@џ@��y̑RY,�A@�Y/[��Y4�H�d���3J�}J,ϯ]�S9�	FJ��lqjH�n6<q�~�A����O�e��s�9��CAs&Hn |�y��l(��f��D���@Inh�w����f��d\�(�_�n�#�����:�.�f�YeQ�+Y5���a䧖��Ȧa=��"W��p�?� �{�ʝ��j�D�ft1v�X^�iD�uGEV;�5�+��?oDl_��w��Rؖ������������ܳ��K)I���ԟ���Z�.��.�7�:n �P~j~Y�x)��7���b<<�-\6*�3���/��-�2
ج��TX0���=���-l@ki��_��!:�LI�0����i�8)�<�����>���;��5pC����u~9)�H�y��>���k�(�k�[*?D��k����)�6�`9K��ǧ��.��� ����P�y����
�.~{Z��x�������|��B�L��L[n�����-_��yDׇ]$6#�4�N'�ZoU�b:|�>�N :�2r�,]IP��0�\�_SJq-3:5����M>��6�.����m���gg0!�``�����W]!v���?y��\���W�����F�K��������0���so�Q�8��Ҟұ�y�*b#l�ĸMG ���i���L�#%��Ս� �$ٷ�%�˞9t��K��hұ��>p������GW1�{ş����L]�����q#��N�kC��m3<O�vR{P
��{t�}����ʛ=����K�(�o�&��C6�m͗^�=9 ��4B�8�0zw^ۡ�Z�y��c����ti��O�9��ߌ�<	~$P��6�C>-&����*8MY �!XG�K�&[��[�R��+?�J����t��]�o����)�݀#=�bHp���y0�YZu{Lܞ��r�r��:���BL�LN�A�&J�3F��}�ߛ.�nJ�«�Š�+G@X��(�<�e&�a�<��s��x8<:�Ʃr0&(N�4���&7��5�=[�Q�b����tRbٌ�C~�vI��~�$A�s�2�X���Ĵ�t?M�N'�wN���#�ҲQ��@�9���Q�}��@���E�ZIbw���(G��r �$MSS�+ ��515����MF2$г<�D��:"`��=X���p��qw� Y&jz�m[�����k���nh�\�3ƣn��F��q{~�ؗM��=������?Q]%�ڝ�P ��a\�7�NB0��Һ�px�������I��鋷�4�Zs4ӓ�,O��9u$�,}jr�,��z:� ��-� �g�M ֳ���ڄB�]=�������u����i�f���?}����y���f$��� #T��&�
h
CP�	Y����ͥ��T����X�_����y9b<;���!ƅ��Ɇ��Л��Ԏ��^��S�{E/�	֦�m�MFi��(�*>q�����=�Ǹ����e�u��
�6}^�����8Lw��D���lW�;y��`�����o	����Ɠm$��B[6�K82qk9��
7���|v"T��K�CKMs�X:a(�z�,NB�h w�
�ڽeԤ9xgRr4Q3���u>:��{ZN��1#�A��m\[!O=	�t.r��(:�l&5���wͰVvr�QS�j㤀#�z��V'ctly��B�������#�H?_��Z�,�حy�YI	�|S�Ѻ��<M4А���5��U��"��͵N��u�4ϼbCݮ(7K�Z��lyL�"��M�]?O,A��9��-��ƎW��$����A]mN�i_��G�l٫<o���U���W����"5����X��_�8U�ڊ�lٚ��t<��f~�:��.j�z2U��eO?���{?oٷr���%� {����s�ɖhQ�q�l�c8���8�F������{�i�ӌ��B=++�z'�
�o��"g@��䇪y�ε\�̏�o�ˍk���E�@�@�{���q���:,��Q���/y��̃뢶��˾�U�un}s�9XTx��#����bM~�'LՃ�" �2sʘ�Y�O�����ۏ��������H���^I�R�q��}�Ozkk�>2
��T��<l{�&n��7�C����s��辖��ֵ>!�5��;���(��N�9�>,�%�&ZTY�u\��OT�UC����H��������:�����SD��Z���"๒�ქ�*ґȒ��MLv�����s0g�sa��\�bO7�*�|���=W�T��9�4T&;6���Ph輛ޕ����s�=	1pР�jJ�������	�.�Mz�j��7MO�p���_�(�~[3�r�mz�QP���R GvL���d�:r]t�]=�eL8]
�F��k/#��>�uJ��O�L?�o�w޿}~�w/�C,)1Z�ξ�P��|�|�ګn����#�3�
�A��TC_:!m� 0@Ġh�>��� �]J��IewQ�����)b�G�y���'t7���	m�1�G��~d�O#1Z�N��R׳��c��Ld�{�z�#�ȕ4��3��	�e�i�6)	��ܺ�˚�H��"�W�|��B8�?����R�~nVL�Dا�9�ʺ����)���Cr�����#8�nK�*M�q~�� �����=����k�-�\␈�!�	3�x�6�oD��õ��9Pk^#7�� ��t3��z��\(x�&�-�������_PkW��T�G�?��e��P�H=Ij Nۓ�����D���$���7�����>k���^Va%�*��4v(�ʃDD���oP\�7�����s���kN��<ݝ	��d�b��v��/.��?&��~����$��$�.����|��%z�(��#�0�lٻ��_1�������7!za/�I0�+Ս�t(��}7�<7�(�x����-a�Ż� �\�0,��3�}�o�O���*�e�1��>C̿`�
�%&��Y�`��S��\�Ww�$���2~���7������� ��y����~'���<TЫ|Pb�1v�4�':�h��_J%wJ�T���5��Z�f�U^^_�i9c�8�W[�i�*�(�3��������r��(�gZ�x����C�?���-:��E��o�la�}�6Qy���}r���lg�(�2��BY����F���IB^��~�~���v������CՈy.6i����]z��?���Sѷ6��xP$�O�/��n�HͿ����d�F����NƱGz���rJ�aW��>������.y�"�s6��I�ƾ(o%�|��$u�?3�
���^b�b�����U�ū�a�X��� ���V�����c�Jj�����h�4���ͻ�"6(Þ��T�e��ȫz�B��6*��"���r�=�Ⱦ�]W�fܿ�J�O"�I�!�2�n1����ƃІ$wAA�p�0�K
���i���ڋ��|���t����� �����{)�=*�����(u�D�*�@V����4ޚ�d��i*��3����I�_x|�w���8�� }(�&B|�i~9,�y�s>B��m�����AC���Z�h�ml�N	>�ԏ�����-N�b8�Hx���2C�,8�O!�?���o�!�U�"�=�_?|���c�lY�M��G��K�lųf#�; ��d%`)����)rU�[��#/I"|-�Ӟ�z��|m�u9��(ި��I�n%�u�>��t��}�aiP4S�P_+�R.�k1��e�h��"u���}=nnlQ
�����M�.c+ ��a1r8�z�t����"I���������44�j$4R�P��*cU�'|n�i�ծ\�����γ�~�ZFi�m���{�'P�\� *�E����c�� �l-5 ����GB���G='s~ELH#��  i;Qid_ʣ���-�`�"N�n�v	�֞,cI���>,WK�����}&3��Ō\;��I~����&
�CO��G�i̓��(W�h���Q@��Yb�ض�Ѭ��C�%r!|��d�����Y� ���߸7K:װ	ģU�j�ǵڱ_�$W�8�h��a��]/!� ���؃6k��h�~���*tࡕ��vd֓�4�0��>a�p ���	 �}�*�淎���A�1��Th`Q�����Y��g����`5�~�4���sdC��5\��(�V)D��Udbǫ��M�����Z0��cj����и=�>�<��o4%����30����}�M�)��Ix�m���u�P�+ϥL��f\$�Qb�l���y�\��U�ce+�\�r���H�R���E�Z���߲�:E����ySB���F&����Y��c���jR۰|#l�J����"x���Ԥ������@4�a�2�[ �esU�~m���9���ľR+�^���%q��W:��Ɲ1���?�  B����훫s�CI��~x��$=�@�mK҅��p�t������,e㤀�1�L��٫ss�Y�;��ń��q�m_���wDV^�V	��I�h��u::��f���2���'����ҿ����"!>v�����DO��T�p�ɡ`ܭCT��P�!�%��������KT�?������>��πt��|4WO=<�GC '?�`G`�R���ĩ��\�'��2Ư��U�ٔE6�ku~�8\0X���c�]Qv{��.Z��7Ф�ߊ���Г��Cxku���H���zM-�o��Gn�-9�#fJ��!8�>�.g�=�P��U���u�\��ǡ��j�(VYU%�o0�$�p��k>��>�ԧّ]]��
�e�4Ǻ��GyԌ���Y�(A�c�̇�l!�n��G��Բ�J�>; K�/3���`�z�Fhet� a�͸�BDC0�P����Ͷc��yQ�ۿ�⥡9d�պe�n��Na�=o�i���y� p:e����ƫ޲\�oA�cc�{�m�7
��]e�K gU�Sx(̈Q<��3^A�#��I<D�x�Ah�3�1�7B�P/�V�Z)��H���53K�s�������G9��8�k#��	������=�y�I\�Pо��2�Xz��1hӦ�H�F�D��e���A��P��F�PO !�}#���!C[X$��<1HJ���P�^�[w>(��;�9��U�e����޲]ekz��LS�YG�O\��Ih���+0�Rrv	2ku�L�����d�[D'�cy	����Tv9�4Q�}pÊ���Þ����Nm��"�s�;���,A��b !zC�ɇ\����Sa�$0��e��0��V ��MX{b��Ψ�	�s%�'F��ۜ~Y�Nw��v�+P�t�o��~������_f�Ni>bB�s7�]zK_yC�H2ǂ�����S�1�@r0D �����N6>6&��(��4������m���zBD\��ZdcF�O?�a$pG%�~�[�'�*[�A���B�W��,�ֹ��|[RD.�ۅI� �@��R��]Me�/?%�
Ο�����:m/j�H�t ���|�m:�c��K�$C��n�Am����,�
��Q�5g��a3�*�y ˣ^�<����o����4u�Jk��y¯T�z�+���� �O67��{��P�ӎ9�W���O%~��gݶ�?����q /����@��W�>Df���Q��
����A��b<Ue����k�¡�j���^Nf��쵲-�Ɗ���QA����N�jg#�K>����t�X��i{�K�mmn}_���PFP�H0)��!TR��I�c�DB�?�!��훼`�*��Z(d��[2:�<C���i�,�[. pʠ�`���f��\����r���H%����z4�$Rk��0t2��R^kj�M\v��B����X���\2��G����>'��}}U�����*ᓽ�}�s�	0�x�4�X�NE���L�	׻�~:*ۺ�W]����L1��.�����Y�t�	~*cRXf��j�����Ow���֮��o.��q�ႱB�?�VU��G���xL}���.#��s"��y����1�AP�io��KƜ�a�f��Uj����������A��~b���Q=�=��l$�[��o�s�݆�vu܄������V��I�$v�Z��l0~!6�x	�,��;o�3�$����-����0�ZR���@f�}��y,>��4�����Fw���{L��*Q���m�d2C���I�ۢe|i�&D{JP�TT�"��p�u�j��{�a��#������K�YX���5"�	��]�&/V
� E�9��T)8�Nguv��;
v�S8n"��P��tnvu525��)Ƴ����$�19ANm�{K4�K�����l*e������<�]���)N���m�TC�2&��c�YQ��ڷ^�X	���n��Sݯ'��M�15�>|���C(ӕ�,����֜>M�$����+��^I���P�MFG�Ҍ}4��@=I���eW�V������q�>��f��-I������0�V�)��&�R�73@��=i��Å5�#����=6�Ia�&�GB����k��&�8s��ewf=�<����>�.�.��z���������G���u,�=6F�����
@:ʣ����|����w��h���"U�T3��=����qs[( �N��	ǫ5t9K��r�y�Z�_�*�p>dz�A��Tª�\�������p]� ¬'*��L
rr����p8��6��Č�����'��n����]B���/�ZG����d_ա���S���.�n��������!� ���T�N���kE� �>Zm�r�����"82�z��=�ҸrS��0=6E��򏣴D}�U蛈r�/Q�M�"���D�
޽o�u��d��/�gy��={��@u��8�R�!�9j���ULN�+f�񥳆T7,�p�ݐ� �0%�S�~h�{4/D�*v�p�-Ħ�G�W\����{$D̉���zr/�Ѥ��0/2�.�M��\J����wϖ���R���m����x��\��d�52g�X��-�q���@��~=���ɐmŭ�㷣��W�k�=T��!@>��L������wih��M^r݇yC(��!{�o�D��,J�}J�`��չ.�vI��j�7�˰�������R�}<������	��v�õ$�/zW$cM�QfD���v�mF��[�L�F,rR�3�-��ݣ�y��h��L�����Op�^y?�.��-��N�u��ۮ��S����"������ˇ�1Yd��1
m����E)~U2��0ys~+d��O��c�#���Qc��Z�,�/N��b�:������fGbO;���x��+_0xZ��ey�`��E)���W��:"��@?@��=�@�vʇL�0v��}V$E�_\=��M�.h���!�2�#xx���~�}{�x��Ӟ�ph' XN��{���(I�18j*�q�@b���|בf�J�H����F���Df��D��k���%�TuNߏ΢��~���WU|.6H�|�1�"C��ߣ���Z$����[U�H�F�Im݇y�T��͐zU���P)O[Y��<r
��[���Qs�K+�b$��W���plǞ��>��G�޷�9T2C�i+�{i�Ј( P�	�C��@=W��5�^�NM�w/"a���L��ߧ30%$(�a�eЅ��\<	���s ��y�����̕��ў�J��>���)"}1*�l��`r7]�#>v"���$Zӊj:���x׊z'��E�AR��"�y��� O��8e��Q?m���jq������/��L2H4iP�Ucb�	C&�I�GCi:4
�O�	��q{���ΐ����T�8L�yi�%A����+/6��[�s�
�.wFF��θʵ���N�& �i#B��Q�$�h_�e���n�A����[��[L�<Z|���c*�cf3��D�aX��[�1sl�š�8P��f#��j��N,Y�8ś�� ҖY}�Q`h&��JAHVE)�����ʮj��~		��X��Ҭ�@��h� _�� ���]�c�o��=����ׇU�V߃�OŲ0�nC���0��9|�aD$��v���R��U`zDoI�g
q+�ߴ��.�����08�:�K��l ��\?|:����b���3����1��[ղW�P��}%��	Ӑ`֘4i��T~��F�{�Nd��f�b,��y����Q9�,\u�b�^��� �SիS�e�����q�ӭH?�T:y�����2�on��O~%Ű�i��e�'���u�ޏ�J]��!��FÔ U�݄(�)�_Y~d�y�~���� �M7�fO����5�k���E�,0�ׄ�n�w%�O���4J�x9n�(6���t�ʽ��m��[$��O5�2���'�a�`��%�{�i���-C\�)�[������F^񩵆�Bs��٤`�;��Y�S��-a�'����?t��I_���3�"B�����@���t����=�x ��f������c
C�Ph٣�����+�(^]{�"\7qUB�L.=�t��!n��/��XBj������(R���,^B*h腽���F"�~d�8U{��!�;7.r�����虋��܋��y9��A�Ȼ���H,����ݩ�dÕn������g���d����'{$܆i��(��b�<R�/�����n-��g�8��h��
��k�I���r� |V3l������b�8�ժ���/���G˴��6`QJm�xG W-p����遐���$���+"��� �V�jg�L�E�k��h�Uv�����i��4Q,	���D�
Ս����՟\��Y�Q$9x��?�����tZ���"��MFh�j�N�J��^�Pd�$\7g&������	����,�����G�8q�d�q϶��s uk==�@j�p/��ׄ�=r�E��6���`��H¬��Z8b����w�Hp��][
�}�P�^�wE�����*x��:�ɴ���:.Ԏ��j����GE�~=l�)�O��Ճ��^�:~���x/r/>���A��f+S�fѴ&�_�K������s�$J3d�V�im����g����B� 5�-�ǃ黑)��:vݻ���;����"v(vm��g�E�������%!!q�:�%qh���'�O��ت1�F���<�g���4�Ҙ;�^���l?k�&�������{M����u����ڛ�;�f%�#`�O�廇���m�?�&�n��o�s���a�h�D�/&�� 9��}˙[��z�CD[��~B����z�~qk�W��'�>�ZE)�;kV��]�*,-��@�3�5'���Q�ā�c�P	����y���/����{��' ��l�B5�����X)0�T�~�"+I�n�%`������6�ꂗ����-5K}/���V{lIT,\'Wυ��c���w��ᡄA��\��_=��v!�L��Av2�x�q�&c�E��z��� h�Q������g:�Z���x)����4��(��K;y�R_Z~*����ϟ^��0M�%�ǀm\�h���U�	��g�����m&ie�p�Qi��7��  o%$L+p�9��\L:�7�?.3BH&�(3$s����]W�k,"M��i��Y���w�C�Қ�fJ���}l},������aQ���"ܲ�����FV���5B<�������fȱ~����/��
���b��B�����Rڐ��)7`��ax�@�z��<�D!9�lI���,|<����Sx��.9��vwaF�<���<R|7�3�z�u�6@=F��AZ9�04��@Ri�L�����7�ܜD+�E�#�N�E��!x4G�f4FQ�K�-�NhK�p苅œ�PA<�
���� ���cKD[���K�U�#�����S��|�i�TϨE���~|���9��0^�����n���W����N$44�� �g���@f�	�V@�4��Bb�����C�ח�x}_f6L���O�?����(ܷ�f�ێ|g�b��>�Vcu���ͥ�-�z�]=���ҵ������Pm�a����k�ə�;�=gf��nֱ�]! }�����l>;�M��钴;8�R��TL��2����� .��U�x���`��N�B$��Z�n�]���������7�V W`�B=��}	�^~1Q�#p����]�5�r4kk�I��tH��s�0ؚ��C,g�yY�������GO���<�$=�#��0�h�L���xF�~A��y��q�h�v���t���E¸V;����W�㕷�t�O�?��*�c��Bh@f�/_�;�xC��g�׍--���q:N쨳S�V�n�2�\s|�|�1�w҉�Z�ъ��1�q3!8�Na����
���	�bi�F���	�~��Q_�ߐ_���U����ڽ����SbX�u��2��k�������|���~lޣC���PqRM�����7)P�%h�z`�z��Jd�T��ӹ3�G�&�f���^*B"E���J!e����Ag���c���׎_ 5N
_��� �]�i�1���1)�O� U2۴�)�ڂ���[856�Z*Lҽ�q<w�����;������H�f��,dT��@��'&��{z��A���7���N&e�37�l�䠛�R�blڡa(����˩�D�y������]1�̱���`+��EU���/L���g�v��������B]�#O
�V�4�wi[�MGG�'��E�@c��"6�5;%$�~���,���%�@��>�J��	���7�ǅ��(w�����4�;�8y��\3d7i��jr�l�uY�y�^��Ѹo�ܳ?W��c��Y��wy����{�P��u��R{u/>���ptK���ܫ9˾6]aw���U>t��|rIFN~v6�1� $�1�fw�%I�eU�jzv��W�C�ѷ�vFF�Խ�)���#�E��dK�ʔ1VW?7j�O7jRd�$U v�>B��>;�}Ffl�qt^��ޞm0��	k�.��t,��,��3@�{Z	�i(�`��l����ki�&	)���7��htX��t�<F��/tG���o����/�"EѪ$
�b�;���Ī�ٲ[�ެ��Wj��a��=@>��M0�U����8 yke�&�	�&!��|�e���p��;�-	�i���65U�Eݦ���$��t�L�S���BNrt���������CC9n���@��m��M���o�X ���.B���u�^���f���c��vLg<Pg���?�?�`}�J /��bto��v�Ku}k�C��}�V(Ka�d��T�E��� �	�cF�O�A�w���<k~�ĉ�x�z˵�p�]lc{��0�����B�Z�2!��-���9���ࠎK󠵩��RN��<��]�bv�}E�R%���Y%��t*U�B�V"B�	b�x�fζ*���'�5�	-����U^V�TN�0ܸ��D�zq���jDϛɌ�nWʦ�T�
_�����+H���uF[�9��7���a�M�f$�Z^=$�N�)��cP��|���I~�{�B{�}���CD|�y��/�}���>�^����o)CKs(�B�xb��?/�B��dq*�	�<ЈMH�����247������w��ӄNhUyX�?>�R:o7qb=f�}�O�r�'�?�`P��/�DD��HF���/�'X�HgDGTob�7i=���s$(�{�zX����������)�9�"����#? �1��ْ(���� ��&�)0�����q	@���|�i.Ed������)qn;ƷN���r��L,i�1����9�W�u(r.�� �:2eK���r���2[��GS��`�]T3r����=��f"�y� ڧ���� Ǌ�%bi� ZGi.�1�K�/���G��{PB\"�������a�~��4R+��� �??�:�X����}��W����x8�����tpȋ�=S��������M ;��^����"�A�����Md�i���"��9�m;�3��kAT��H�a�׋���%i��]P��2�f:kg" ���1���T��R�rUV���ep0�6D�$0C7z#�qC�q��.�}�`H�6�6�6�^�K�Hq�P9�H=�9��"�{ZQXLgN����4Q�̥�z�˪���[�4Ef~/��<`2X�,7\gb�q�ȉv۵�#���8)�Z�D�6�ѵ�*��KR1r=A��fP���n`�_�1��[���r�.�{&2�ZKe���f*(�����d7"�.d̅�udUa��b8�����h��Ae��%�y	tR
�Moﶖs��\��U}�Ȓ
6pH�He>%6~�숈C!Ö��ɛ�F���p�4=�����W"�;t��_��w5P�c���R���-$�DP��4��ܻ�&�:��2A����e=A &JߒM�Q}�Qs���F^7W��f���~����"�*��������e`�fR�Ҧ�����dd�6��&]�����N���Җ�ܼ�7;;Vk��j������H����\���P��Cfr�ӌ�	�!�D�S�J'^��E}+`��!��0+��B��
"�~����)mq��Q�aԅ�q��Q�3�PA�0��n��F(�^.�w�L��T�>�` U�
Tyg�ւ��r.��e���XH��֒h���w~���So
�J�>�S羋�$WX�g�P�OG#�C��W���H�h�'4���08��vO�^���[
?>��싍�s*�J:wOu�qB^1�w"�?s&��FZN���a��4Svt���(Vr����Z�� .
	��S�3E���b:$�)#^�('5޳u�bY:2����0jJ��x|k��f<z���դ�����U��ai���^Z�hp�,�1I	�z��#���I8
N}Ӎ��):�:6��x^���J����5U£�\uqV�u�'��4;YL�e˰�2"ٌ�碰v��Ո�#�/�qXa�3�}%үU�4��P" ��΢�\��-�.���Ǆ��;9*i��K��.�y:7�3`0^���.�)n�ܔ/��x�;��R<��߈uq�/�>鰃�UxM���XK3T��0f���72���>U#.X��↋�@).�*�c�a�S��	ӈ�fd�HD^������]{�!���1�_��x�wOj~h����a1OɔB]���R^^�Kq~d[B�3fa�51��3m2��)������}������W'zW���@�Qm\��D/|��[h��/�1f��aGؾ�Uܤ�~/��F�""H�՞i���PM;仄��.���l�4'Ǝ�̿2��~�m1v�'��X�����Ĺ�����'��,�"�}(��Ӟ��܁_�ͭ�)���D?����&�%cik�eu�2�`����[
����Yw=�_���׼����j8�Q��$j/�Az]4.'�y�Yk>�}��ώ�N��Fލ_�^�aK:���5B^�G8�V��2�B5����!��������ŝr��_��U��я��£���=]�T��)�F���x�U���c�����18�!B��g���������!����*N�V.�(t44���v7e�t��:|����@�~��8�K
�&�#j����zk�}ԏm���A��8T/�`F�%�ȟ2����Kl]x2�y�_�B�9��,,�e�� j�De�Ķ��uS���E��ĴM�6S nK��`���������8q�*0Kd�MdO��ڠ�[�>��ٓ�C��L��H���j\F�H�oI��1�yBF]� ւ�9��a��B+��X���f����O�g�J��:����AR'�8�O�dv�K�6�׀੤�UG��Ң�i#좈���(�9���,z��A���H�H���XxA[�b:v�gU���7�@����r�OƔ���$�%h����I��0w�M�Rk�7:#jyY����q�D#�$D�.��q�K;��qAy�B��$CeW���%�B�r��]>���$vI*u#Io���tȮL�S9/��bg��Wzy�/��j�h+R̅�TP��U�@s�Gē�4[[�;'2�۞[�aqJ�9��,|q���'���[����E��b��n1n�P ���-$�4����xn�*L�/�Sm����S��t���d''i%�K?�L�������Ȧ�Cv��P\�l,�C��a�fQ���R�u	���J�Ϭcj��^"}�I�}���<vP�Yٲnz��FRx3	N#MI2 ݧ��$��	6���yР�-����v1ҶE67æPX�<���͜�DCભ��#p��P>2��c ޢR��P~�XCv%1�8 |:dw�����-П�꭛��Ī��2G�U��S��lm��5X�����56������̾�~��&��ɚvCw���r�H8��B��*��eQl��Ҿ�k`��r���!�U�$^�S���f��t�?WG��]-.�f���v�U)��GF��yho��x6�l��FEX��[���Z�N��fU��� ��Z*�AF�s.EL��m�l#�2��T���_���
�Cǵ�ɀ������Y��q�~1�U�{�g⁭U��`=���u�9�9� ��g���}7'�||'��Ѱ�_�A�Ffl����b� �Gb	��.YV�.\Y�g���v�J��{l��1=��zh�?�e[L<�j��+p�)j�C�,<W% ���43v�J��g/ H*�՗x���"ɟ1�����/��S���ҺdAg���i{���OVR(l��i�I����)ݧN�d�s?J��3rH�<�:�ȶ�)>&��4p�	��Ē�ԉ����"f��oI�}Ѹ���TEH��������#���Af ��j-۲B
7�*KN�^)�e�I��������!ŗ	�2����񹷙^	ttC]c��S�_4}�����5�t�L�^B�H9jz�1��Nݟ���;�y�w�kF($PP/�p���T���Q��~�!W�~��&-Fi���ru��� �4�����=�Y��z�GAHd��خ��
�%��L�f�*M�_�q��P{�D�H1G8!Q��{Q[�(y��ޜ1��)�8[����"��q=&���/LȮ�\<��S�OZ{�<f>���h�7�O_L�_N�|žRq�֯��Ame�KLh5�q�U� ��8���V�����JS�k+�߷LLj)v5V%�~QE}��m;�@y$6m��_9��K���瓺=��g6�A�z�pv�r��H�А�� �����e~�,����Î�W�O�_	Ni˱d=��*wz�Gx /�ۣl�6�����{X�D
�%A?�c���R|�-�������}�Q��>�~z������6on���,�7�TY��՟+�az=a���"<)l)��0�t�q��U`�lk��:�7K��,)I+�@�g��gK�j4�ٰB���U��>�^@��p.M�Q�	@<�s6'y{_~v�5N���LTdj��D��:�`�����T��ݙ��	|���{�uNs�-�,��lD��Z8���}�&R}i�C��v�8��<��,a����klO�kN�zx��%1nW�XW
r�8��i���q����������k���M��k����ƶ�[�b�\�]��L�c̰LO�f̏�$�x8E����</��%�MW��M�
�ǽn�O]�^���;���q>-]��Kc��p�Ih�z��:),��@Mp��,�����ón����<B}=�_�z���4��j�J�����|6P,+�aɛSX:J[B��[�<̇���^���<�	���3��vD^��,i�1�@�cO���FUtI����E�V5�㖝��Y,����{�P��������6�s�'9=���2�e��C0�Z�tt�[�s�ŔG�h�L��?��串�&�z�N4=���y�1��z&���P�B�D�=��n��p9��ha@6V R���3S�u���Ѕ���\j���7$w�$ n͐PP��t�����\i9�8{�� Uu3�9ώ��0�2Õ�� m�U�ʭ^0U<�9�ka"�<�ʲ���P`5����	(�ٵ���hOiu��T�KR��3�[�~���KA�q*E�����f�$����@�]'�t`6��!��b��d���QNn;k�ʁH%CèJ�?tR2�0���\�&	����S/ȴ�������7r��7����A4�u{��H��M���׉��mGh��t�f!+6�v������F�ϙ��\�)=��;��6��gi�Fc����6��'�@��U��,�RQj$}�c���c?UL�F����x#�`���2*��Y�Cp��N����C� �w܂�{pw����ݝw��z��ڧwuuuk`���ޙ��Dٕ_�&o���m'����5��@�b�)n[#^6�ۈ�� ��C��1����cps�&"(�3k9	���(9ԋ�Cz����.Q�0�!���*�v�į
Q,��B�)^���Wz�ݡ+ib��&�_̷ܺ��v�\s�!��bY>�0��6��g9�KD���%&��7��~���WMd`���/�҂j�����%�Y�>�s����nM}�Q���(�B�3�u���7A%�Li�߰�,nmI<B�@�+5 �1�t����g�����G�� �d���I��*b�u���;����V���B��B>�A ĉ@�~�B֓7fQto�T�-gIk��i�
�VT��oS�'fh���GEӇ�p�fq8_���*m���P��2�����:ŭ�r���7�WY�q_�1��%A���3�+�������g5�GW
����cjQ�Z���ʏ�;�!�s�_�r��xB�e*ڣ"R��/m`v��$"���8�hׇ��m~�B@ ��(�2ÃmN+ݲ�K�٦���?�l���|(Is6���L��?-�'m�I���P�vd�+U������gO=r��/�2��YـMCd?��?�����:���1�?�FeIhO}ܡ	�,�Lb�c>�Y-'��jٗ���|���cf�Y
R��F���T��$۾��\�tD9KW�̂&V���_�d�B��3G�r��׺ i�	"���q��JY�1��Vat��dt�ڱ=�1����];NY?��un������J�L��7��'lR��0�w/#g���˝J�p���T~
M'a3COR������q�j#0��[�=�<ϡì���)�]Z�v�L��c��������R`�Z�ؾ��ZI
 ����زA�a9eS�Də���s8�`8�⮉�9���KR�z
���Ք���J�����{�2 MיFf�:����o� {eR�veK!2ו����o����o�H��\QY���%�?���3Cp=7u�4f���3�m�/��h�Tk{��v�rR��<"����MۇK~��w���dq{fB�=�Ϛ���R��v��sЖ���sva�I�$P��F���>�r�p�4�/��
��Ci�������V�@a��Ֆ�#�|$�ԥ����G�Ww�ḇ�?��Υ�5�V�a�#��fi��3,l�8�`V������n䭮C�R}��/m�B��nSp������� ���	���^j͸E�v�ft���:�V�28�k��:�R��RH4Q2S��G�y�2������hɿ�Bsmaͼ�r)���G��rk��B�2zO�-��3\h���~_�E��P���H?�~ݤp~�ID���!�'��E��K�zj�Ioa@��J3Р���QqF������wIU�D�C��_o�������q]����!��(u@��W�Th�Y��x�r]i)�Eu���.��'������'&��=IЖ7D�"�1o�Ԣ	���*����.��<L�����X�����c��u�������>a�D�s;>�$z�8�x�p�Z���d�U�M$���pA�p�`<֓��U�I�r��c����4��F2�޿f%��A�h�%��`$&���
qI>��C<!Œ�a�}']�mG~O����D�a��8�x4+�i������KoR��ٌt7�������;�Mq�EM��fF�h�g������D���5�-��sUY-m�},އ@eu���ײ|�$�m0�@�[ۧu�Y�����!*M�c�#\�t�z�����Z<!f+j��i �\���w��,�� �����ŔX����#C�ϖ;>d�2v&��5M��̛9G�2H(�[x�;di�ޗ8������Z�����	�p�3�[�!س,|l��{�c=S�L)��ٗ9q���hD����< �/�2dRu�1o+�:R6W�@w�����lEN<�=�i���,By�{R#�@u�G�4�/[%�}ٞ��
<�L{β(u�w��>9W�=)*���Y��<= ��݉�]-��N�B��@� 
r$����/�p�0�_���@��0�I��y�*BD���4�������K{�H��� ��;��Ә]�9G��U*��-H�F��at�eJ0V�3�P,�e+�k�5p�G�G��Ro��G���q�ύJ1�x��+� ӫb��(�Mt� �n�,`�`
�u���eN+��
���eG.������~��.���6��E.̗�t�#�\vi{5:��H�Pщfc(�o�W�a�׊�������Mu~��;��
���/���9L�g��J�!Fa�7��m� ,g��� ���w+�K�i�!tw��+���4]����K��V5��w�'��ЙwP��2?֯�aY��+KbH�K.�i0BX���Hb|S�X,�+��s�K�Ʃ������}C����gk��y�#���M�
�vu#�(��EK�B��C}�Y1��U��ey���a�4���L�Q�3� U��F��{�S��B���a�9zdL�R���l5Ȥ!���b��N'X�ʈ,�=ev}EI^�(��w'��h�z�O�����n�n���$�qkaVV�hp��H�i-@Sj �h��z�`eH�w����Q���3�ԛ����������b4˂)IO�b�m�`��	�D�
5��|��l��E'@��J
�`:"����U��h����4��@G��%�{p,�����3�w$k&s��}��G-/���W�a|v��8٦���e������g�3IhMY�#�dQ@��|����C����߿�Z����[�)�(حЎ�/ ֟L�:���R����5a�Z��ڑ�󁬡��qm��0ց����%�H��LԮ2�XK��Q�#���b��>�o(�Lyѽ��yA�oq��' �^�l���}��k�	6���9���6�%��qr�������SFr.|����;�e�y3�W%�i��Ps���NR�\��ý����;\fԽ!�n���Dm����q���
L&=�V�e��m'3a�/������= Ɂ|��Ky�;��[�����>[�!��/�k������gC1�&�S&��~�kTЃ_�j���@��#��ޙV�)���.`02�[JB	<Qḱ�ЂXh28g����HB �&�O���e�e�
�6�\N�_����7��	�}�|��?8{ʗ��!:f
���"��-#(j���m�hk�R�d�6��OsQC	�h���G��%C��)]����k@X�}��H&[���{��W�Gx���M����F}p����ŝ��T�ࣜ��R�JU�Fk͞{�yS�V�,$�}c�=EJ9쐲-��k1'N�W�����N<�Tl�1;���^��9�bz�F
���x�� ����d�D�'I�ߗV˜��aL�UOZ�����)I�;�X�\{��cˤp2!.%-�9V[���B�@��Գ�B���d �``��'s)�e�҃�S'R��7��|%�[�4q�L�DO�F��&�p�U��0bQ"qoi��ab%�֞���a4�ϣ�Z��`�n�l�kY�<P$ҋǙ��N����ԉ*.�W�9���jd�[��䶠����`�j�l~S�K ������#k��NP���&'�Vrk�_cٷ|�fx�r�����u���?�;�LlE�H��"Q�u&M[$��U�1Id�FR#nep��`��f+����VP�l����w��]Y��IDsH���e��@�i!�������5��֊�Js[��`=I��)������� �H������E���������*AΊ "��iؒ_NJD�k��Q�#��&�R��������D9V��#˾}h,l����ۛw���1ջ_�W���1<�_��5����[�5&���p��0<�;���ʸ)xL�F�xt�|Ғ��<c+����]�;�Dp�Ģ���S��S�0@������vr���__y��N����<!׾|�vi�j��#�ҦL���/�T��c�i�"¼�-�<���������h*�׮�_h$؆�(���lۓ�m�Y�5}5Y)zݹ33\7��%S~m�B�Rr*���b_[V��Tx����19u�	Bv�?^^_?U0���^Bs';{y���5Mr���2�mƝ��"C`�G�3̐3"�������%�.F2�:<W� �No7��T��d֛�q����>�e�����۟�Qu�A+�gռѻ�е���'z���-_�~ҽE4X����c8�zC��9�ڬ[��N���B�_Zm��9��7�*�����jy���ps� N���UN��))	o��Z�5���_kyX��<�Q=]�O��(�B�	e*O������-��O��G �M��n�e3�t��X��m�� �T�����'�ڵnƽi0�8<�@�����sټ�㒜/C���w�$^S�#ܗbr)��c���<�
�k;�gkm��?L�Wv�o�f�s��N M*w'lfY�Yd���k��;��9�	����q�\�b]9����^%j��E|s�^�ʛ&T�Y?�\ѯ���#��@�|�ժ{�9�)2��4x��KV��?�%�`�y��r���"�˂�xȪ���x0l��iu{0�G~�
��O7��i�eN�;�	7�&P����	8����⯉$���83��=_C�XY_\�>�ۗ0�sw���6��1�ָ(a4��P��W���ęF�]|��DӉ�<X��j���.��h�<�䤍��RK�����"�qb�AZ�ҕȚ�[�M�ȕ�5����傫#ǻ�g�7j��s�����"���n�k&��@TDR���1�����ʐ�jƗ��(Ѯ��	D7*Q�Ym|~�}��B��6VY�N�k ��1&�6�Ã�@��2�}_��э&+�	�.����f�~�J�QuD��-o�]�����'�Y-=rϪ
Ő7�!^�m��CCf��-��>A�alEc���P�(Xޑ���}�mi��:�z�⦶������Wt�#w� ������S���z_r`(�g�W�Բ�������o�o�4�O��f]^g�jHxr����+T��]ɟ��/J���
�矯ѩ�Z�/��O��܈^�8�cTO��2j��:�*�75�ǵ�J����ݥ�G�pÞR0C��1�T�&�Eҵ6V0֒�|s{��.y/�_F�i���j��P���^Z38@����s\�i���W6�*b� ��'�P�f�����{�N�����^q%OC¾�N�V�̝n�
�MV��k��&0���{�аj�i����iw&���B�w,���pZ�ø����H���34�*�űq��F(�xUh��ҒχǑz37�JT��hn���i�K��7�-�� y�B)�J[!�������/j&�X*#b�ރ�6AƷ�~�P�����۩UYj�3��w<�� �U����$ӝ���W�m&�4g�?��[��D��8͝p�l&���c�ɯ{���)ۇ��|��Rb�3�c���2�{��\F���ރ< �]'w��ܺF��&�{��b�Kp^n�r�N��F?��{�$�9�S�>�u�2�����Ւ�(��#�Ņuچ��@㽛�R%+�)��[�Ucc楮��-��k�l���id�pw��RiK~��.����M!�V���-mh���?�	@/.2
{xR'�w������}g�G���U�S�^c���:8��
4�L�jr*'㰞:5��:�9��+�?��V�x�j*��P&�	X�w��F����V�=��0�U�����yO��	���<O�3��{�uo��1?�c��5x+�_,�oN��6�9�9ۚ�����ʞr��SWe�=ފ����}J^�Ĩv�$�c���d�B�_�E���g��je�����(�X����_
LE##�2��+{U�~:�dS����{���ׂl����q��_�m�	ϿZ�� �+^��E�����aRn�|��9�u��rU������*=��I"�N�p�b��ӧw����ot�n%���@R��$�^N�&"�J�a���~��I �v��(H[jsn�����1�x�`�RВ��1�1�`�)pV�$�t�Z8PXz�	(�8���j�u���H]����ԁ��O�}x��o�Gz� �0���v�K�Te�piz�m�N�C�u� #uy��l+KL�ڜ�҆�^�3�:Z���1�PL�{c��+#��H�ac����1誊�0b���ï��f�p���o.�逢�F9��h�j��<<�'w�fl)����r򻁳�5��س�^���X9T��ޟ(2Q�cϵf�����zn�S�W< ���*���g}c����
�{�#���Ik�T�)���P�b�e��$WLw��=��_!�������B�%�)F�ò�	WU˝sϟ�O��}\�GL�O�Ԁ�oi�|,�PXqf�ˋ���J�3v"����o!�Ih0�SU��&:�\B��ʙ}=m�l�o;[��'XS�Gn�Œ�-A���[J�\k����R�H���&ZQ������B�I�22<�Ω+b۾ln�/	���n͗D,�VI����p�T��Q�&��5����s�5���g��Uq�K2�Y�R��"���K�:���N;�,1��	�_
ܰ�)�零��������L�@	yl�������
�+dC8��p�rW[yT+v/.EdF�	�#SR�8�쏟=hq"��:"���A�Zur��gQ5��1�nq�t=�4�7�k��b�@o�#�L�z8�^S�����V���M�'P����Y���(BAn�4�*��r��fpP�˭��ʅ��e뎄mNې�*�D��oz���=`.�@����L�֛�a1����:��x=�L�Y���}�/'\�5���۴S��5o�07�M[N���ʹ}d{�1�,�KH���I��\�Q��G��d���ʶ'��R�m��$��M
�jMk�GJ;�g�7N�k�}3��u9��mw��Ae⭥���=���C	Sy�y,��o�2��G��&dG�΄h�� ��*p�*�b�F
�$~�������퐮-E�0B�Ksw�����A���9���[a��5�u��������j{���-�57�������4>戊�%���C������ν�t�c.�l�}���?u�� �*�u�,���V�|�>�
�Dw1zAr���Rn�s-��q�_�)�&U�f(��Ox�	,M'&"w$B���?�ޔeyC��8m<�:&+�ff��g/|���˄|�9����!"�r����V�+I5KwN8�K8����;]<��]U��w֫�zb��������(T�v�$���R3p^�e�Zᵢ�Cc"3Xvbh�v^��6y}`*0��ص!��g$p2�6�2Z+�Dv*b�/|��wz�yWY�������h��8q����-���c�#�^`6<�5@�}�84Z�[@Nq{�5K��(�w9� �IY�x�W���~u��;��>�9���+�fZ�J>@�����ɥ���M�e���m��@=:���*���|[T| �ko;�r3�Z�����L��6?�'�ڝSL�k�h���~��p���1�5���k3�#��e���f�qF��|��sћ�$�4��i��Pa����/u�ʼZws��ה��Ɗ@pz�<��Z�Yn�0���o\��н�@�=]JV��u_����͹R�����p�����QU�Ժ��g�X��6R}�Yb��q�a�;J��s�	��+Z�\;���`�y�mi@��m$v�膩 v��'m(�Ȅ/S!gUcSsښm�($�ʞ�l�=Vg��Fo�w/Wo�{��P�8�

z�A�u�uP�w�	�/!oQ/�7�g�����B�����0��9�G�=�L�r̖�B>v�R�" ���6_r^��shm M������T�ŔU���:�텠;�V{G�^s>����1����=h4��j�]6Q$���k���6�j%��&�p	��tQ����ls�<bx1��,��|��ᬋ�P��}��vߎ!��U�9�U?B"�:�@�^��g������j��O����t����%Go�OD^f���fy�&�O�Y{^�(��̨s޹4������	|�9R��tx���:�����<'g�!3���E
�HQ���M�8��
��^Z^�%`�NW<��\�聥��%ʝ8V��f[Y1�ҮԳ�ġ
��ښ��n��R� ����V3���?@@eI$?o��їP������J���I`Լ���=�=��E�����՞�a�����p��<vU������z��S�Z[1z}���܎q�Ųc��$Sd�=���"�ʔ����!�6��q��0�W]⧊#;b#`A����n��d�vh�Lr-/����5I�i����1��*L乘�"z��z��8�����g]/�er7Mjqۮ|�y�W����n�\ƽ��N-7nL�wET�)��\�o�W>��|ک�D��E�����;K���\�7�T�1^ӷ�<ˉ�Y���F����X�=����l��AWQ������y���7���ũ�n�j[��Q��yT�|m^���paBZ2U�]�S
B)�y�I,,xt4~M����Yd���|�s(E���	�J���X���3�*�'�K�z�������Hw��%��Lkȳp���TSXc����t�/K�,o?mp�;[�Ø��m`��+g<g��:%�h�� ��{:���/EM2��c����2C��� �!�?�s��j�65���
����/���U�uD������bl/m�P'(��>�}ى8�]q_Y2��:�����o�����հu���.5�ʫ�x����'�����¤vu88�"U]L�;�c����蘭��z���W�G�e��uEK*K�y�������	�v�������1�?�Ѩ�v�`�5�b�bmV�7����$F��@�(�C��}Gze��4���$N�4{����Tq�o��/��u�KD�.ٮ�5g�-�p٤��]Bn�;��n~(ޯ��:KS��N>��R5� �!�z�C�%�.A۽�R��ؽĕ���٩D�����2z�ч�
^����Si
4�u�M{7��ob����-�jX^�H��R�DmI�h�><q��h��_�\b��!�;�O�\�k�H����<j&艈���xZu��hmsK`�4����)��܅��(�p_O�k��YC���#�,d�\�R0����3�j��1˪�Z/[+R��#0�U�>����gCs�tu��݃�0����@���ꚥ�F7�x>U�C��/�F"����_&eǦ&	�9%���K�9�YnV�`�+��L��N�r����Ai�k����vn�~	����>����+���Q���c��e;�m[ D�9 N�+�/`;s"+R����K�ʯg����ܠ2˝�
�����׉lN�D~��8&�k��kx��Cd'�.m
�����ld��, r-��{�0�\����B��6�-!S����f@�����YTA\�����o�=����p=Q!�#\Y����-|�y5��\��}}X�]�%v���X������#�_��g3)�{/>33�o�4�o�K�t��Y�!O�J���ea�n.���!n�s}�^I�n[]U��]����L�ffˏ������f�p��M}��vKMN�6�ON
D�V��c@���vC����q�.�ʘ����jt���R��ހ����jI�3!��Na#�ėh��U��NU��~qO������27�k�1��9:x���K�@^C���f�Z�*h=t�Y=�NZ����ր#Q�L��^�X��[&?� {�:��^[v\�"{�P�*$2>Y�!���@f�[�r[ٙ9���f�m�V 07==��pt��ҵ�G��57��ɝ<�m�S*�n2��a��\������"_���=r�Y���\W��i�	�7�"<��_n�w��h)�Z&$��T�,>�V_���Â����6�	�����+�C�k�N�Qn0�
<���W�	u�`ݵU�����V(���1��w�9��ƿ祾��^��z�FH��>��J�:h�S��j2@��*�)�AA�w-��5m2���C�N.�3���cR�ǡ�W�����Q��<Ù���A�����.�Y�����@f�eh�]�;�b��(>Sq�A*O+�G�_,oe�^Fi����g8?;�!�^
͒�c�GY�q��i-'-�ce:��AgH��K��-�aܱ��$z���CY�F�C�OX4�u������tϸ�kZ^���Xq���1�4�#+L�VZ/���-�B�����[�\[Y�� )�ż1c{�ϭ��.����G Z�g@2�7�.��N��@mn:S�z]=� ���i<RG����CoE��,-3���3Lj��[l;BM��G�v��`ԼX������͐���>����]+�w�!���Ʒ=>��?O#.���Z\���$����N�y�Q�NDZ�w��Ŭ�9V����ufA��X��8�)S1yF����m��c���e#��ӵpI��C��9<�r��I�^�z���	���R��~0?I!\�=��)R-Azښ��x�Y����b�_}�ӸC~��β��ކCI��x��.iUm��T��p��iu��a�rlR��ɵ?ڰ�oA�4�""��nMÆ����b�őW��K�������s;fΖ7-*�!�۴��X�1M�J��_J3�a������;��cB���/���e�?`�獤��l�޸��@^�<�h�/�s8�bvM RԷW%�ɒ��z8͘��Y��^�}r7��S0B�����`n����������Q�zl� �6���lӾ.��u������D�ݵS(���O]�٩��:�g�r~E{����I�f�h*�:��J�Ȏd7�#x�?�׸�0�Ͳ~s0�x��"����XF��C��I]��OZz�-U9�?�R������X��i9\�B?W&�>Zz��#���tA����&�@ik��Q)(�j/_J,XJQf����*!_�s|���vٷr��~v��K/�Γ�/6�y�]��+,�[�1/tt�==�!ԨzLh!@�)����l�.'��h�'�%��`�:މSTSi���rȃ(	�A�~RO�}�b��7�<��~��w��¾@_i�b+��X�i��.a�5��)��Ւ��B��]�fk�@�^$h���#iR��2��y�j��c���H�-ԳZ� �� �6����}��
�m3j���Yq<"�.��>�$6F<"l���h����\���j�' Yr��|�+1*�3m��/�Pa�?�C";�ڗ*�\G��-��HF�\��R�Y�G��Q���D�VǶ��|7�D���9�f�wf��x�{YN;/H�x�fk�(a��ӓ�ӆ�QKh'���o�5��m}<�`�_-�r M���3k����y���3?]`�
J���]8w�.XCυ�Z�Q56A �r-T�f�u�X흐i�|D(U	�՝�sԧ�=�PV��ej9
�E��+���4�dp}������_�@�\w�Tٿp�y�u��~ƙ��JV��_�G�Cu$Q�r��fݓ���oG-3|3�_F���e�/Oӛ>���$�n�ÏRZѧe��� �:&���e=�ČpZpV��+��;��C������軪�,L�r�{e�B`h9z !��·�k@憸��ݖ��w��y�{�W4��y�ƕ�	�%C�4�_|l�w�{,-Q7����0�ғ>J�n�}�$�P�{؁�����8U�0e6}�� p\�_�ɥ��[�TSy�14l�j��8rP��W�T��SC��j�mJ�ǆ���Z"��R��_w�3
���s÷�a�S�\�a�'���F$=\8�v�u�SϽ*�C��[ߜUH�,�b������L
`��?WdF�#�op�F�j�e�V����)�&4u;D�WH�t	HL�qRF�2Ы�����|�!zP���_c:M��[a�S��B��Fo���0[֥l����ǜ$9��[�r��yf��o���f�x���$���':*f�v+xh���@�=�1�x6�U'�	���Cʢ�d*��f�R���f�˩_o^�Bվc:�7E	�J�|i�ݕ3����M�6Q;��Ш;�28����W��p��$<I�(x��edk~�Le��Ku���S|/5d_)��2�	��GB?@���t�|Vk�x� �_��b�p�.%#8�L���Jī�*JӼ;�|�m�!�,�05�Η�Հ?E��8w�� ���[�Y(��s�9���0�1h�����ă�_4�j�ԝd>�����#��9�O�'hWK�r��h�.2G)��VJMq`J3�����/O�X�lb�|G��e���CU���G�5晊��E�'����=�V�Ѥm��4g��D�|�@N������k�7�m��oE���>o0N�O4�GK�+��
����O�pu҄��9���-u�{��!L&�MLr�PS"ڸ����ϖ%����#�Ui�Ӵ�ETr��v�� tn���3,�h�_?f�0�C�irt'�q)$���J~L6q��h]ԅ,��(��R7��D�����A���s:Z6^{f̤���5����zo���Ѩ�\B!бӾ3I�mLL~=c�F�e5�#�E&��}����#�ǟ�g-yTH��F|��8M�H��"P�X"Q����5� 0L��ӕSm�;̏�w����,P��tӄ�Evg1�{+!=0�\�ݭ���#��5W���8m�֌����k��V�Y�0�z���>���|�K��t5�]���F��ɸ�[�ɦP����S�*��X���˥�oy�C�L7ad����X��ܰ���$���\�~LsŪOа����+�@|���0���#n|U����M�(7�'�<1z[��:[���{ 0�=×"�V���5�e�4�����ɻ�4y"�V���Q����׫mr�'0�6p�@�P�DS�B9�"�s�E��1����|[�O��?��(���<F����p��,�5E���2���m)�~�f��l6�z}����N�v�@��ނ��G�)��B�J�`����jQ�}L��4A�rQ=N!��&�\A]��{�jӦcԜ��1{�3kg����#���L�Ãz�j�S3��uA�拄dR-{�!������a��઻�����<�%l��GI����+�^��p���%x�' V��G��+Y/��|���m�7�;���q�R�8s�FiBM90赜BQ�Q�L�i�r7�rZ6:�`E�m'{|Ih?�Ë��f�,��h�A��Nlz���x�C���]��"�@t�]����]��q�#�j�*�� ����rfV�I��'M�XIw����/,!���x�I�ʬ� b����1��(O�O�nJ[�90sc8���P�׭1�Px���1J�m�?�0�[�FD#b?@��H��ʨ��]`ǟ\`�{M�������L��1B0ie���/�c��Hu~_?M����w�M�2/N����(�Ď"f�='�Xc��M��k"�ʹ��+Á�+I��ˑ��M�����lFZ�����7�]q��CG⃎�ۣ�3�����}�kԍp�%�zB�0�O��P*�`�gW�¶��HV�x�jT�X�E�Y�iҘ�� �����b��� ��^�G�/�����tr�����J�f�g�����f�wA�ٗ[�JO�my���
�Hyq>y#��Տ��,�W��bB/��������l!/$q��A�'�k-��D�sz�Qg��6d�Cj�"�����a����'�KJC���8�ȴ;$����o�YwVT2�mlJ����2�Ԇ�I=˿�|��iz�^$=B2����ED�GOCT>�p1`��3h���v��/�\~�� � !T��F�!�k�d�	�����ə�W�.?z��#��ڜ̊��F�G��_��� +��'g^jB~�"���&���ot8!FC�H}�E�%�tբ���`��Xc:1��� j)ɂo���
�:�jo��� *g�M�<�p�4n���M0����g4Gv5�r���b�x�)uE��2�ي��q�	H�S{R�l-����d�JU�)}���R�	��H)DeO�HEAV��[�ҧ裦xY3��7�A���$�T.��.Q3+������Ns����p�H>�����
�lI~$o��1��Ԣ�y�M"�IFس*�@ׂ�"�2�+�*�� �m��M�y��I)�������.,4����3kr�PMoU� ��Ez���G��aO:��X�'��$P���A������k�S�rdD�Yc,I1
2����@���xz��B�����΅~F��
I�W�f+c���%�a8L|F�w<��%�;�e�Ы��_(�x�0%����ǒ�1���h�(R�1��$G�($�)!L
����aHEI���ˌig����ݼ	��KB�b��1Y\��	�AV����ON�'6���0�#8�h�Kn�"���&:�o�>=V����i2�J�o�	۵����9CB�>#]0�,:0��u	t����S�1S��U�A����J<kI�Tg�jJ	y���y�!m�96≡%�!U����Ć�|fx�(H�.�z�DB�����ʻO
��J��B-e+�ޣ���[mo�'�\� �rO�&����we�=�As�W��ca�~h����$�􇉪1�U�^s��@E���G]ʙ\�w`%�9֐\Ve�l8@��} �}3�H��I��afPc(`c�3����2$ �>#mH�)8��HR{�R!���R	.�������H"<�>$�{��������ʧ��~D�=�[jTvp-��b@-�C��5�P5�s�Z �"�a�������G׊����C��������	���th��l�M��rf���z����FK* ��B�e<D�G�w�*���>���4��Z�4jR��OM*s�B����U"��� �*����}a��ը�q��R��z�o؆��+�J����G�����> �wZ!��N�x<�xD�O�ـ[�L������T�,���[Hd��-bF�I��t�X*9PX�+�(�T���z!'j�,��� 8[�BQ�ǣ(קK�+Ө����L��u'{%���t�z�7��d�H('���@����7�/<zNhPן`<�e� ��e� W3���gѡ�	�GR, 
��Go��{M��\�6RZ�/��6[�B2*���e!�5�C���l?:����Dra�kT��GuY>�Vm�������_���d5�w�"Q@i"���U��z"
 �KY�kY`�2t����������|�JS���u���g��=Ff�_$YA*&���7v�oG��H�0�D፾��P�qI%����?��.)��H�m�uXQ
3��d��S0������8?*l�u RЬ�.��>O�(�������;���ӝ�FH+�M�Uhgᯉ�s꾧�DO�$�}��7�RN)ّ+$�O��0���D���! j�䀵��s�����G@ �FI���f������H"��4ɿ4�|�j���Q!�v���4��p�6K�+D '������bBp������8)%;e`x�j��Yv@$�I��B��d�y��Q�L�+�L���Ϭ����c�!2���D�RB}�y!��
����}8���1����R����#y�*�N@��	�,l)8��"'uA��T9����@&�����(�'��TYc�� `�n��L��I#�X�_�:�C��j��7��J	�o��d"��L�{��(�e�Lmn�%Lr�~�<*�������Hu�hk |&)`����Ȓv�}�!�>���)� Czʐ�?�ㆎ�������,�<�D���!�
�X��i���N���~3�8��,a�%��*Y�j,*BB��F�Ci�O��0��������-�2{���*&�����OD8E6a���]���}��ޜ)���������_/�6����g����;��_�b�����sqr�Z �d�t�m�0	�#'C巳EM�����s��M��	��IC'����s U��~ُ���	]�����#�zA���	��ی�z9�m�ʪI�/���ݼj���`m�2�K�"����_$�Ws�Y��M��������lI��xL�S�~q�z�_?��S��$��ERȘ!ύ-2�Ʒ���>J�w)%���;���L��*�׭�*�y�ڇT++�݀��rGq$	�E����#=�P��8�z�CZ;ȉ�1(oE�(��3��>R��4�f���3`s&@�?���!����l-��m���]�`.)�	G˯����9��M��!M�#w�]�<_�_"���&:&V���g���	Qg�|� ~ �B�Z����\�?�-�P*A�¸��A��#�G��Wd�	��o������ͪ�ܱ�)R�4�k�%퓔��l�d�/8��&��ܢ��eƱwF�����X­P��K�p�J%6�аZ��?d4��=�N�E��U����4\eX]�����) )}i.��%��)������Vi�K��t
����|?��3眵�^{�À�/�E /�`]�� ?z��=�;(Ӟ//�^Af��m�6�>aV�<٨e���	ĔoTVM��H��z�VДHR
��{����r���t�>~��:�F�@��b̓�K��y0�u�G���,;BF�b?��Yb#�%���5����lK��G�4Jwp�/r�.2���Oax����4�	0�I[�6>��Q�g�wC��j���UC�s���<�qe7;�x&O��|��A�b{�ĺ�$_wFi�^N�3Oipm:N{|�B�US�ٱ2�Ե���e~����c���q�p)�^�~c��$�����V�h,�ǟ�I�I>��)���a<��|���&��h�gj[i0CV6n��ga�Q��xC��U�1z��R�i�nP��C�2: r߾�6���zd��
���G�"��J�@?9t&,b�~�`�j��{��T��2g�8|��c�){�r�([T��Ϗ\��]?�[�d��}�)K��o��F%2��q<I�2�n�������X�z9O��+[H��!���|6�e��Q�Z�t�;VSşE��i�	�7�W��>J~�tY��fG<T|}F<�pa~��pr&[��J�(��ޘ���(�%���J�@}X�#tf[/��,5��������]fR�э��D=��Mf��P\��2��a_A`��Gz�-���+�y��ԿC	z	S'd�J��'�<3���Q�E�-��أ�n�8����t��ABP�k̲�h�Y���y�`�f�X�kOe]�l	�1��-B(V�VMOq�Q�҄���%)\���5m�%�:���Hy��+`ߛ�=]Ϳ�)�*�H�l_�l~b-7�[ѹyl��w��'BUI �}6�?���DV�$�_������o�\]��"�������"D��� �2��M�s-�9�m�,���v������n�U?vV���G�	l��x\XS�&qu�r�^	�\K�iÕ�Nx��dPP]����f��'&���(���We���+�F�N�܋!ų,�[Gm�w�����F:������^耵���k�NhbY���0$�V�~ک�K��WQ����!2j�EAU.w���z ��.d��"iO|�<�����p�5Cx�p�&���R���n5y�ʬ�������}�����>�Vv�M���t�$Kꎨ˂J���6��z�m'��'P��[a�]�(?��n��,/��0+>�7	X��{O<�rʪ�2�T��il����m*��`f�EA�%s�̷)�x�2�������� �B:��O�j�@QG�>SǱVZ�yv��ͩ�)����5]��o�_"�Ff���Ѝ�R��
��#j�*����H�*!���o)ݮ��s�.h&@$g�s�ʠ������yy���Wx�S�(1���w����G�7�����r��(��s��;���Ϳ�LND�d��cB+��gV3T6@����HܼV���|���l1�o����z����_��:���Qfp{�^�E7�
���v�����BY	��݋�����q	y�}��&cd����8)�麊�#t/+�^�k��n6cǳ��F�3o-����ӌI
5g�L��4��	
����!(� g[��1�&۟̒�Y�����Л�&ei#�������7[���k�QV`�4�Ϫ�|h7
j�������:��jCr�K&~T� ��*7�D|���o��#>�.%0�6��ߔ��L�{U�Ԁ9(M��|�z6�� �{��*�|�)��I�"�<ƊLIN�X��Wo2��@)��\|�`4��Z�fX��������� �ʔ��.d�����߄��� ���Z�o�RQ�A��D����y��U��xѣ��C60N�?C3,1_O�a<�s����!��	:��JT�!f����\A�&t}q�Ek*�=��]��`<�A}�G���־�YuP�r�˺����w�*{�B��0����c��ԕ�[d�tU2s�T���~�2K��ĺ�� ?	27VXw������#p*d2���2�<���1a���+�������=���y�2S�;�1l�	k��J$�~YA�A�E�C@z��u7)ɭ1ǉ�9@3�g�ve+���A���c�C�z�)-Ocvo��t5(��Q�f*]�O����;:��4���%��'��Z?OT�g��$�X���W�=|����-�/cq�F�W>:g��
����e�vi��Z��bP^\&����P���y$�fq��{~�s�[.�&$M����a�4qֿs��+�3Q�(u�B��!t��d�L�Z��x[/p��drT��ʙ������f����ҧ��9j�>�?Q�Bqyʻ�v�O�x0��ޒ�p�	�*d'@rxŢCd�uᱧu���3��Cd~��'Gͤ'�W��t��C?��D	�-7|�j�6t��"�3��|�*e&�����l'������a�-�k��`~s�c�E���_�(��L�ACSce��]c|�(����TǇq�lQ�n���V�����q�>#8\:������fG��`��$k�Zl3xS�:l���tˎ�~[��۷g�Aŋ��8�9'�߼^[C=��7�b%�� 4lD�TbO�g'k��<⑏��(ss1��.pB!��J���I4�s�-�+��@�e��2�h���	(�~v��G�:��}V��}��j'U�,�Z�<#b��\�S"�Iu7dz�*��V�'�A����0p���������+�W4#�zX�8��ۿ�{	9�6M;�&?/���zEh�0�����<?{�;C�q�����ϛ�h����|&�d�܃��r8��y��o�ˀw�����n<����0��s6@G35r�#"�m�u�ǭ��G��\��cp���}�zS��YW$��-e�Z/�h����	������8S�n�O1m���gV�b�zj��Oⷽ�#��7��� �W�UQ�-���ְ��#T^Nl+���[a}�/�x2�l����J�gE�<�ͿK�G�=N�7g#�xM݄1d�����m9k�ZԴ��t3˿@j˃��R>:L���c=�K��M�`4�0�Pu��ew���(:6F_i��b@ �t�4I�4��,�N?m.
.J��Zym�ޒ��M�s�%���2UA9?�ݷ=����~�G�o�5v�#����q�hL!a�H�`����[w\��ǝ��w߰�����ϟ��]�t��w��u|�����H8�j�=,mz,�j]i��@/����d��>,��=�����Z|Zt�G=��`��<��zĀg��Fg�v �
݄o�o���gg;�Ҵ�������ߖ US�ԃ��*����1��w��'3��V���7~�1�S�>g˻/�F�{n<L) ��d�6'��>?l����x���O̯^f�N_dm���GY�D{@�/�?���K|l//�6K��nK�L3�M6��nB|!��]$�6��ȶky]N��B���A�,��!˿����r0h�_��@r{^j!l<���e��k�� � ������Δ�˃�Jɤ�6��租_m���R��!��ڪ�Vq\�"��r���4�#����u�E��:
9�h'���ӫS��C��Ήo߀�񜽏ϗO;��H8�\G�N�6�g�m�|���7S,=�J9�h2L�q�"Ү۷b�a�l���6K��w#�8�k�q�<�����,���9��f��8�jU;ڷ��J4��~���\���D�'0u{L���EBZ>;�g����½$Ur��^eC�Te��,�i��~�8�w��մ6�n}�e�t ��󐪟�a`��_;���eV�h����j�Tg���\���Y8L��׺�x��_#JS]�!���(�R�W#�X�PC�]7���) �����B�wN���/+��T?<WU�\���v�������w�]D�9٬5p��FcQ"�-�\��@�?���_D���C�Q�}l|������u��:I+�q�{x�-n}%{�x�iZ)P�����U�S�
6�q��p��N\����l���y����ui�)���W�ůݯ�Gr�@�fy�8��SG?��� `��v�+,,��Z;�_GY��e�8ҟv�^9��ڧ#��� ���W��\���g��]<�^�����
�\Z��g���ܶ6H5bKrR'���[h��c6 "�S���Տ���ӎ��#M�_����h�W�}�i|p�Ii�(����Zo�{Q����з�)�Y#R��,2K���~���w#����߂��e�R;}�P����)k7�G�69���{��ߏ��>�e��Z]d:�Ҭ)h���ϒ��ݯ�[���4/C,`c=�>����<~�\%D	��.wD�Kv�wv�-~>E�q׆���|�Z}�0Xr��(ٚWX�"� WلK�ٛA�j�:^�n5��Yz�\���vs��%�Ш��pѧ5U)�ں���L�l�t���)��1�e=�Ì��P�$��%[���և��U=g5��<�4H���~_����ٸf���ꉇM7����!v6��W�+��(I���<R����S�E4"6����оǛ�5b}�J:B���>�Ds�{����#J
���f���a�A�1�<�e�
ѹ���ev�N�� "g�Z�UTx;��@����~�C{�[�v����}���xJ���\;[����H���e�"M�[�;��U�sY�����K	�|��pj��]�킎z����`�T���i�=��G�ے<;�����sقF�V 2F�#�4����_��t�d�ȸ�U5�G��{��>�y�j�MsUgy���k�|����c$9f�V��X����]�]
�˚����J�(�m���s�T�����.��7����z����9����X�#���=�|�'���
�o����f]�������4�<_Z�D��ܢ�{����S�H���yިe= ��<���q!�|��YO���S�M���GU,^�r���b`��m-fN��"��w%{n�w��2����ܳ��z3��";��.]�AVk��/g|R�]���ZL��k��������- �1����5j�3F�T\�Co�N�=S�����E�)�V�?�/�a�t,u�*�+�E���BS�'��I]��/W�JH0G��Q[��q]�փi�7��@s�Zk~i���Vo7��H�8�T��ly���n��]հA���eGn��J�4�ɇƽ�Y�4��\ �J!'�(;�j��+op�Dر�P�d܏<{)x�}��ܺZ�>����p����4}O�Fk��]�p�|�r�{ڳ���~g/!�t�P����Q����;�ՁSQ�.o9�kLNQ������΋R��X�����UKJ�tE�y�����N��_�Uh��8��/X��<�sz��r��k�gY���9rq�b�y��!J�8��Y��;����he��p&*O���X�F
�\M`�r�\�B�9����?#f�?.ܮ�n[y�Jv}��l+>�t�*���ô��1�4N���Ut�d�1�mk�����`i���f=���"�=�v�*�*�cm�8��N�[*Û���=Iߧ���,�y�Ш" c�t�opW�jg9�ݪ��9���%��(�K��ilG��n�]���_z���y��Jh߉K�"������:~.��v�oB���Y�@5�w���Eq=^��w8���?7d���J�z% _�N�C�e��.<zh_P��|*Ҙj�oV��NZb��s�/���t�V������=x�(A�vg���ਯE�Nw�*`��~����u �pOTpAIj>�{����J�~�V����'H��!K����6��}r����VX��������`�4z�:�p������z��;���{������>]��CaJ���*8!��Q�Ke u.k(N���VJ��K��b3+�✛�ގ�BI�Ikzؿ��yF�^�%�r���xO��[=���U炒�΃��+�,ed8'�QȰj����H����c��kO�9:S���B`�RLs���A�e��z�d:/��Q�e{�v�态c� #ɮO.c<�$��wa�C]�X9�j��N8���Al�*�>,I�7#��:�4��[��M��I�N�������+�Tz����h�^}�9�hsH�KB��O����An�OB�nWcT�-���a�ȵ�$��o����.a�Y��F��_7�{e���T.D��X�z;wq���֍���5����{�<O\4 7�T���W�P͓3�F��g�מ� J�/�w�ש�SҬfAR�Ժ���\t9�0��;ݓ8$�*�!�! X���sd�c���IϞ\`�C��Aza��4������|WV��ɿ�x!���U��A�t1�)O��ƻo<���N�o���`���Ds�n�q������hz���������M�V �͊�fkS�
�O2���F�P��J�9]�9�F�,]����-a4.!�E[�k�4��H��L��T��0��V�锤����诫Z]���kuXn}���h���@��nv�
	�Ln�<��k�xPf�^�k	w���s~�Z�ak�C	�V����g:��ulihQ�-�<��|��}��94
�C���}~�꽁���Đ��a�����Ć��c���F�_V'�Xyj�c07�p�T$L���Ұ�!��(��y\���>{*z���J�v_:5��z甇p��v�@GG|���k������E��8ӈ��!f��Q���u���[�ّ��˶ G��E�+U]��ē���N�L=�Oеc:���a��:�e�o�

���@>W"5�N�4������lz1s��T�!"�v�0r�V&є��5�3��i�"��	�!AA�+_�dq����5w�% �tEV�����?�F��&�]J*�9J��)6<��u��S�
p��
rK�o��{��k�`dwJGÀ�|�q�;S��.�ג,��ٵ	{ϣɣn&~�f
��P�FR������D�%�t�~�wf</?��%|��E��j:��r�v�Cs��n�a�Z��e�;�+��)প�#^l��IJ{~1|rw�u������ֶ��K�xk�/.�V����̲Ij��d�j�	DA�.l��ɶ�ϊ8u��� ����Vڮ�|�0|��}�m���-=-�fK��'s[��}k2i!!^�S>�����U��-ei2v���<L��\s�y��za�'- ��]��Z /0JQ���G���\>"�����'uK���ʹ��ks�zqPI��c�]��TG~:����oi���[��ZO���T(q��#7��&g�a��v������G�l0�ǯMw��^~���Ai$@���ց��E ��'�L�g�o��n=g�=����_��aL���#��ΌC"`����e��g��cO�]����t.��ώ�N�Zx���&���o7d``ӭ�O�,���>9�a����;˗ˤ��Mw&�vm���
�cb���\�4|-���ޑ��Gm=�z�:���Nh�/v���Y��y^�<-�]��j�������Kn[�X�$�z�GpBZWP�Y,��),wb�b����ϣ�׹��~x��U�#db��ϫb�<�4�zzZ^�`���m���W��J��(CY˂
�����*��o��~?����d^��^j���5u�j]��ֽo"Y	v�z6}���_Ŀ�*�Ēgm^�Iֶܞ-r��?�t*"Q�Kp���I��j�C�VŬwi���'����H�q5�%~zX��F��/��s�S��T����S���Y�s�p*5�1��%{���\z������O�����;%�+�K���LG��Ib/%A��^=�;�U�_ǾU%;(���;>~�\k��4*�� ̾��a�u�[����a�����cW����|�񤏋��U�A�h�g��/&Nd���zN�usO��pV�v��9�|A�%����u���C>��v�_Dǚ���4M7��=��f�[� &�t����A_+��MlVeϣȳˈ{��>&�v(AQ��1������MW���l���Jg��#Fg�qpݫ��)��g���+NͿ�,���������Z�FkՓ�{r=X27�'9&OY����kA�Z�"��̻�N϶��.M�U\}�o����.�K�HA��˯�8N�}�p�[=%CWĽ��&�)�'q����+ݖܫN�c׹�&�����l|%�����2�ۗI�ҭ��v7�5<l��g����4�ܣ�|�r���8�Lz��vX"^c� W��&:�;<�hqO�㐈k����/�G����R�(��;����,������b�n��a2�d��j�̂��T5Ƶ��
>+ ����E�5�z���xN�o�����n܀*�@�C؄GW�cY#��X�����=S��u0��s)�C?~d-2�;�7�]�u �(�m��Q�Tzͅ4�T�e"�*�˕	�AO}�2r�i��3�ѕ�'w����ǅ��3,
@���hqc�0IL>7ߍ��=e��6����w;��p����`A^�2�;6΅�v�sߥZ��H،�囁��^��Q��4'�"Ɵ���,������1�xM��[9=.�"`�r�v�z��_O���s��ZOK21�B��g��y]m��#M�˼k/��YMAEA���%�k:�\�^X!��x�C��\i����� ��m�fƊ�\A��\��)�'��=�%^��j�����9�g�	�Տ<�+ª��6K�a�N�z8��是�i蘽eh��M�%u�z'��Q2\�p逳jW\�����y��/�I�:��u��ւ.��t�7P�=nv]��g�[��>r��C��[<������}넄l�8[��d�+-'w�0Iu�F�q���Qe;�jZ����gf�������輶3,2�NY��*�j���L���#xy����s[9(JH�Rj�\������&��H�|�z���I��,�{�L���W�����6������*���mN�p�X�+|.���ug�K�:	>�7݁�+=DK||���˔�Jle�n��'M��m�g�����6�z�Q����12��9�uD�r�O2��Jn�L��Os
�U�Lfi.�T�_�L��r	��k|t!��v�uT�,���<�Bo�0^���Cr8�s[�S��X�2�tE�L!D�WA$��9�V��~�#X:8�6�k,�C���j�b�/����~�@z�� �y!�5B�2�����!�5[��=��|�6,@J�v��[oށ�W��� AS���;��ŔuRO����o�C�,��Y�N`{Im����:���wǭ�[�|L�S¯H1T�'�eK�O=L������z/#���z��!-�짗��ܶ���%�M����fq.G^�ց��D�y����ɕ�}-��*���D���a�QV![@C^�e��Tk�N.�\��/!�$T����їF���g�v�륑<5�����[.:�C�\�˙���;1���w��!�%��3���jS-�Z�xѕ�	��Ϥ�4��;g���gU��IH�cq��y��طxѨ��F��{C��@p�K�n���2�w�Q #���d�г�Qa�S��PE<�9�&G��2�����ݪ݋��R
c�k�I��JRV�u.t����!�/v�v����yq3o��?�; �\"�7�N䲬����啖Ä��pXQ��a��\]�� ��IΓ|�l�߅N�O�I�fs�"3	�*��|3ܷ�>+[�����p��/�9�&f4�[)�3�}9W�4�!!G����n�>��a^�Zr�W��G��5_� 6Y����GExy�$���^�,'��n�����J >�{O�!ω��Sf�Kְ�.d|�	�P�.�I������.�p��m��A��5��H�FF5,��=,��� \�{��O�B
x�..��#�Aa����:�̥vG(�{d.�VǄ��#lZ3l���z������N��i8p�tPb�l�b�0~6�����R����m�������GrQl鲿3?����2�r�O�`����E�l	
�Y��m���.�8��ˏI�8��n4�ދ��������j���n'gn�z��rP ���U�S�� }�4T�U*�ߦs�[���p��|(�GH��hh$�rM�k��qS�7�����d�sr-��Q��~Z�s�����ǹA�(���(1�HT��@o�w���Gyjb2�X �\�[/���H�29l��S�/��5E������}��g�<���èfܼ�(��6(�V�� k z����l\��	qp�� ie��f��D4~3!�Dz(�E^,=4&"w�c�$�	�s���p׼'��k���3�y�4���2] ���g���k޸LAf=�c���� cߢ�G�	�ͷЮ!�����}�������ͳ��l��H4�\5�W���|��PT�CTS��86�Ӗ-FB�$ ��H��x���=ZvwKJ����
31�	���{�B�g�d�������xM��iѹ�1���ۗ��=὘����-3��_cH�
W�@���T�Lӿ�^�
�K���x�"�Rr0��!�k���ls��Hy��B&��w �6��԰E�?M$����j�Zp_}�!}H���֩�&k��^:C��%y�Ux$�Em��%���>(�����6{Z���4��!)����{����G�$c�+�xgߪ����~���
��&փ{���$C#1�	�T����(J���?�q<�S�o�����/���sL(��:Np�a���gh��!���IZ�yE<�$<&� �#�K#Ko>��(%���Y)\�䤤�B��A���n�4z�-�<���8"]DQP�K���+(�c�ݘ��,%�1]�+v���.7v���CRT�bm��!�ܚq�1m�z�e�0G����7G.Svab֑	���?A��_jѺ���H|a�kkQ|�[k��V*�/���m2&���+j7q�!O�K;�ƅ)i��a��ޣV���`�Ti>�l��8V�7f���fz�v@�E��dr�S�N�Ub�M$�04*�߰LXJۣ���95,&>^�������e�SH)FL),�y�
|E#`|��F��U�_�M��&�5��f��Ptx �	g,3M�r� ��=�"&In�'8��kA�"1 �su�cb&���m��R�Ӫj����W�f���I�[�����m�17.�R�CBe���Nڂ�p�g���f�x=����`D��	6Km�O_T/h;ge"�4[�k��b�7M���	�:�/|��}eӴG���`�D<�N�2���$P��ު���YlG�c����Z 7�bM(�"��Y�:n%i�l�/�='�u
�W��I�&E�"M����E�?����]�b)�^��д�P�����/2FdJȜ���ʜ��ؼ�։��a;�u>PWT��������wW̨�&&�Kέp���~�*[Y�u@{3J �h�rL��x�����$��σ%����:.�0Y: ���5�Bjr���9-!���0��ʵ -x���}V\ �@q	�I�u�P@����YZ�(	�Z�Q�x�¡��?���Т�p�#�m#+}f`O0�0�P>��S5�)�@�$��xs�B���߸�v���w|��٤���6��ԅ�Ya�����a�/(s��O�=o�K�ш�5�
㧘�<��ኼ*&�
��r�d�(,<�f;�HsE�ӳ���s���cb�.=�*��  +��QWZ
��zo�#��L���p^LyH�������XԌѲ�b�޸|M�cLynn�#�
Eh�Db7��n>�VG�X�Y���_�;:|Ӂ��oK��r5���q�k��ߔ2Y�x�`��d�e�8��������B�V�r޴�C��!!�֔�m
@��n���!ȿ.��\LS�DU���ig޽G��M�pa:3��|�T	)|�E0V6�"�;�b��֒C	��Y�5%,�3�#�����l�n���(�+�~ϯG��]�00���ǆ�ge��ZAP�pL�{P&A��I�ZJ�8!�(��@�6�� u�;5�3�e�=�S?�-��iQ_����zO;�ğ��{rd�!�4��$9s���@OU۹�!�T�&�R�d���nX�H�K�x��?�-�U�Mc}��k0���H�p���C�o?��s���k� �sx�P�*�Q[ړ��W�"������X��[~/�Axg�V��S�&5��������a�_V�k�A]x�S���W]��d�MT���0[�~ ��w�j�zaĤ�r�zd� �-0Q��I\x/�T��cP��G�����Wt-�}:!c#�<8�jH肾j'tD~���4`���v�/�r:u��Aɼ�?�MLM�I��z�1�ϳ�q"Ǯ<g������S<q����/<�5`�2�<.� _�>SHN�ziǻ�������4�u  	�p��X�G���s��t���7[�G�$��Ɨ'�o�
�Hn�L�H�^B�P�}���U�2�4%��̟��cm�EoUN��Eט��2~G��SH.���=��tt�O�S�>�2�й!E�nb9zQq��u�>D7|l�B\�<pf��<C��ˎ4�5�,?�w�Q��[8��o�څ�p�)FX�hB���_��?
⋿bGX+2��� uM���]����J�)c�����W�'����/��[lHj��p��~�4<0��h��`3C:a�9:J����Q�`zQ�$|ŀ�H�H�"��!k����pa$^�X�:�Ht1�`9'�	K��њ�� �� �ų�@1���_��sW�<�{])�Pq�"�8፼>��i��3�  �8�z�`�<�f���L>GCL�Ɲ���{d����J�VM�z% "�@�' ��p��Կ����K����;:�$��fM��ϩ���.���Ԯ�%v]k,$�t�t���̉h��S@3��-�s)R[Ro�չj-*�c<�Mj������T�>�at�c���c�`7�5��rO��@��ó���}�����宲&FQ������7��#6��骬0��x�IBE��^mq�	>	�`�Lե�y�d
G���M����I_�����7�9�+� f�"� fC\��Y���%����k�$�%	��2X��65�h!,#p��; ��.6�LL·H��1�G��qE���ޜᯤ$F��s���=�����
~�Z_�����ԭM��H��4|��b�5m̐fq��s��椳����:�@�����[�W��*ygý9V�M�����EOT���~T�^�'g8��	���O���KMK�����I�7������!2K赆����b� p��{�Ь!��f`��9xO�q�j�uP&Ԑ�,{Z���pZ��x����l}�5���
�U\�� ����%�����9=���ᒺ��
�0L�ŢUZ���Q	� ��<�:���6-*�l�B�=ɖ!� ���N��)W_���	�|���yn��IU��ʺV.R�4t��e5�K��ЛG �0�7t{���I����),������U �����]rE�lh���o��U�ȃ�ԍ��/�a��GHtA j�	���-�����w���*6��5I^A����2�G���S��2D?	(�%��H߹uH�SJҁ�Ş���
:4�v
��P��2J9ʠŮ��uQ��*<�e�@7s�~�6y�� b����6�V*���	a��ZHrKny��)y��[�̝�W���A��F�xE��kZ�&q'�~��+2��D֜a���=��P��܇��۽��I�6�O���_�d��4 ���u�N��1���q�d��;��F��Lp� i��5�w��{*�z#��۫����
�Ϝ;o�u��%VN~�cZuNq#ط&�;-
j$����F�;��9 �������z`� �?7g�Èq�	�ɣ��W�!lb���&n�KJN�{Ģ�������5mo������=]� =(���3�A<S��;ɌX�SxA�����B�T8=}@0S�쯊(����u*`8��\����P1<��V�RV�{�ߧ���Tn X�Tn�۞A%̺7ce�~m��Ƿ�w�V���	?3�E�'OoK�1���@1�8�Սo�qR|�Zp)S�Lza��G1��޿�m�fl��~1D�/���$��^o&�+J)&�����S@d$���/�f$���4F7^nn*2�����M| �PLk_�5���J@��z�JHw�����x��ҳ�X��
�*n��~��4��*����L��VA R�����v�*`6�T�{t��<z��K��XJI8�H�
�=l�*|����g�,a�0��u����9>с�|!h4�o9L2⪋���_~^�â�?�m+Ui�&M��V7k!YQ����c��_Dꟃ����~������̈�"���J��D_�n���:�D8�׍h��a��[�ie:���4�H�S��5`���)��(J����}+��So�4�R����x���ɼ�\3*Q�|8zj�]mM��5���s�89�<10f=��`�C��>�j6R_^V\;BR�q�np�	��/�s7Q��p�m����y��\�vr��Yɦ~��G���5Ue���"�1Ko!��I,��"E^B5�VPB��v�يTi��Q�j,�Sr8� ��L\#f��1�^ �]A���B_I�� �
�e���=� cB��i���TI� V6�V��-���ȝ<�	�D�Y^�����*I��:�Kˍ2,�P	
��`�D�
��\�D���m�rg+��w�xa�a��j�蝳�1�S7���ί�bmn���뎘��/�	u ��P�W�&���+�t��߂c.3��R$s勳��2��
Լ*��)������P�;J{�n�y[�dU�9?mVk�q��gv��d�G�U-�x��0���%.����C�w:�.,����=	�N�׻��+�U�ĀrՂ��k��"%8~���1��Fs#>QL���3]9��ۀQ�-���{p;�����`�)�U�p��S谔����ͼ���L��@.,��+^���G�YE����;$����Q��1����,�J�e�E
�G�S�c5)+�iR�"OrZ�?l��p��~"���̂�^��NW�Bי��G �| ����'T�j�;\�|� ����Ͽ?.v����>{�[�G�S�ŏ��7A4o#�U+ߖ�)��m3A&w�i�,dF)J�ʵ(�����8�̸$�(����HIN�$qe�$n���,�[&!6?Rԙ�S�5"&��ףw�*K��>?�}��Of��W-��O�y�������3	'x�.��T��q�8E�QÊx�q.拙Q����ݥ���.��u4���C}T&,\���$��0���K���X��	�� �\����|�kJ4J2G�|8��ƾ'<��A�#�3p���`�ň����c���Ǝ���B�d:P�6��Rżb���_|�����M�p@+<����	.���~+q�4c������%�Tepl����<T�i�3�/1�(�c��$m��1�6�`e�9_|����"� X�0>�׼�yt�$��� F-�*���v���LM(q�f�Q-�k�f/�s�FC��י���P��'ʲ����is�
8�m�=���)��3�F��A�v	�c��$���`̬��:����E��5=��'�=|���֎��"��IS���>t���Ņo<�o�X�,%+X�Pd ������k�*�����T��n��Z��̄�Reӎ"�Ű��Qxx-�1S5M���&A�񾲖�����`���M������?�_����bI/����r ��.��y�*e�A���('+�,�U�gc�< �-�z�{�k���G\��>I���ǜ+r<�]x��+My!�%ur��G]�������Y����ѡ�Q�Zn�5�b�f�R#�N^��P�-���a��Ja��A�d�I�~����/̪��1�Rj�(X���Z��̄1�p�hnN�	�[����[�[$��d��9�̟�5��A�3@0����A��8��50�@�󧙺~��ar��@��c�j��#a`�M�QrS���G��-'H�J�>��5���D'K4h*�L�LC��K��n``��L���|&"�-�G�]��ō�b�(�-�.��3mG�vQ����=�F,H��ސ�Ql����g v�Q�uY��w�hm�#Y<��$���^|U�w��da�Z�RPJ)җn�����E��W��}[E ][��?�.�
wȭ��*0Ldr��H�Զۍ��K+^�!�p��]�X�Y��l�H��w�䐦���(���E]��t���& :�G`���x@�Hk��T)�%'"$j��rt�瘝�ҝ��F�iX�Ŀ� �T	D�\�f�p�?�����Wq��
qFG�G$G����z�[_p[�٢�u	Szk�_-*���bq�ňI�Z@3��~c��5)�@ܞT��&*	ܢ�?mǢ� v:�w��Q�잠-�|����̖1}�t0n.�d��߅��fr�-�0K�A�L�dN����JF���ٟ����2|�l�'����)�h��c�a!��������n��$��+�؆9S�I4徕�z�6r�an����>��(�1��?7�#D$��������Y{}����|ޟ���=>�m�mR����C"����Z(�xJ�^��L7B��[�3�9q64ˋA��H3����w$����Ź�}Pd5@�c��-��W����y����-�y�}W���@;��u���\d����;�CB�g�g8��!g�i�n�nB�n���6�ˡ�������ӏ���������i�򔴑�!� ���Jw�Vm@P�߀f��o��i�!�ȹ�����p�4���ەQ��jz�r�C�5����+ݵ��s�����l*����2fF�����r��ڤ�g4��v���=�x%p�F�)[�Ĥ���χך.��Q}䎘�m#CȺ���Z��X�ƍ���G%����r����"�E��p����!j�Ӕ��9�
E�Q$�0Ed������$.6e�Mh�^��Y��d��IP�ܖJ�N��ї�q�.~�X����z w�-b��:��8�Q�6)�E�7WI�2���;l��4��j����ß�=J)�i]
����Sݘ�\s�����:�-�~�&OD��䗹��I�]������2,p~/t�MX� )��#]�]'A��8QX)��f���m�8%�'���c�]�Sj���������0�PeZL<_�w��Ke�$� -��Y� A�6����`g�<6L��Pcev���d$�e%QJ�Q+��˺����lh��"VPŧ����G��>S2N)/ѱ�"f�3���DFRJ��L����k"�󛹥͂�q�5V���x����쿳�8Tů�P����M��ڌ�̴��,��/+��%jѕ�b`!2����h��'�����Ua��`a���L<$$��_*O������L���P��sTc���� <�K�U,������:�0?� u��HK���`E�?�U�}�_�&��#@4�c�,x�1>$.��g����8�N0ʱŲ�I}����!F��P�.h�/U�s1wS��;���ޭ��9���K�#A�TS�:��R>�Z��5ób��0��H1* �J*$�峗@�7�p@�LA`z~F�I��'�*]�����4{Z�9_~���O�w�B�����p\N�i�ߢё!���4?�YBNqK�M��z�6A?��	T��!�B�{�!���Ypw Й�o��\�<�b���$sX��j�V�x�yItϾVF�5�~��y�)��~2���J$ڨ�""�!̯�W��mkq¡��9���C �ꁧY_c?�;ֿ��^-���)�*��H@
\�j��	l���`d�쇽+��w��X�����%	_�M寋��I6T���Yҽ�ikx���_�/��^)�F�c�n}bpӣKD��	�ϻ���ȡ�U����y'|#H�w�p�% �fv�,/.�^_�l!8پ�U���e)z���q��ƣ�$\�>2mb~���ܩ��L�.w���b�c�O�}���{j������T1K��ި/<72W��w��Q�F�=,�H�`�!Jo_@��.���(�ao�%Xx��tk��Oi�L1���%8�Q�?�YvG��t:��_��}u'-�/���_���R��l��9y��%���.S��-s
�0��a'����������k�pv���F1�M�[|��^H�c�c�OE�U�	���% ��0ʙ#�g�NN�n��7��9�@y,[˩ K�|5&��>�߾�,r����a�>�__x׍5��c�򃎨c)��+Bv��߇���黍hȨ���F+\�}���5�N�ɗ��fF�D��a�d_b�m��lm2�\v��V4�tD��Np��M���E�AmVrYj���Xc!7=�C��5���0�"�V�� {2��'�� �obz����0:-�f�>{���`B2�ծ��6������9�A㮈�N�# ����
��N�ʍ<~�G����q�P��Pyjx�*)L6�moA�e|�e~�fGMb�U�K#s��cm�r-��t��@F�?ߖ��Z.��� -ܞU���M�=�s��-\��}�4)�|\^�j�|`�6ѧ�������5R�k����_i�)�*đ�����-��a"�b��zS�J���n�(o�3W�̉pAq���@�b����-�F!8�{�0�	�m������a�F4�'%�3269 0D�_�HP�,<e�GY�RdP��lS�ˀ*IZ��d�pH%]���Q5�����S0;Ҵs��U���U���xF���.䍔��g�;O��Რ�0˦���qmm5f��\����J�\1�e�L�$�`���wu�J���?{�Y�^�'�#���6z(��ojN��k8�.7>��Hv+(7��
�graSק[�3V9�����0r����6d�����8?!���9�Q�o����x��A�!�"�ݷUe�M�/_��Z����3��hc�̾����ti���M6���6��Kȧ��n�a}�]�G�2i�fH�:��3�צ~.�F���j^�뭟[V���/��
�aN�0�%��2�vl�n��#�Cֶo5�O�.�<� ���Gb�.nA�����]i��ƚH
s��Z�0n'�e�A�
�t���IN���z>75�uU���H�5�I�K.g6@��"����٪W�n�����ߎ<��ᆌ���[PW}���4:��L����n�
�4�?���f�/�IXTw���&Z�2LN�V�v����#�6����bUkPZ�H�l��s�)xɣn��sO"��J'�l�i\���ٌO���������E��ŷ��"%a(N�#/�GY!�l�.)��|�7b�����=î3��P��y��;ҁ,���|]�����)�>�G{o��Dv��q\���+���[��,K�襻J�`Țu��ւ���2tѢa����}���+�4�]�$*O�Ǹ,K����/!Ț�i��MoT�=�+����JAV�`�K��we�7��� ܵQܳ���U���ˌ3��?s���8�g��$���ǆ����`ǆ5I����u|[�v�@9����J�wo��ӄ�I�pI���י��� �m^ʪ�W�x�*��������30�#_��O��L��^�(^�*��	:��땴���/�r���`�V+���'l��N{j�a��A�B�Wxwrr�v$�/*t�f���B�����yCm(δ�T�kEP�;_[�>>�.�<flf�!�q�y�C�u&�_�2p)9~�@���c7�_��,N
���L�?w�N���95(���� pv(��57�5NR��SR�i�Wiu�Q��3G���jsv���K��\�"�����7�e�.%�z�3g���I�(�����I����t&�m������B�QK�	��w 	}u���S5^Z8��ھ�ПW��䖅�7��l&W1��}^CX����y�������+�1����'͞�7�]��F�{lb'�\��/c}3�*���PK   �yX �Y�9� v� /   images/2a0872bd-f672-45e8-b778-ad7a0f52371a.png�|y<�����k��S&[d(�d��0��%k��dY+B4��oe�	��Bc	ٗD�K����w���y>���^��a�>�\�Z����ι�PS<{��)tVYI���@G�h��d�nv �;�P�t��������}x���3%}'�\�CX��G �A���mm7ㅟ'<���V<ƾ)	�/���d�Fg��֎�*-ϭ�s���G�BC>�� 	����$L��k6�h�7��u��-�Ԝ�w�Qya�nyƩ|�&�dW���4�� 򏩡[��9�qz0��S~�j�o�~���*F��~��;�0��e���Lп~�%���v��������p-�u�`����t��������v�ϫ�~A��B_캉=��74�����g٥O�����Z�����A�����C��쩨X��)�b�?�ŦM�@�q�F��	+z`�����;�!���TdR�9� �μ۞���r�~�v���dY����k���C�_��/����K��.��tS��+�_9|�<E6�xj*��?�ߺMO�[Y�sb�y8Ҫ�����;��-�E��A����������C����c��
���߽�#��>�E!��%�:���9:���鰙�j��I���ky�xF�/��tZ�K��	���|k��g'����=��Am�
CSj�4��+Z�1����R�|͉0�����hx�p�ǟ�Z]���u�,�)6S�Q��*����7Ӵ V��m���n���/߄P�aʓ�(�K�ƀ@�Oޟ|�b��M�p_��L�ް]�N�c��:+DIc�I����71���T��L�C?be����=j��sj}¥�ITj}Ս���;��L�A�L
�F���3<=�]2������T�p�$�E���B�5��n�@�|��&K��l�'T)�6=/�u�!F��z�}��s��;~Q:Eb�^���Sv3g�7qv�1��7�
��_dO��P�oH�ȃ8�G��O%T�F�lBI)�>D�-"B��ӻoEG'C��Z�m�y;�#��%���\��
}��e�J�.��N د�rÀƽ�@�#}�!GU��#���ʗ����CZ�i9@�������R;�$��o���> ��A
->:�s༂�q�PW��ӂfç������yE)��ܤ�
�RW᠎.��LgZ=�5�.�y*���HY���"Df�;*��n�$�MCG��_�
�����<+r��h��ч�O�3�<Q,��3ӱ��NK �ޏu�k���8��C�27+enS_�7�ﾕ�)�?����R�
��{��<���y��-����s��5[�e���*�!�i|ÐMR�9S�>J�
�D�D�
y��f�T�+�y��;��HD���ӯ�&>�'mƳ���b$01Wc_���d�|5(����rH�pc����_G�GO�l���#�YԖ�vFM,H���h�ב@�Ws���R��6��GB�����|�{��l�5s���8t����_I��$l����)ތ�t��8�C⭢�u+���U;�|z��s�����0P�Ĺ4��o�B^�N�b�<C$��*V�
������rJ]��,G'���X���L���wg!8���Q���vE<U<�}c��+;:O�����HN�=U���[hU8S��2Ҳ�m�[(ҙQ�C�I���9�R��.�x�VF��H����GM!��c{��I����@��_�ѐ����#��GMR]��D���{�̹?�##!����k�_�%Ex|$���𻟘�xw_���J��<Ƞ����W�z@��Y�;���{9	=���|�����o˙�ן؊I�@�:��9(z�o�+ͼ	��∏ec$K�����F����@����=���75�^�XQz/`�f�i2C��3�a�o�%�g:Ϩ`�_�ֶ+ ��oQ0�4Q=�w;߳�>@�}�V��m}@�9��=���w�3$S��ʜm(ؾ�5��޺�L�Ѿ97l�˙���:���H��a�F1�F}��V��
σw�������!�\�d4k"]nf���$f�cy��Ț�J�gɽ��P�lx�`�PT��8��1��'��D�O���\,�;{�>����~�1��q"��8��K�<�+H�2<�_4�YfᲳ����qa���8� |�=1��f�e~�%���B{X���{�(��Oq��^0�@��!���+����r��O�_�.u��}.e=wy���c"nGJ��a�A�9��%#������|t�s~��k(���>���]3.�_���{.�����+��T׺G��Ç���u�o-�=`Q�;O��w#��!z����C�]Δl7Dv��O�_�z.nB����T����%�� >�t��t�7$6t�OXyWk��$F	�����2GҲ��}�Pr�W�D�����Y�K9�#rz$�iC����bb�R�m\����X��M<����w�G.v�9YEM���Q��t<~L�d��D��4�rzd�����:��L�?�Ģ����$Gr�:-��.��-��G&K�j-+UW�c�X �C���+��*��w��$����P�U"�3]�:>���^h�P�,����O���B�p��ĺ�,ح�<sZ�k"�f} ���ݕoqR��d"e��ڞ���o��]� L�#=֦���\�0����l���̪��N)��o�p>��ʓ��}��=��S�~Y�swIn��f������J�9��3"\����cz�vc��[A���,�2�"l[K-aU���<�=%��DǬ��5�� ��;��z:��^������$�oS��,�9�[��`��Ę�G#t�"��V��+ۧ�R|<�)�I)"<��+R=? �c����|y M>_T֚�
Ζ�Ş8�v���v��  w �0X+$�xuT8Մ-��B�yS��-Wyz�(����S�S[s�Q�x�NF���`�*��}���
�9'R06H��h��{�a��n�L�[ ���6�\���D�x�S�`p�B�ҝ�ٰT����YA�|9Z�^��jn֬��g����o��u;���pC���;�L��E�d!:�{ϟiY�B� L/���.�L�?4 �C���3���V�K=��t����k�S���j�F��'������9"Rq�=�o�]8�g?���#�����&c�.i��"N��DN�g`g��]��4��;��x�� �VC0-�>�΂��>��G]8�]w���D�Q�I��"����m���|j%�"��@��U��	ep���;Ο�)^=�_�O����Q��(��#�)P\FmѬ�L��J���@'�KG��/���(,v��-y��iru���L]y+j��{� v�o���V������J�L��B��_&���(��,���2ױ������� �3�}0kТ#����o(���VB/�K	�qRV4Ou\�,hG߫��o�g�Oz�z鄗���@r�\Po���#}K^*�M��xP�-���.�~ߥ���֖9q�Sk�r�YPR
���즕�ѻۅ�0'{��{���7�,�d��rGP(���b	v�g��7���Y1��[��8�!���Toct1�!�ˡT��Ŕ�j�DB,M"�4G���ʸ,6D��ոY�L̡6Q�4��7ȃӨ�������&F\R�i������&������\��	�.HWZ�����Pcv����5tQN��#i��|�	1��{�<�S�� �� ��n=���X����\ �;t�f��Ka�?�TAq��W��"cӝȦh0��AB8�|�����E2��S����:���ݼ����+�v4� �q&#�6vJ�[X|{~�����^)R�p<��]=/^Z��mN��"/�p�����;�� '7�D`S���٭O�\��R�UP8�������y�j�gR�T�oIA8E��� ��]�b��'������a����P����0o�J�#��x�C�9|��4~�׆F]�ab�SLC�<҇4XILAf�Ce����ѿ������<�1����g5��8i�2Tx:E-έV+x�H���.ev+'�.&y���y����[�t��F�2:���]ip�O�����\�$Q���T�Kd�J]���&f޻4����|���gI5@��~���i6�`)�#����|���L��G�m�0:6�PcgTK��(y����]�I#8�����P[���� dm��C�|�|�]n^�|�{W��7���>l��ųM�{l�0��M���;��択'E�_��z\��,��u#w���r��	|���&����Μ�P9�B�J�B��x�Ov���	�H�0�}��C��&a�NI�4x���t�����G��"n|a�����b"ى'5I@��T�����
B7�%S��I���LH�>���8EU�6t��>�H]��-��S�ܦ�ތ���GQ��������h�Q	gR u;0�Ú9��{��gI�%��Ol%�I����&r4:jA*�H5����9�	�V���E��~�����u�  \���HhLeZaA��9� �'TS��1>�Ck��/���l� �Qc�MN�M��w�x�G[O���Eƀ�Y�-^��+����+�Z���S'5�ݻYQu4����>�b>����=�I�[CM����N.���oʰ��t��{Y2�@��t3C)�3Մ�}QZHF���2#*%/��[���[�<y�fT�)��g����1����Ѝs�&���ӿ��R�n\���K�}�h�S$�ɇ��XU�הz�T�����m�]�&S�/���/�_��ʷOa��5�e�Y�q��Q�@�9��'�t������S�������
_��"ϝN��F'z�[k:�(�� c{�(jS�;�j9f��~�B��O�N�`^��h�k������� M�ͬ"T�F����\�)��|����Z�Ѻ���o��ͪ(݃{g(�8��Κq��3T�B��9��$=O"g�O8U�4j{�0�m2�vHFjOf�'i���.p����.�X/Ww2����-uo�!5i�auFk�mG5��	�F�VP����[#���Ċ^Q���D���S�姴o|5���C�Q�Y�ײ���09v�_C�)g�>���v�Fr���X����%��J
�3=W�G�i�P�}m쎋a�&�Z��d`��Ძ�����#�ܞKې��M�'��5���'(g�n�Tu��|��W�`��M�3�G[�R�i�bYY� �L
�����H��c���=+�`R�����b(�9bG�Ջ0 땴���h�i��u��b�>��6��P�ݠU0!M�Y� �:^S���7�?�$g' ���<�(�~�	J@P�X-�2����/�f��JEt"���{joY��Ay�K	�z�@R����O���Ĥ0w��~
pZ7�C�9�Ks�J����`(����9LE��0���B�d_�;e�9?ʞJ0f	�����5��Z\��
T>o�V"s]��l?���MO��G�J�8��;�B�,tdCkg����%ŏ�ڊY�N}���)���(�X[	�݉���Ϯ��ʒi$�	�ѻ�
&(��+�.����6�2�Ol
�ۧB��.<	����o�����S1)��$\�k]�q�1� ����w�R���q�>�"֮C�ϕ;��]�'6���ͨ<�^֌�ԗ�=�u���GE�Va{A@���2�.y/�+c۽mM����{b��ɼٞ�+{o��Ӎ=\����yu�O���3)��M�s u84��l:�M��u�f+"|֝��#����B��o~��*�	���G���p@�7KFP4a�ܥޮ��;�R�����t�
�!�~x�yH�N�Iځ����b=@>(���#0q�i��"֠��!D���:�7<�cj %�;~���u�-�*����fFZ}�;����sSł�o�v�k�!N������������'���"S��A�E��"m�J�ѯ�׈�i(��ށV[��t9� ��XܧG���g"X�iU���O�|k]���q�՜(�S���8Bں&N��S: �'��i�E��Ƶ�*;��#��;������6��� c�Rd|������fXZ�t*�V�U�㼀
5�_E��k�u66�6�h��#/\Y�-�+P{>j��[�=H����%G���̒��'��q�*6)��Y��~u����:�*����S�:� ~vv�]`���=�W iEݔꚫ��:+�]�4%���@�o���+��nZ��Y�/m;q7(��w�f�:Bގ
 GY�UӴ�݅�I ����>EL��A� �:K�犪$���4^޳�s���s�W�X���6��hݥx�xgO��@r}oJ���9Em*ۍHYym�&�I��.&��A�?�S��AZ���)sr�72�3�1 }ڵ����F��0ȟ+���yi$F���F��0??�
��d�1we�S�i�-�Q1qg�d�f��o1�8�2�;'#�>}o�G�U�J�7�CG�'�.��Q��|5{3_�L�� |�U�n��_���4�r����B��n#��q��rr�]Y��<�z _�U�2V�Kb����(�k��1b+���f �O�K�XǑ�8�+<Fh?_��H�c������y����Ð)��{WT�Zē(&��3+��v�7mG�+5�S�m�N.By=���|�[��\������o�Ds)i��|��/(���'9.:��2�@�8��,�"�f��6� ˿��+dPZ�!S�uu�c�5]�����^P�s)�*۵Bφ����[t",�y�Բ�͜�-h0XtL<�<S>�4k$��M���y��2�����C�4��dЏ�@�'i����� ̣�*���J)����=Xu[;��:a�K}�C���'.�GQ���ﲢ�E�X8�:��pY��d�aמ�:����)0���.I=�����!��J>	jW����x%:|s���T['�3��UQ�'@ 
�חu�^2qC�oR�R�
K�Y1���?��z@l�q�R��q�Ά��׆�(�#�O�hoy>�lR��54�����H���y�^w���z�Y�u ��$�Fvn͝�>���Ct��;�RДII��*�E�|�/�����හp�<nMLG����*�V�I�MLr��>}ieή0�?^!40L�ׯqx�ъ���[A}��/���L��Y"���f�����/��V+P���ͥOC��MLZ�g����y������#N�K��2ڌ�m���\C�O�;rMp�Z*H9��W��$�8�W1�iEP<c��H��An�(O��A���� �G o+������&�Ca �`��8�y(��b�l��7�}n.M5������ ���fF	��b~-k��"!=@9 �2�Ʒ�fw�<� ��S�=��f������Ӏ�8��{��h�ޛI�\������6�?�d59mg��ߊ��"#=v��x�]��%AL/���P�E���'ea6�>�?Ul1�i�
#ؤw�6��v�1֪#��ؖ�����U�z�b6���^%��d��{��S�Į��᧱�\\��Cq�)?��������p������Y��5�^Q�C��5�PR>��� ��!�o�&6��Ya��B�pq��ViM�������yG�Wkbs�Û��/b�5J^��u8{���J!棛��7���W�KoEAj/Q���dɤzG��!Z��6��>�G�̛�d��`^��r*c�I�4�／SR�?}?������,�v��Q�\�s0>����������
�U�D\��:�nl���:�ggN�;�G$��Ay����h,�B.���:[ �z�ぎKl-��8�+-@a٬7:�ћ�����.�F!r���y7&�hs!��U��h��1-KX�!5 �DĊ�l\�-;��L�a��Q��V�c�fYپ�W)K��6���_FͿ���Y���-�?H<·j|㈂J7�ꦸi�Ѯ@Ɋ�|x�:�R�ӗ諄Kn����>�v{��Փ�*�:ݼ�ck9Hu�[ �l�?�Pp���}n����0� �)�JS��X��<��h-�H;ƱUA,� n�&�G�Ĝ�i��`�[���J�w*cY 4��'`��G2�����8Qb�΋mV��] 9<=&����.Q[��u�"@�y���`���,�p��_���,d�9����sO����1>����S�c��cV��{����L�x^M���������҅q�ڷ���-@��[l<�����Vr�C"2���>F�Z�Q>�i��x�$�K�Q)D6�����F�|-�
C�vڟ^�����使w9D �]F>4�=lةpq�m<7��Z�Wb�4��D�FL�;.\����t��S{	�ý7rw/C�6Yz��6���H�uW�\�pz˔d4]\��=͉�pq;��E���
u��F[�5(QT�zF���;*,Ed�=�N r��
�{yuG�KkA�^	?�` �S8���h���dQ5��FA��k�q�So_���C�3Ğ�I�R�S�P��e"�:��!nq.G��Q&�@�D��ޯ��l��+7��<֛;�i�8η�c��K.5�' ���jw���KPVe����Qv�V&�:�5�Y�͓�T�EJ{B�����u�nO�G�2}X���__��H^�/�����jˈȌ���4�{��\A�׵f�e��Frs���/O<��_�!��6��h��9�ʼ���l��jY\�մ�������jzI
_'i�:��E!Z7D��e�&0�@u"� "���|�7+y�0����&��8���AM�;?>;�lqv�����Wrޗ��9� (�b�T$�)��s�Nkz�,���
 |� -Hq�|:�tdX_N��	C*t,��I��I��v(8+�N��O�����!�nn=�p"��� 5&� E�S0)�F���Ϛ��Q�)�H��h6�B�Ɨ^<.ER��&jҼ��H�}���v�.�m%�bF��k�{K�G��;HGO/��~ɜ�D���/Q���p��
jf,�8L�iyD� Q�0n!� |QH��|�Ӕ	����\�����F���u�"�Z��1jXb�"�p�{/USZb'L�N�PW�/����ո�%j������դk�wNi��>�Z���]����H~Қ���!�@�����ۚ�4h�yVx�f��2n33�o
��)��۱��^d����=�JO�j��ZA��p��1�� �ko���U��?~�翫N
��� [�x��X�B/I:��P>�����vh6/��)_���y/�.Q����5�*7o	��:�	H�D�(��#z9����l�@�)�M��5������ �uuPl�w��O���V|srX�V���[1����S�v�Q�B�o8E��e�#3hO����j�0gD�>��`��P��[0�"]!Gq�������}6�lk�9�V�5d�l|1iL���G����"S�P0iy혒ҧ�zd��'
!�m~bB�M���@,+�����i��[���P-�Ȁ�s���'ʬ`�>�F2�0�я�RL5�Қ���f�2�f:l�0����r�
}PSV��'/[OQ*���4�dj�����ފ�������F�uo��e|曺���G�%:���j��-	���j _������6�k5E�#Ĭ�Γ�{����G���w��4�N~���?�<`\�3}�cf��N�h�nӫ��B��.x���Ο��)�GW��ϭw1�m�S,��N�:�ݖ��i�Sk9�N�Ɲ:4(����j�QZO���3������2���).����m�]rE��IC��Q� �#Z`Tlnz�@S�_�����_:�3:�w#䍆��hќ�r��ڞb5<�N�ќl���"��h��ߌ��t(l�Ź�ʐ����Q+u=�B�������>�L�j�v����n��|������8�f��F�#�(�5|q�~��\A����-E���I�ʹ��?�3�]{���o��y�%�0���7���,,6�.c��,�鑷����,�����e�d�U*�������0�'���P��S�� � �F��jI\�C���aPP�\�^q޹�̕���-�L��\ �`��a��ĭ��@�R��%���>F�g��$E��$���Zh��1�|���^/���(fvv�c6�o��R�`��o�L�5���1�(��>au�	TJ�������=a��h�1���� ��No�nv�6���z|��#�K�2�J�c�aT6�yȪ�<m{0�q���}c�:�T�S<�G��u%9��>"����ǐ��E�A����1��~�X�v��f�K�6��yo���S?w��`�@y��6n6��j�?�M7����1ź6�b��{���gk�{���˳kr	�#�w"�L���cc9=���ϐ�ڛ%%��9�=%�*���H�W*B2�ݝ��(�K9B3MڴkҢ�1e.�}V��zN&fǕ2XU���I�ovò��~�0j�[]�64����la҅U߳yFx�'
�<Z\ ����>l�w�k��b�|Q��i��EJ�x���:��y�䎤9���/��/�]��"�W"���|{�#䕕��n�0K`Z�����5�K]������|�O��`�{�{�M����%�;8Tt��D�9�$�׵��rɾ;|(T�- ���'�A��.O��s�?fW�ӮXُ�ƙ�����8��,���ň?'��ͷFl8�u�#5��G�tq�#iQ<�{>���hct���UIr�$'(ad_�@?�Zw�\̨s�ۗ�!�y*m��E"�n�T[��%���!g�7q{��2�R�������j�P�,�| �����@�}�ut��0��<gT٧o������D�<�>��Ϣʢ'>nIɗQ�8Ǐ����x�(�Ӣdj���|�݌jNp�'d&Jc��j�����]D��~��?爠��v"F���ٟk�GZ��C�2Z�\��h�>�y]g��%����r셭Q� D�Q6�/zP�kx��h����ѡ�h�ڞ����
�� �U�� n=�����|���WS�<�4����dî�=�j��_��9���2̛q6y���Y=�ץK���#n"���?�>�	VTvx1�Te�x�;+�}Ҽ�d���l7�^�UZ�������+��k�����P�3�yWmf˼�w���$�~�de��r��򘁅o�2�������\J�H_��,Je���'��y��CZ��'�r^�R��w2O���3��ªS^����
��
'Ӌ�i�G�����^djw��-z�s���wد�,]9�U˽-��?o�\�kظ��փ��Ҫ�p"�Tϒ�ݠ\�mf4�	`��NJ�HiO��L}Ik���R&3�j_l�5(�E?�(-���e�.Ox�X�����Ɨ�<ɚ&���y���j��L��o�)�;1" _����>��{O�r����5x��-�q�I��/G������k�_�+|��9q�q���P�K_��KS�� �����:C�P�P΄d��g�OW�r�;�>�p?�H�*N+����\�������)����m
�r�a�G��2a�t�?�1��@Uw"���ͭeF['�[X(�$��Rֶ�,�TݴR�!����h������~{���8�a����黵'k!{�8n������K��%�v�j�|>: a^�O�Z�L��}�@pVh���d��q�6鴝'E	#�M�QV�I_�dx�����`�?��/�E��|`�/���ˆ"� AfK�IJr?��CoF5�E����B�p�C�m�Ҝ��u;�gLF�Z$xkK��U�\õq͛s�����tq_�i��m�`���f�q	H�O�{����C!7���H벊��2aBM�@����H�hg?4�uo����n?K1��ڃ�"o������'��tO}ضv���3�q[��}�q�i��n�+�ݼ�F��@w����z�I(� ե>o�0�����?�WJ�vx�t��*���ok����=}AϨ�j���Vrc>�f���)�޽b�+��2z��OfO�/{�)��CL�񰒓�����s	����h�x���܍~��շHI�%T�+v���Ļb�|;d�S�jLR�_�h�*�tX�00�y�����js���u�=�a �*��l��ڊS��d���B�j#�Fw_O�p�Y��ꬫ����ы��Vl�/��$�. D�n���!0ă��Q�c�;�!��kAA��g��^t�T2Aos�����Ġ���>~��g7p&���f	�/f@e8��M|�+��WF�;���2��|4�Y�eA�9�԰��$�mr�SO���0r���~�*㠧��ϋ��*���~������DJ,������6���Jr�����b%}��¤�!%��js<�_��.r:���h�� E�?�WQ�t"v+��M���w�BX�+�!�[�Q��T��ZY��3�re����?�4�e�A��E��y/��j�v:�j��5��މq�s��Dh���/�+�v��0�|	�����Zb7O��-�Ze�7+N�%h�K�;�>C����XF|P@��N"jU��*~��|��l I����y3/�����D��J������λ�Z���""�����|��}2r����W���v��"�i�
'k�7C�$I�;�	�F<�i�����iw�Ap�t��=�?�r�,�眚�6~��Ƀq�k��wƟA�	7Q��+���o+a�ׇ�m��̃���9��e�Ol �vQ��N
o&8�;K��5�
�g����2 <���(���M���=�FG4v/�L2����e'0d7��H�
��ڱ��޿<�ӯ''��oomc�ʸDD�ڤ�D<4�>m�L��R����j����Z�m,�15�8�	qS��/�V�k�^F�I[��~b�;ieȔ���x|�l]V��i�ӭ�$1�T�|�H:P!{S�$��}JKct��^��J��,��(��ڢ�':�N}�r|g�}�)��ء�1�͟��݈�]��2ŷ-��'�����$��?��ECb����H�(�����=e��k_T�W|�nx��r���q	�^D3�� S����<�	�֣���r$���[e��T�t�T��Jr� ��<\�x�#{j
�ow��Q�޿"-��sY���� ��`���;�_Y�I�]�g�폱�}�q퉪��~�bMD���S���,�3�.���2��J򯾪������P��Ў�>�mtK������������Ff�ݽ��Fv��8o% ��{�j9�w�Ԋ7М�����a��tQ�PM�ĵ��kh�^���V�C���W2v͹�� `O�J0yTpOf�P�g�* nY�ت����Yh����U��<�(=&t�/�s~6�'hB�QE��9V4���x��1�{�r���Ƹ^�W��<�I�Z�c;�^:{X���s�+^�^��3UL�b$�֯�%Q���/�Gذ��1�?��	#�?�gj�m���|]�"����@�ߧ�1H��\�������J����� ��"t?3�|����(��E���ܱ4���7����֣	�=��ٍ�n�3�L�G!n����7pͶ�5A���bNN.V�	���4���:��CI��p6Y�K|�K�%.���{�\��9��%�L��g��=�U���J_(9tX��m�w�sf)r���kS��
vG<.d�����l�YqݒH�o����&&�ww;��`Kt�y��8��lW�n���9)��]�Bktno���k�q+���R�V�d���.1�4��`���}���D�H���u��I���K��ί)�,gb���Ƕn/�ٙ�ɧ��(�0b7tH�J]r@�����2zs=���{p�oCN�j�qk��n�N�@�ky8�5g@p���&��֑j����m�?qȏ&o��tbR�?�� ��k����8E��X3��5���d�,�U�3:��a�*7W�l��>Ϝ�*9�2!�|/��Ɇ���D����ɉNw��������za�c5m�E�X煑�
��M�^8�ۉ6Ӡ������LÜ��j�>3�ZV��l}���kz�������R��*k��$���s�� 9j�*�:�����Zw���X��_C_(#��#Rk^�hղ]-\��y�=�w���G���#g�c���ǻ��ޤ-�Yh��:��Q��a�����bJ>
o�U�i�/.\)�{�`�1�@�婾ѢǨ����vo�����	_X�q����|z�I8���GwTo씴��<��[~"�զu�-8J).�!�Q[���ɦ���e���}E_�k6��7�=C/�\t*kʓ�=6��]�1w{ 㞟z�g}(��<��_IV꿢�dQIf��g�e����D��Г�x���L�Y�*+�c;��O�|/� )���_
�;���H�1SG�+�?����iك���{�4����ț���|�a�,�J���2ޘ˴���q���Ƃ���#t4EU $=ڈH1:�I�pg Hj�;#&'9��0I��^OӞO�NeȁA��nn�/���e&��G^�Mw3;�3�Rq�0볷�i��F�2,'�A��'q-_��оҮ��ܧ�d2�b�_�Xs.1�v��6h�4vy�*Yx��j��Е��O�[z��5��ӽX�X�Ҿ���U����yW/|a
:1�T��G�~m�S��-���Xj�z�|C�m(��p�}"�2,W�V��F�F��6��+G�L�N��sX�u��ğ(��>6�wf�l'��r�����m��������7ղ�S?�Xp��5�[w�,"��: ҈|
��	y$�3��Q��x���`�p)��J�u���_"���3�L(ø��'ܲ'`���)�ǥW���9+����v(#,s(��"��R�
�%+>��/�n���9�Bh��aS���ق�4h����_�m<�g�>S{����΄�%�i�f7GƮ��{q� 47G&'���"]A��)6/�������<ne�T���?:>['P��!��*��i>#�_0�}q"��"f�޻��p�%h�8I*��	��
}�R��j��I�NsI�����<N��i�b�F��Va~�8̄��]*;�8vo��"tݸ{+"{����E�AGm@��Zj @1��sk��wT��x��[J���>,D&�_�<z���T�YR���?���T�[��9[�l9}��K[]biw���ҕ|��XٰٛҐwiQ��@8�p���R��z�;*��賹*�?��q1�K`���0
�����]��{"��Wn���w�
ak��k5����Ϡm�nF^��u�wY�`��o+�V[;6?�gR^����UM�C�5�|U�T`�� |���]TZZ�*�L%�w'�3���<!��D��`>v.��]�I*��_�5�ʨ�h����v��h�����7��c����[%d�!A�: �C4_�dO� <n�-c^@&�F�h��OA���� :�N����Z�*d�ܯNg����"����gD�1�5���i��s6��)c�sp�斋;���P^iU�ɗ&c����y�s>Y����5�j�%̵�bU�53��Ur bM������!��h�&����̕��$e�����w����X���D����+S�)W _�DH��ö��R.E�R�]s����?vJT 1����ae6qb�h��K���8/$����9��c5=�����N=P�Ë3����Zre���j�A���lms�v�ej�����R�pGЇ}��VĤ��3FC�+i�tK��������A�J���M5�+��r�*K�>�� ����6
�7�8�۴MӆN�9�}z^�;Two[/�|�L��3�s,�L��w�+�|�Yot f
R5�⭻+W{<���=�����:��&��twj��b�IjV�<�mS����M]=5)5vbkͤ�`]��.}#��y^-����r�*41���|��_7��5��|1X��9���K�v �
 �{Y.��!W�-�n�tԦun!$����6�+/�A�uN6����5s���W��=|�K�'I���B���-��#��~�؇X���t��dem7�Gx��F��h5�WU�3Ѯ��3���S=og�������~`jKq��V{�m�d��ي.��Yȃ�Ln�J��������_�`�0 kY�{�!Y \�#Z�q�h�c�� JH�i�
�RYvw�.���>~�_o[D����V�?�Nzt8��f�*�2;����EuC��2f�8��������=A{1E�����z������Q\w��ND���������79*F4=���ß�
^㼐����iڣfDN�tG�`;��g߆?����vwTWYS|V�����X(�K�n�A4{Ei�6�&ڈLBd��]����Oa#J�n�iٹ>�=rT^5)V�8����hHMvM����p�����������VBm~ֵR��,7��M>�N�'��bhqӪAB�����n������fE2,;:Oa͹����/����2�$����?or�U���1��G��{עD.��5�1G�7N��D�wU�\p=���s������6�c�i��R�)�&�m_��Z5�����8_�B�E�(LJ�*�sV~��������M��w���e��Q{��l�F��i|ɭ�q��f]6;x���E�=��f�=�ɀ����x�rl���{�����%x���e�Z��3�qh��l��`��ig����b�I�p�X�ُTT��p`��_������.�xե�a"��y�U�v��� 8�����Ɵ�n�6�9R��L�J�G��|y�rY�Ư�0��q
W	����p�m�[<٫�_7"9�P�n�4b�3�� �[)sJ�����k�d#k���N$�����M���;J�v�G>f����1�c����M�g9�����ӧJXzd�����+ * 7�K�?PG�Q�o򨶏tv�@Y�6���.�t��C��K����Дp�ak�.o����e�u���*둓��gaãyHe�]<��p����i�{�~*�"���[��5��()�ock�?�&�=q�M Ӕ�*��֍��9<�<���9%��G��79����wҘ��������n�s��@�HO[��_H�^M��P��ٞQ�z����8��Gz��t WF� ��_����{�D��+���&�<�%��@��;�E�vX�IU)�9��Bz�r"��>��������ܨjMid]�/w�\�H\'D����O�&w��{����8j�1kU����2�����Wć$|�6G�o^@�7j�8�5���3Ƭ��$��1XVwס��o����2�VVa�bM�>g�%5V�M+_���s��%L��X��J�h]NN6J�|��(t�^���NR�wե����+�ݶ�������OE�'��L�r��TdMu���Y����p4V�zM�:�b|��˯|O�Z+'�`^Ϝl>�(
���Ù�*�R �w�˺v�Ś�5�Q�*I�������n��٭�����,uO���:��>�C��m\Z �i����=�;��-�%�����Ҍb�k�hB.%)QbEe�n�$Mt�r-׺�6�C5�.�B�㭪ȋj����h����3�-����[4�����G�T$�RZQj�H��t��$��0�!1:����t#]�I7H�`۽����H| �W�s���y$��̤�$��X_�j�5SZ��8S��4�@��>�W��;ل�]��jk��O�'Ĩ�C�B��/�}ۮK�i��r��nxS榷 )��r��e�|�(���; ���Es��z<~��$Ʃq iU�FL.���n������hB��V<������)�	���\�Y�Ra:�&_Ö
�	)K���� �V�N�rN����:�y����Pk��wUe�b�xA�U�h��𷦇	�q��f��C��x��v�m�W�d�Ot�L4�2�V03S6��ccAd�(]d���$��n4=q0�R�����������6�2��'@���M���	����۫��r(��
A��U,� ���p6�xg���}�(�[���b����ɪ��Mi�0�x�E�]�O�y������������y���)@1���J�����K����\�5{�,�A�=;�h��LM�K�g1�݃�>}k�r*�.g{�RG��d>����+pl���of:�#�~S�̛I(�}�#e�$`�a���{���X�z��ػVs�Ň�
���R�1���������11k��I��>�2��2�i�E�d=���������r��a�o?ǃ>�t<��5W�s���z �C"�2��A!x�J�j A�x��x���[�L�v�/�,SZ�n�W�^0�6/�y�e(^�p8���5W���m�0.�4hM�Z����~����M��2|.��87�D����	�Mj�ú#�~]k������g�>�}��ZG���/(�`�5�[VE/Tܕ��C�g\T��{�k�l'�đx�xw4��tY�ભg$jj�HĐ��6� �IIk�t�9	M��>=�#�)��ߏ;چ]�I��CKK<4bB.��>p�3��㻅�J�~�8P�J�K�࡭?
oϋۋL:�ހԢ�C�w����0Ι�k��cۦG�3 ��/*����^���*���_��w}�U�ؗ3�nhOX�U��l�E��W�4�$��ciEٷ��)��F���K�8�[u���=�%�r�&:�-G؏�dG#�R�h+�
^�پ^�	{���l�7�����U�?0�U�0��?�sc�{�o�x��vmE.j*����A�${��y�@{�+盋��m�!7u"����7Jq��i�	9�<��-�V��$����صD�� �E'Vo޿�$��T�R��W�Qv�|��cޙk6�]����U�+�H$�DKL����/�L�+�� ���]�ˠ�sL�湒���OԖ�/�Y�'��L�DJ�����-�ŉ���������t�շcΜ/��91U�ˍ�쮧;T�{<{�D�f7����?u��]�'uY��{	"��S;��bi���9)��xy�D�0X㯉@�h��iݎ��R�P�K`ҕ�-Dɾ���Ҟ��:�$� ��3��@�g4��0j��a�1M���J���Q����<�ْ���%Ϛ�|>��k�v�Ad��=)�cE
� �?���K>�Y�V|�ۊw�v.j�CJ�3��B�$��͍����<|����u����:��U�h�[�A�o��k�԰��A�fd��嶱̲l/u���:n	t�)�ZQ����ጩ*~ ͥ��}~@<yj�2�sQ�z�p����G'Y�����(�n>��u�N���dN�爫�h0�D҂��������-��tޱ�����(����2X��!6&Kpe�u�7�,�04�
���%ī{2�R�ql�� @6J���l�s�D=��d��m���'9kS~�L����6���N��u�T�~3�;�#c����<��oi�eN�^I���f+ܿ@�.�8���ύ�y��<?N*ʟr8�].5��x����$�2v����3jZ0*��G7�"��Z��8�HcNdC驢�|3�����L�����Rby���sh��	�Z� ������*��`��0�2��G�R�j�*�t��� �M	���|Т�X���w( {�Rl}��w�EB݊����Y5%��	�~�����^o!'Gt�]���8Wv���&�Y����]�W�emC�#�e"N�ʻJ�o?x����9Ix��r�
�	Q1��/+(k-w!q�7U����VƘD�Kz�m��2�����s�0��pKJ-#�焈1��7�]�[������8mԢ^���ew�Xg�t��#I'�ȼ�=��wI�r����[��3��5A�^�rl���w�gt���2ʆG�4!墮����Ӫ�P�#���6�3�=z��I�r�i�bn�0��A�=�jI�Y�A�XT��A�'��psse��.���h`z�H(�1��3o,/C%K%�%�A(a5��}��m��k�g����FW1b؈S}�ݘv���_A8?�'`�+2��&�:K
����7�U�{ZY#��Vx�؃>R���L{���y����/3^mj��%ۭ�NzL�����G�)hAL�b�d���G����E�N���Z �x�da�]*x�� �Mw����p�>�vQ<߀�æњ��*�3GS��ދ�M8�������j{5:�m�`k��ش%�2�\%_���#H�G�\E��XR�k��2Ǡ�����K��W�}-�XvF&�1ny1A�m�Wٛ�7����ˑXZ�4y�ċ���"����U��m���~cM.�g���ίFGf����cA*�w-2�TR�OH�8�������@��@ڹϜ��@�.I��ګ�nF��M7:'��r�pB�x�E64��?s�b>j8��,����&D;|�q�k������[��F�T�4<����n������q!pF�ؘ�����\n�a7]�K�X�%|ӚOz��ĵ�IL�Y��%ʓ�q�[7��S5��H�`�/_����'k�i?yS��[cT������ۙ���}v�z�4��B�!I�q�_���c|q�T�T�H���Ѳ����#u��Tg����bJ�/ݘ#G���l���gwc�gK%�[k�+����1�� <UB64(Z��/[lIV�[m��9pCB�{�<�:�����S��StB'�)�W<q$�����:��a�9��
�6i�nx���� 7"�9�
w/�>ysaC���>G��zd�����u(���U̧��u�b��G��ѡ����_:�dk�������NE����h���i���/j�GN���핑L�z�6�c����d3*;�7�fJ��D�����X����-����Ő�v��.��v���>#��=���,�d��)�j����j��A��\�,rVt���#���V|��y����z��bd܃�QGm���ޤO�8�{�����Ȯ�ʺmB]�ʿa4���D�I�<4������\wo?4�ԛ�ܺ�p�>�y�fxAz��Q2ԐjXtv������/��Fǭ�_�޴n��#���٬�)�6���7�h�u�jb�x���,�F�4W�'�Wc���Wf�+]�1&���4���_���7�.4�2�uҤ���7j�\v�^��8eIKZK����}��6�o,�W(�kt: �O9U?=��_t������D�h�~/�
��u�p�F���j�m�� ��c�Y�K]��^�5� � ��U\&�݋n�no��[,�&�C�9nO[^m蜒�Q�%�?z��"�o��v������}�=*3�w��3g���8���d��.IDz���+b�T�)�,������զ�p���	n��4V�|�����~�Mw�ʄ��ߒ��+�4E�y��6�$_Sǌ��&��Е/��]��E=���>6\~ ��fM��_d��	D��&+䩜��vbln6�;�jB�Z��(Q\W�5�,�ä��ho��+��t���0�0�|��O2V�a�k�r��#��
.-� ��y ��&��S�7�-�4P��?�3	Ч���+�g�Zm���\�c��O'W�f��hfYp�`b<��oJ�T���!V3(����G��N�%�/O���0�!$���ze���_
m�b8���p��e*U��k,.����_���f�p��ӳ�l�� �5��|���&xF�t�{`�a����P�K�������xߒ�T����� B��G������9H�2i��z���f�Q�?_!������TR��[�cᅬkDU8c'�c�+�&I������=m���9ec�/;�0�{�$��yV*�!f����t[����X����\]ޡ�`�������}]`�T�,�Z�^#yy�
�e*kK
4�N6-�s�@�C�Z�̔�~kf�sIw��w�޵O0	b�o����c;�k����}#�
������&�͞���n|v���Q48�&;;���"8.�Κ����Yr(����gRS�l������H�h��>FT��ן+��Fa�;X�}�y$���4Q�օ���<н���1������K��F�L|��^��9�D����L�����d0.n���2k����d��}E��2'}H���6����wc`u1�ܷ��Z��[�H�2�KؘZdD#����̛�Ͱ�.��~���'K��GI<Z��Xϰ�!��x��D5��Z�6��d��"Q���~�����ktz����w�w̾���õtO�̂n��f�t�z���|ޭ�B^� &�3�0"�āѷV�g;���tNl���qi�&��hͥ^yʗ�ʡ_g�C�l�]����}p$OY�n+[K�\kF���4[��Z�>�:�k0�ZG��.�k�=��-w�����ִ��K��9X�'���]��tD��x��$�K�3X�Ϋ.�8��Q\�n���·�SЧԿ�Yļ����k�Q��8L2:���QewK\��r�2+`l0���<�
�������z3fdMGP]��n�>�Ѱ��<���*�.�4λ���7p�w����9BW7��@z�vURX�N����jR2���� �gk�#�>��E$b�U��5�ռO*����EJ�,?[>��_����(�u\/�)�,�+�c���P�V�� ��ԕ�p�_�?"M�+?&���,���^�	��Z|��t��J6`�/�Vd6���+��E=��2��t� S��m�b�����_�k�Q�������.���	|IB'��i`���%����%3��EG9߼1���w�V��b�*)p,�)�<�P3Pp[ê3J��Y�*��U������v��R�-O�Ƴ���1/y��|'�q�C�a�f�5FD��(�Ɓ�'`4X���u���0�zd�ݛ��j�R�?��୑��֧Y�/vJ���{J'i��9?�`�����X�	Ul����#�ҧ�+������&�-�Z'����-Ɔk��"a%���J,O��j1�7<��br�B�r��|��i���	������/��m�����%����?�B3����0�o6H�՘O0o�e�(�dg�y�;��֡��M�d��{={�7�(nH�3��kX�����V�N�@�L�.�� ��_tf����T/;Y@)e�I��$��n1���l��ɥ'�K�Oa��F\u�.�؈#��
��w��Z�=�3h~&�b<823���,��S�8��@Q�y��i��z˵vo�����Q��1��3L�X5�, mvW0�'6p��>]�������@���Fg/ mt�00�Z�yżD�-�{�d��T��"�K8�ʁ�%��ϯ�O�!.[�n��﬛�5h����~�#��FT��z��Pkk��ǹ�_���iK���\��5�rm�u��ba�:?��`�/�~X*F��(���ц�q�<�H�I���T��jF篆�m�e��vN[��..�U"A﬒/ �+?=ν��Y����{~�A�Ou�#�BL\��G$O�.�\�O���V��_�2����~�)���	!L�g��U:�ov ��%-+,s��9?�Gu��1Ĉ0Y}���`?H1���3����^�q;r#3yg�q�9����`!��3I���.j�9�I�-B��w�
z�:���aƸ�S(d�9��Y5�Qo��s1�^�Bhŕy�S�s�m�$���sC3�<"Ȇ��B~զcw���Gր[�VwT)5j�XV���`�b2�/��Λ�7�
��cK^(Eǀ
�ڹ��Q�e��iT���MO!����zc��ް=)x�3~�v���.�֓�i�4 q����(� dx�3��b2�C������7���`�2��!��-t�y:�m�_s^��j�dTHzJ`jp����c�b0�����<���� ��i}J7�W��x�7���,�{�-vZ��a���#'ν��*}��6���]�+l�}١�y�S�:>n8�:��N��([t�w�l]��.G����Cb嗩��s'��XoM�>����6�hT,�8��ă�ǇJ�s!FLa)�֍��$��O ���Y�-�b��΂5N�%~��9o;��<�R�^���ڌ���oz�ȑ������~�����[��s�����81���r��.^�q܈�W���h2wY��.-6[9�}�	��w�<}�������hohz����Ns�Ӹ\�G>�V����8
�=�+��D1q���a-7�Q�������O�Y�����L���*Au=��25v9���c��s�: v�@=
lj%�dfxY��٠a��Q�"���J�S����"g�_g��ĜI�Ul�bIC2�2�	��la�z1�x���W������U���=m���+;4R��k8c���v?h%��)���K*vU�ĩ^�Ōx�❊]W��`�]��}O�m<�2`� �/�F�] �׻���v9?zENŀ��7;�7&'.6q�L�| �1X�|���D�d+�ag��p�H��v�K��� �i�� B�I�Pr\Y֥H�-���IY�ٶm�iBp[&�>�y�.Wӥ�]�f�l��&g��3�y������*8}�2RyK���ջ�+�\#"��f���r��+�`��k�;�$]�����>�MJ�Nr�f�8@��ÿ�Fn���t�� ���x�׼p1��"��`�)�{���.�X�=�o7�2.?S�v�2���\��>�Al]X�QEbX�]���f{;�\�fH��9!�y����6�lf����~����g����W��M�ֈÉ�M����AЉ��Kuf�׀�;gQ�?(�)��Q�B>j�s�7$:=x�V��2�����`� q��W�o�"�j2�T��:�Z��	���J�cZZ�kt8C�w��]������i�4;.��Mr}��N��i꒙��=���P깽
�����o=�8�-�ar�ձ~�V��-�ν<�-_ߛH�@1���Dߜr'y�mE�����Ǟ��pƚ�E�	�Xᎅ3���Q��@M����~�U#d�yGWܨx���F��yN�:��zƓ��P��'�H�md6/�M�����"�>����^|��﯆#�tL+_�$-yd';q>��ig�b�:Ј*��=I����e�Q�D�:�����M~�Ģ� <����s�ɠ�	ƣ�VYI�VЬf�wr�����ҳ��H��"������.���N�P=瑱Զ�hL�p���WV��=ޟ�̈x2ܺ{O�DQS��tW�ӑ��Z8�V�y�@���f�H���1h�Pw"A꺂|z�Q�`�Rj��������V���+�������fd}~����I���p�������3¤��|����nxW�G�ZOW�1R�韞\�Mf[S_��eI1s��5EY�$��ֵ� ��{̳u}w1�����Mµ���(���u���_����S+�;�s���2�A3��v�֤�R�A!d�cc!]H/ߣm��z�tY�PV��Q_����}O�k ��W ���Żы���旾p�EG3����ny�������:��o�P	����
�o��NƎ���8��MP97����U"�*Oq��K'�
���C�Q����-�έU����V�+�3�i���]�濎��g��`�=�_��D'1���Cۢ�*T�w����Y͠jŐSfN���%M�ӯr���n������d����kvk#�輨����2����@��O����d���ד����sk��~��xd\��T��m� �q�c�[L�m�[55r�I,ݳD�2O�:��A [?w-u�@s=U���_d�v@�̚Omo��L�S:$�AB�IN��3Bm)�����]B��^P�7<ǽ��p�CH�mCv�5q��=������z�x�HʨS���5E̾�SOަ����qX�'S�v�7r�@�D��e0��d��d���)Ad�J��(���#����z|�qVpߧ��Ae4~�b�'��_b?�u�|���J*������͊ÐH]�lN���PEp�U�����>:��]C��hG�l���tfD�h��^{�*�����4j��ɁW����-����Tn6��f����(�;MH�1��C���d ��;ɸ��k�޺Ӹ����"��L�~�D���נ���Q��U������r�$I����`ߞ�E���i<.�SoNK�g������㛫�o�����M9�̖���F��v���SG�V���Y����#�K4���ήf�K_�_WJ�R�\�z�Z�C�$�Yw];����z�B�?�lh(ca��"��Pe@|��Ŵ��^�����.q�p@1�~{�>��z֤Tm9+�U/��&�I���t.��X��w��'��F�a*gD��p]��_�o�7&��ˑfgA��N��q�g��j��+{�ɦd�a�"1g	n}�����:[B��B��9 �r�qW8��f]T�SIt Eܷ��TN��~ԯ�ޖ)X��-B	r��yק�H��W4���ے{f9m��?���0�7��A7�	�a���S�vZ2�\F�п�J-�x�U�E57�[�;5�>?2F0����W�DUtuM�s �T6%\�����X1e.�s�fMJN�$w����������x3��ዦ��dk�ؤA�f�G��_��
h����Z�	*W���;�Mjw��#EvL���4c9�Fc���Ӟ���ǒ�G�ہ��eK�<����&/���B����H���T�Ur�G���>�4`���K�+�J�o���,��Ng�}��Ϩ�>23]<*$Et�_��C1������3���q��` k��D��{l��7C���.k�֥�|���!J>�>�/���;B�8�:v���^�,��<͡V\i��=T������t�����"�Yϒ��D8(8��؏���_3ȩ��#�kQv�i��q�/-��K:�0�N��Ay���\���V��	��f>=��
�8���<�=�@K�D��6�r�:&�jl�>��Gx��W7������^�j���ӫ"�/�` ;Q���2с��@�hё27���+���,�ö�Z-�V���G�����lr1!���e�d3�$Z�����ܫ��*�#K�g���'tL�gOvsG8'���Щ-q:�l�G��kz*�v<[i[���*��8��D�ݦ��<?��0�i�����`�#�k�P@<i��lo��%jMH�����z̬��eM$0�&� �y��̓�\�h�āk$�\W\e�$�����w�8�y�^�������Hs��j{�p�!.�v�m[|��t<L\�p�ݭ'ʬ��>�YA�l:���m��_��w�6�M�S����hP�R�F�s��������%�V�&]Z�l�QuA8��ax(��Y����0J�߿��n%$�F��>�[1�`�2�� O��X����I�J>l��{Y6Qb^K���+ؒ�)��'_K<|�aww����bQ��h�d�C��Yֲ�qsO_�׊~;X$�A��%WjD-�|k��qd}H�{�R��	���97b�Ԥ��}#�ۜ��q��g�3��B�^��"#���^Z�� ~�7�_��3T��?}�́H�y1���X��z��5v//%3�P �ξ��c����;�4�c���,�J��Ҋ��ԝ��p�*I;���o����1���w���[e&��Q�2�\�d�6�vJdvV��Ɇ9R�;�H�⎲���}�Xc���i9o��%﹆B�?8���~���������7Z����@,g�3^ ��TI<t?J��Ȱ�e���u�jZ��Ĝ�J�Cj�p��݉�B�3�TPm��o�xN�I�Z�:��P5�Mϝ������>t�)�����K��^�����˘#ݮ���ed�q�K�����TLs�R��^��0	�W[L������e��wF�������x0�6����:lflJ��IG�ͺ���1-o7��NO9�g���?H��1�4������}�rh�Eg��V�GγC�c���0w�t7g�eZ�9��`!<�����ѯJ����ϴ�h����o^bfB��% ������+@ҷd�¡w�D��yQ�G6�pG�߹V`��r��?�T�J��ٙ����z�AV<&�-��o�3�Π�M���wY�ڳ��3`�k���2���X]T���{8�q������Ӭ�S��+�mg��iz����Mt�f[kj���J�S��PVMx=�D�6����W8r���8(x9���E�#�H�qP;��g�6��x����^��O8���OIڂ�Uw���)������n
e����F�����>'G��{"��A�Q���-X�	���ξD�ho��wAw����A��W��2�h3�ձ�����a����2��U�z�.�k��$'G���^$��0w���9T]ß�����Ŕެ��[�;�7�2�+������CZ3�N?�<�ؾט��R'�7��I��f$�!���[v	i3t�����ѐlS8�,qʈT���^G���D��&v g�B�0r���)�Q�ҍ_�+��j��7���>+�.|���C�Ҧ�`
�����������K�o�pY`5 T�7�l�<B��h�4'Ϊ�ev���v�	n��p�w�<��v�;	#1 &-��VO?^9T�q=�f���y�J:`>���~A�,~�?��)�?&��/o�m}��/�3˾uK�nz!F1u�e:�����]��;��x�E�e���i�zZ��� =�2�P�Sol�{$�P�v/g�~���Cj"�
}�bI9���S7��W#�W�P9��㣷3U����oV�ss����P	;@�(C�����_��S#����n�u)4B,��.ࡌ���15{ ����1i�( �xB���b
XzH�	쑆�ݜ��'�Ɠ��O�>	T"�eV����R�sn�T�����*}��wg�a�,�i�$y6ui�����[�?-e-Q�j���=�۬4�o�~�s��ߨ؃)S�t��3�"c+��	(j���c\IEvx���W����ĩ'$�V0����9��زn2��yry=1]���+�5ѶE��݁���$���S0 4�rb�S3�#z�"�'l���Gi��csFM�UHJy���Y��]�-{?���Nwy�=��#J�N����M֝�#��,�L�h�j�=���2n�ߙ]߁�9jp�D38�g4���mj��g�mm�-�D#{W;��BB�V����?��GZ�}��ۜ���Ǚ��-�;�?~�k;��\d�z��A����N�z�����Ҟ9�*B����]�G�-�v,S�8�H�	u���������f��ԮdX����g6n����l�b��F�pOӳu�gN�z�Dz�-
~3Bw�s��I���(Ϋ�S����-l�MaY�&�(��XJH�{��hvL�IL��9i�4��e/���j��5���󱮱U�oF)z��E�X��v�:z���=#�������q�3b��V���d�*�O�� 񆆊����yz�P��4�����RH�O!��䒃7�%���_�Ӭ�Y|��1>�Mc�Z����I������^<aʭF�yœ�T�~�5�pM�ӭ�%�HĲ �"��h,�B���{��WTê��։z��|��cg�sKs���+c����[e�&�b��Oo�26H0�h��V�R�<�_k��K��̙��n0wg҆�O�&�4�Y�}�$r�n=�"z{V!�+puw��[)N��[���=q�M�2����4�q�[�����,t������GTT�v[F��,����dN�~Q�oG��̒��.�������K,<���}�围��$��&o�:Z۫�;ԫ�Z>�\�C�g ��y_7�C`ٙ�G����ו�%�i�?��v�W��+�x�-n�צ��&��C��!��%P�����{�z>�����SMe�RD�6
B�9;��מw���JxY=���"*r&�q"U;B�U�Nh���n�Q��|���z��K!8�����=�e��11��LOC-�s�ulRL�:�Af�-� �����sy�_��!��b!x�e<�����=ۙc��x�Q�$�|�+F��B�؈B�QTѰ��|��z�0��8�(ѬH�ޡX-ǩ�٬�� �7r� ��e�Ƥ�+�tΙ�k�
k��)�7��j��)�_w���Z�q͏��/�ѣlX�D,[$��Dn�u5�&2Ne.���уx���|���_;���~���O�u/������gŚ���9j�ʴٷh>�n���2�>��p���9w�JO�w�--�/=3�?��<+K�]j��|U�^>Tc�������2sT�H���İ+67��q��2�t�'�F<i��� >(X��'+�MR7�1Y���o���9*TC��g�׌��J�ۂ�� ����n�7X tS���P{��o�ᇮ�G�9z���;�wUGO��zR"4F<����u�77�� �5�:>`��0{��G��F��h���U�ӱ(`��a%�E���9^�8�u���nv-��֕�LJq����=q�-3-����հ��"�n�ʜ�������C���4Vܤ��@�÷�[܆��V��%R���I���=`f[�Ȍ�Y����ky�1q�m��]!��M+EgT�+���"Lo�͑�<k�� ���>��7�I����U��l_9�oqa��F���������m�'������,Le���r�$g.����(�6 ��F����}����p�3�h�NvP�@5�m;��g�� }%)�֓��R+9�7�Q��q}Tһ��v��=����U�L���&./C|�ZEa�?�q�E��y��o�)�l��[�qw}6�t�U������*Ts�r}}1�����u�Ɇ���U��6�Y���8�r�FB��u�)G��;9 ����f�0���I��L���e��/_�>�e_��C�*0�B�>���{�`���)]/y$�а�hvR�2���i�poޟ�ɥ�x�L`�^̶�y�޾>�%5x:�N b�\�bs���_V&��*���+����v��ٯG��l� �jj�v$0�Y6x����QU��O�<��VeՐ�����d��ҚڴܣG5�r<��oz�U
�&�tt�L֝��ȇ1k���>{V ���̜�ק�|�����u�]��GM�%��`C^��Тy���oM�q�F�.���j�	`UN$��\7�K����΢�Z�fن�i_��̨Ɵ6���ݡ��_5�T��a�t�4�T���������k��\�S7}��t�)�����y�
�q��,�˼8��5�	V�S'1e��{<tn��D����n���x�ы�q�h�_;��Mig���F,>J�n�I���%��/ZC^]5�!�����!΃i"�@=�����ɸBYy=����u<����[�w ��ӂ�0UӚ�;*]��Z;��I0�T�(��%��A	LGKCD�p��3�5������|�����G.9����W����9J�:���bg&��IJ$��s��i��y�b��l�S�YD�}⤧�6�����X>ݒ���G�1�[�z�|SS:~9��W�]&sNf���Z�(6G�]��Uiw�U_�͓�][�| 6Z�S�)�ve��	KQA���4���7���O��7?9��u]���4�~���H�9i3�����]F��]�+L�@0lS|�a�Qm�ٶ�~!|�M������"WW�eX��iS*������܏�;�����(�i����ڽڪ	Rp1�V��Ҝ���ޒ��_�^�|vz����$[�KӸqC����P9��E$St%����A*u���޵4����r���S���8g�Sb�������̥C�س�K)Y��lLK�Xl�G��4�L}���3���~�oR�ux��D�P��q���J�2! ����|[6��Y�D>hoh�4�9��<�8��=��S���z�/h��o�+����{��͢�t!�\�5
s+��n���.�PIi����nӛ������j4NC?5��@�t��AA��ǉ�*�"�Ȅ���Y��ɲ��i�9���6lg�3������]��̐�E[�&!R�K6��sn>}���a����%�����1qCo_V����4�daQe3ł5��(	��vů%����p�Y�-��\kg�JZV:Q�h(Q>xs����Nl��&� _�W���f�5�7���>8־�4�ǹ>������,�]����.���.�b@�ޗ����Vr�-_�j+B9a�ߜ� ��wiњ5�����'?me�������\�4�JWejy;��R_�m���ͩs���fa�S�)�$t��v���k<��z) ;�B���ep�}��V)S)}.���iI|2qR�+v^"�T?	#�ɊZC������*��ټg��^:�#�3�ea����Ň?��(��uEp_��>~+S\��Ĭ�N���C�VCΏ���| �R�*Bе���s9țd�o���hs,��ۿj:7t.	A9�l��2[t�T�D�%��eX��;+�RtE�S������\�uh�T�'�༒�e�{b�]�dW�!���_�(n�/�'L�z ��UM�����j�{�����/	�q���厸y�6x��}E`H�+y)��=�����o�+�Q��{�~C�`��I�u�#�O�[ꥼ*q>�I���ɂ�ik�|K��yC�|³^� ������<�8�<��
	eg��l�N�ሑq��V�gPu��=��Ӹ����#ɍ�K��M8��>�$�r�3��k]F��y�] ��>�^�kO����)�㐩�0p���g�_$W �%��S�Cgo ώ#�I;��?�f��6t~�]�;�Z�Q��F@H���z2��Z%�H�:U�D^8#0�T����J�|�mVk]y�;����T�������5(�z�s������4@�_��������A[��&"��=������2}(0�:�V+�Y
x��,̆3:��sA��Mv��>��]Qy���3�ܿ�OR�;N�7��Q!�*fa��	:x�(`{���v3/�� NJL$���&?[ֈߵ��l��B��N;%]�6�y	Y!�aPD縣��2�8�\�RBA�k����0Z)!x'G��e�j�ׇa_��;P)I�-ݓv
ѳے������C]xBR�1uw�o͕�e����j)H�9"��������/��kp��x�.�情Z�8���~?؜_k���d��Kʄ�P��q��*u�3Yn1�9�78�;�^���Q45�Y�_78�1�wB���t�����W�Z�0�'����f	a+R���],<f�#���S����U�|����A5^Ҫۡ&��_j��8��� *��,;����^>jTl48�wl��|!l2Ĕ���H)W%9�"�Z9R1�"�H<���vi����Ƈcn��ͳ�}]�fb8OG���𗱣�u5����	��>TO|Q	>ӧ��/:6:����mؖu-�	v���-��ڒ�'�kgG*���E�?���?	ЙĲ�eN�	9C�]Q��p��K:m��.%�0EE���Y�}��2�-s���?j�̩���F�	#�of�u�u3�d���e��oE�~���P��7��(��k��8���0>�0���Ժ�����%-�x�@r>�!Ҍ�6/1ߋ�Ի��y� �yy~Zt���֦�	�?b�S���~4c���t}�)e_�Ez=���q�w{��E���Лa�V~ѯ}:���6�aG%�Q<e �D��������Z	K�c��_�tO�ts�4����lH�q��B�����x�'Ij�)����i(�L����ڦ�K7��;UVNs��'Z(�z��_���9(#���Ӹ����n�j����T�8V/[ܙy���� nߎU�u_�~U��a�
�ߪ���T�m�-Aq�Š;"Z�w6��� �L�{�ҥ���5ߖR�x7)�� ��-XzE��}��ܣ;�C°�/ҩ������}�F�ELm�e��#4���'�,/�m����(�H:%�s�?~�/�!q1�xR�g��o�Zٷ�ua
���:��Z!�Y��g{u`o�nL���l�N���b�*���Ҳ8��46[ܽ�/�l��HB�;x��4N�}lJ���z�:��s�^��[�9[N����:
����$�a�Ճ���6k<�v.����b���7'�,M���Iv���Q��� ��oD���
�ݽ�����iV݂�ͳ98n%T@��:7'\w����mg0~�':�͝8��CW���{*�lm);����F��W�g!+�N��(n���3_3E���܀����尙����n��?����]̞�>�+6�uG=d�>:��a���ŉ��!�B!���F1�K�k�!��#��n�)�$(���=�#����@m1Pb-"pa9Yr��q�ռ��N�E�7r����*��)������=[�[d0o�_N7�Q�02ͱ������9�v��ϭ)#�� ��Υ���9fZ������6�����^j�8�Hvw���/2֓�7�yf��g���5^��x��	2���?��Tވp2�\Xsz[�=��?�0^m�Z�8� �/��Ę��>�^	����:����z�p6���{���Ok��V{�*5c=S��&�7�75cEJ�Y�V�؄���$���x߿r<�~�����<�q?.Շ ��N֞��f�b��/�q�.QT^�����{V"���}K	2]���ݵ���=��n'��!���d�2�m�]mǞP�5�"F��y����'lytu�Z��4:�Ve��e�{�k��ھy$�ˇh�҃4�,�.�/�D�s�@��#Կ���/�4G="I�#�Q��>3���]^�q3�ƞ����+��3��v���E?*(
�r��$4w,� �_7?���1�>:^�Z�
����(���żE(aG"qr��:� ����I|ֱ�@��(��������6�����o�Ӗ�]<Iɽ�Rrr_�zK+�?Nx�[ֱ�/�N�=�(R���sd��D���44�r��������V� ���]�_�Q��M��e��G[R�a`�P���B�k�$����������|�S}L}e߿��\��v�6#3/�_������.#7�'a߫k�=/�!-�Z�v03�V�#۽�xυ�!?	q�wT�-���=5�a��a�x�ǭ��	ۂ�9�nK�9�!�E�ݸ�
\D�oG��saP�俯�K�YYl��.tm����p���.j�]P��H��(G��VB� ������]&e��EE�L�_aܷ`��D�����y�W\���P&�`9��+pp��w�^FI�[5�������睩�P��v�,�`���<�~�y��_a,>&��_N{k�.z�.j-��>��N9�#��D�Y�v8�9K���Y���h�c31ч���}��-��gC^�������簯P��ٔ���?M���� ��ߏ�Wh4�Ǟ'o���+S�4cf����	��P���� N,-7.�A*��w*�ź�U���QV瀀^�1�2�Ep��-[��#Ƙ�F�r/�h���/����������M%���>���{�9��D����S6�Wӂ����tM���p̑�լr����q�̦U#�BDq��m���Q�G�F>�N[P`��|~����.�0���2�+��c�=11�����Y�d��܄�����8K����sw�x��u�/;��S$c�$[p�c��$;;(ٗ<+���^]?�B���e	����pU�K��w�e�
�U������;*`0h�B���eq\Cq�ru�� ����^6�dX�S�,d�g��o�]�B6pd��f����px֭���ȃ�J���tO�h��xs~�\1�R@�^���\u�NR�SX���nG�Yl�}:mq�A�+z߸������=O����ޏ��n�ff+�ٟ�b�
�4��t�o�y��'�Տq�{�𾗹5b����o�ӣX�7dQ4��Qs���3�m�]�k"뻣i��\��"�`�
�JG�w�[���/�j�N��;WB	n�h�� =�}{��*��ғ�,�x.�9��L���t>̯�X�أ!y�ohҖ]�6\b���uڣ��J��.Mcr\O�6}t(� ��(�^U��f������	Lԃh4�VJ5W(L(�,�ŭ�c�X�{Sf꧎=�JS*�D��·`!i44�%7el��f3R����
��l b(�@��VF�'�k���N1I/�� �)��4=�H����5i�%����{GO�0t�v��1Q�� �s'Y۰�X	��p�"�U�&���g����K��E|-�d�@�6��uA� |��F���j�_bƳ0���=����e��)m�|����1(���^�I%eT�_��͗�iW�>�2As�lջ���JF�M-F0���}kբ/��à�p�Ѓ�_���4�m�Kc5@O�W/�_��������O�f�����KƝl��Ѧ�F��^�#�]R�u�,)�	��>��vk�AU����0_o���4��qa ��T�;�S�f��.�'�[��	�2}!�B�uZ��z:���jB����n�&X�薑S��"7�����R�_cY���4�cDwf�p__�J���:9X��~�C�'��J�خ=ag�S�U%���v����ŞR&�
��5ԕ{,������T��UR�v5�4����Q��vmh��]2�g�����u���ۏb;/(/I�9�Gx*x�W<Q�c��>['�ߐe~,����!�a���4���#2(ؑx���l�l����	����n�����-����B�X��x�yCy�a�g�o4����r+�RO},?����,a��0uѶ35��"}���{&��X�T�����|l\�[�z��q���Id�e�����Ϙ3=�_�K�d�,��[���{�VR�p�)܏i�r':�o��9��w�
�D�����h�N���w�_�����0h����$�<��#�B	F�wn�f]QK�Ri:=^�>����Ґى�����aW������@�L�c(�A#�'��?�;E����'�t�{"�V b��{�	.��jx�cw����X�f%$h(a/�:K엡���'�F9}��]V���Nj���Ԙ�5_B����{)^N���,�)�!�H�⌹�9�<�#T�zHԇ�cs��:zz���'	׆P���5��F���_e�(t���v�b�b�7�;鮪g��Wo�=��/vH��pD�:\�龍g�8A�m���f;AF0�Bs�h���r��z?�Q/V�~fR@�M��4�!Z�}9��k)��p(R7Vٶz�l�T#}򅩷�F{L1U�M���Ǥ���w�y�uv@�,�y���6f덎�."[6)rNșa�S�e�ڨI���>NO�D���o>�!<�}�Z�Y�}��/<��풮�v�D`���t��]�{�N�a)����I?/��6�[�?vc�ƾ��S{�k&/�|�~���>�
�<�Pv��Hoe��=y�xU��,�
ڶ��a6O���Ѐ��l��|�TM������/\���
,�0�\���~� i�-�#�2ُÁ�sJ���</�	��D�x^�Ϟ�/vB�n�b� �q��L���.�WrS~�O=֠�	�P��uV�`�<JӒ��i8n��LD'�`x�!���� ��3R�{�,�|Ġ>9E�#� qxv_=� �[<�a����,�Ԕ�˹c��y}n7�UM�lYc!����<��R M*������G)�/�O�4@4b*#y�ik7X�M�4KF������+�?&�	i��b�mא4�AJd����������8L��&�2=���l�ە�#�P�(��Ո��Z�[�O����!!�M\y7���0�~�n�2H~���&.1#���m:
O8�w�D��MY��5�]Y{C['�2�7�K�N-�0S�a⑾^
���2���E���Q֓/��ھ}�a�N�:�6�|�ݮ�Eg���\
�yA:��ҳ8�� ܤ�����:�o�ӡ�M5�.�E�°N���G%6�ka�K���[��A�3f@�і��F��j֨�0y�� �_Q���2�62�� ��������"�%vߋ7�(�����1����U7~���>}�E�]J�J�$���Օ�r��C����<d�M�db�����P�S���f? �Vt̺��l�ͳt�a�մn�<^��͒����I�&`b.l�q����9H�p� B�����ܡ�� �����:e�N]�Or�DXˠ��Nt�ӕܓ_ͅ�)?@ޝ'�_�KW��q?����;A�#s�ĆʨW+T�H����[�l��0�h ��m�ܸV���T*1&&ױ�<�DɄ�!��G^�`�א
&�&#ɚ�A ?p���)(��5Zm<���@$�d0�!gz��hҧ��s}/j��p\�*��RAc�%����]VH9�'P��
�:L�G��J.?�0ĝ�>����EHﲯĕ���R� �^c�y w��ՌF&���$�J޳Ǒ�Xe�f���:�/��O�}�u��9�&%d^WpI�ýu��E5�h��&d�߰kIIGQ� �]�!
�n�I�4o�Axcd5�|�еM�ʏ��;���T����ʱ8��������1)�O�+ �'�m�x#�315i�r6rJ��>#5�yKK��9��|t>Mz�
�'@�.������=9kI�]��>	��rs��"򹶱��`i汮�Ca�Ƃ)#0B��fIa������c���/5��eVZ%��7h��r����W���Fb{������gH���	<�֭]˖�=}uq����
گǴ�&Ø7@����8�O�gv��0LQ��u)��O�����VN�� ��T!"b���L_ٯ�GJ,S��y�u(*�`�b��y�4���w+�8uB(D_P��W��Շ���hd�g����IcD�1r},6�۞�nw]&^�ӇE�C��7�2���'�g�=��
�)������{��_�FX��:���]�#��ފ|U�����y:�O�5��핳�e��O�߅W�qKe�}���J����F:9�[�R��O�J��z?z5�?Uޕ}M-t#�pv7���x�κ�?�m�2s�}���p�4���uS�>N�s�;���6O!�����~ye��4YH�
�ր���֞�)��3�S���7��.l���c�Vy�!�X�d�t�����F�𣈞���/�k�1�p�~i��eĀ���q^K�Le�����'%�	7>���"W9]�c]���p�,~����f"�["��1�L���������2���<��oX�f)���o��M�\�2v��пߔ{}�������gIN7������� w�����@�S�¨�H#r]"��o�p@�v�7N��Ŏ�\J@;�q��M��A�֚YRg;κ"�e�_�jS����5�6{lܑ�	����/���M���`�(�τ����^� �.0%4]�U^a[l�'������Fqʶ��1b�޹v��?`#a��N8�Sb�\�g�nO�յ���4�ٳ������K��o�uF68M�콣����t;ɦC/�G�5_ب���-=������hc�'�f���ٯ�o����03��ۓ�C�.v������h�j<��7�5���7��=�n��U�b��	���٤V�\���Ц�O��.ݱ����������U�./_F&��*��.a]V�~]��Xg��0��g��LY��$�½�6�LSSQ�.�!Ǒ��[NBb����	l+[���L6KJ�P���-�-�ᲟZ1*�uJH4��}ǟA�cO�`BSY���jƙ{�$M"��W�I�8G���[�T*}+`�H�0E�s��_NTTO�d�P��mCe?qW1�Lu5�e�m����VI����h7�t��6S�p|��Yu���2&�;,�n7{���e�*��|����j�^wV9�	������$���vn�K���	�G��v��|@l�/��7���(��ZXn
(�K�mg���V٦�ֳx}ƶ�.�n��5�N~�XP�\aN�s^��3u��xfH�L�y`@�$J�$��d��˓hr{a�� ��*�1��8�������o
�I����	�1�?Ò��� M����Q��f[��1ӟ�Z�wC�s�0MƐ����	�./�_\,%�e�kL~��R ��_B]h-����F�� �,m�[۫1d�?v�u��9�n-hT���ZT~W?Q��N�4��Q���G���ƚ��cM*~XE�y�R=2	Ϻ��i	��Vݣq|4C���n؝�=�x�|cq��Ə50ن��u��j��#���۟��Рu��x�Ji�j�
��U���I�.�@�H��3��A|���~����)l0T�_���her��F�lk�B�=�=�$1���;1O](B��$�J�9`G���'<]����������'�^)js��Ja��K�-�@!=jZ���ϊ�{��@�:�t"&e��x!nD*��n�^�xk���%
m����/8�H��p�����'|r�u�4}A��yf^
1x��5_�w��R�T��Sŵ���Yׄ[CQ�e[�\��W�A�����D��t�]��+2>���74,v��휺���^�/�e0K�hl��)[;u�����t�j�%g��.A�c�NI J��|���I���:k����B})�9-U�����4l��e���k��0�RC�)�!A��q��>�F?�c]K��~Q��T��D�u��]�:��D�y#''a+T��:ڵ8�B�E���aluȘ^eY�9j2M�d�j����z�n�Ҡ��j�Y�ŋ����̫F�i-���Uc�U��l���l��'=���a��h�I���s2��iӿ��o��-[�������=Ql7����v�m̞rqy��Go�Ĥ��S��_E�{ P�4we����d!�;B���HK�z4�Yv��a�
i(�g���/�I�NeRc]�p�9/"�C�lխ�k�G���~�2��V�X�~�H���l:��|_�"r����A�*��S���$������Cc��(���oi0�QI}>ag���^6ԥ�@�"mԴ;�i�¡���3�J%�x�%y���T�KB''��k:��K�ݩw�za��<T���۴��c�;�%�]*�B���E�T!E!��lӷ!,15u�eCq:�*ؤ��Rmu� �Ck�˥�����4���� �C��f�Q��'�|����U4{7�r�m?_�uO��0ST�8� �:o��ȪZ9L�TrsԮF��{}���p�c��iF����(�j/���'�
���5��5��3?42Mȓ�_��3��뗥�����#8MnZ���Q�[����%÷��TE&�2�u�J:�?�.Nȼ]��Z㤼�m��7B�H���^{�����uh�߰���Yٍs�����ox��&�U���R(����0��������^h��ò��']Q���E�7r��9+��)Ƒ�'�i�����.uzF�a��(b
C�q�]��z	z��W(��?�H2i����L�ؼ����m�����_?.�-hhP���v��.;3"���-''����a"�CP;��~o��N�i�@ng��r���0��8e���y�S����`8��s��4��E�;P,���{r��o�դ�E��Viۊ� K�X�1�%��P�$�ed0O^&��Ê~.�v��Y�[�?����
o7��"`i�1�{k���Y-E[�J�%+ˊ���$
O�GN��2GN��uJ��4�����ѵ�4�UxxI?���/��u]4�>oe���X���������O�#/#��2�����*�ҳ�^�k����C���;b�[�P�%����*��=A��ހEޯ�I��y%��C��s���4L��m���RѶ,m�D�کѝ��������8E'.�P,f�oR���5�WT����@Y�����́���H��Ƴ�U��SN�x��-�t�]��_4��#���{�J�<���/o��ɍ҄��3T�*��n��q{<4����8�T��Gו�if�f�l�Yq%
��]���.��(w*I���?��lȇ���\�2�_�pӗ��W��uID8%G��K�p�/oy���b��)`��`W��n˳������Q�������D]ǧ|�@�j>�_[(�x�s��/B%�� ���y��|P�ҧl"S��wC����Ny��e���G;|�C}8����h�o���4�l�*8�l�؀ӽժ"nv�������9�b��m�hW-�������&�(ѱP/hy����z����.�$5��d�t�Ə�i��*��қ�s������JyGya?���DΩ�У�޿`Ҹ�'>��6�w4~��`�BO�E]���.���!N`�S�B�wj��cj���}��*�2��^�v}H���-�C�ѵ����ك�n Br�T����+Ջݮ�0x�]��ᛶNwr|�P���-��D�NN#&��)�`�
���6�5���ɜ��gg�[t�0������C�_����I��k�}4��/�w�jDO��z�����q�2��}0V������8�f�h�/#�p���0��k�,����ʅu¡\�6�CkOUݎ�9�~f�e�HIC�k�i�Wس[�zJ��|(�<9>9)��B�<��z�\ ��t|t	br=�qJ�\���NE��ܰ+��CJ���:���	�L�3Mi�c�*�>��N��*�z{�FD��TJo�1j/^�LȤ	�r� J�����ANi�ҙ��ۧ��:��:�^7�< �=3��H�e��	=�;�|��u���[c!,3�i����o�K�3=�m����Ҩt�rfy|eѳM���5����c�j�1�Б���E�7�������)�D�v��2����:�����9v" ���Lm'I����#��. �4� ]��2|d��ZE���¶�;HX���·g�Q��zF"���t�=t�n&��l�����F[С�����#-�_�M�1�(q�����̆t];KI�6�\�#�y����9X]g�d��U���פ9���)߼גh��V��|Ɍ=��?*Hk�\��`�w�ފ���Ơ�$fJ"��K��#�$]�k��0�Ub6����*2���a�M�'x�P�[B�w�.vv;"��/�is��s���w�YPcK3�O$�J��.��h]a���W]9y]�x�K�Xrp����G�~�4M�u	�CŤ�_�'��*%�X|�=���y_�����V)��ܗt�.�=굠D�]u�%ٗ��3�c���T�����ɰ�Ko�<�$���:����x�u>�*��v1y��m�{gQ=����9`sU�ƠE4!i�O�C}��o~ p\(_*�sZ�
�����I�./�
�R$�SN;@�/(n�>n{0�g�*o
d�r�o;1�I>tyyz���D��	��W���^x���~+�~S���X� 1����y�_�%��7�A|�'RԬ&�Ⳁ����
��Jo����j��|?͑�J�1�����������y�*�!T�������~0Z$O�*���2���d�5�CD�-���e�٧�!D�m�������wa^G<֋���ݻ��Z �����:���t��߈L0/&�N.�_tU�'�� ʿ�ƺP�}����c/�$׮��&K�E\�������K`��R��G�py�SFIt�A��ws;�Qo��s���ġ>c������>�̘Z5���GT?��<U�OI��&v����fU1_D���/x7;7��|����o�t�)���s��?iF�!(�Яt���9*��t�'=�Q�a�g@�4�g����8pֽ�c��T=m�m:���P�+����{D2��J��K�{���JRLk$]A��r��;p�������U%M�!�i��:uӢ�S7r����N�+OLe�R�T��� 8&{���C[|7�&+��r�]F3{ʫJ��ҰB���(HD��w`�|���ۊ]�yHyu�W�$>��c�`�N��:sh�bJ�(�{ĸݟ�x��|����u�9ZU���Mw�f�\G��}��źb����WJ��*埨�9�u5L���[���XJy��{n����k��)�-DH=|��l$$��;��~:gLSb@���5%��}v�*�t���t*�t3s��$_T��M���ۃ���u�~�&B����lv����I��2��=���>ɇ{/�Sq<��ģ�>x&���ͷ�S�94O�y͟��g��u%� �?��p�rL%�4��Fb���ѭLe����r�5��V�&Ɍɷy��m{��VG.�籌'�hT�T��P��)&\�z���U����2�]�cmȖA}e�К�d���BK���z����'ްVi06�w��&0<Ƹ	g �Y���ry5�D
���H�L@�l�����w"����TF�<��<��e�o=]�~4�����t$�3��ق,��x7���~�#7#����r��}��ӐH��xH�8��N�>ɗɨ���вp�*X,*W� +�骱)��~�r� ��j�`����`!K+F�/]�{ ���x���L���q�6�|���D}�bfh{Ƹ.[[���.KT�Q��w$�%����M+G��3��B��k?cn�b���t�������6T#}�����a�N�I<�1�����xJ]��nT���G���R�#xO�2'A�g���J#It�{���.ySfh����Z�?���3�I{U�Ϗ�הԳZ�����o�dgc�ؐlt���,ɱ�˸�_
�G���g=�z�k��;��B:4|�PG�!Ҥ����{ �����wR1�;���,O��*֪�PSorڦJ��(���������-B��^�%-�]�����k,��ʍ�yZ����$�/��mUn�Z���JW����Mջ������\�_*P���V�"��[xV��Q����x���zH��+�ٷÊ�8}�M�����ܠ;"���ݑ�n9�c��ob/���&���i����A�o�&=�����HC�Y<K�+�.��NC����q��ֹ�Ȗ�lN��8,��֘�O�RQ6�����9Ff�z�𔛗����f�9	W�\��Lh�%0�C`�&i�����"͗�3&�]v��B�C@��kt��a�Á��駚�&l{
��Nu
�ލ�K*`��fOx|S�I,8ՍQ$Ō�!�qT�*�'�����S�6�������`�L�f�&���3u}��D�@ה��v����j��Q׷-���>��β�N^�?�{H;*��<�Q����E����)���
ɗ�EC01�as>z���Q7CH9�������M8��Z��[=�<؅�)�N4���]}���l念��,��u;��2�DD�^	L�գ����O��(,J�1�x��ß�	پ_�w8]�HB�X���VڨY�x���Y��Q��H�钵�Q�K��8�Ak�y)��Z��ኼߺ�lpEQnͯ�<�����5��`����m"g����ԍg�4��O9�:��7�0آ�g#vy�կ��vL�/i,׸��;��q��f��td�f��������Ʀ���+�����F��|�r�$�C�u��b���[ѐ*6����z�R@5\�]OJ1)��.�����=���9n��`�7�����by�
��=JW���Pz�U�QNl��Ӣ���Jl��lS�uvg�i�<���6���dt(X������=2(3��(�]��9�7�ʵ;��:s(��$~�~�@�跃x�a|{!@l��������Ӳ�B���Y�{�ΠU��b�6��7��a�Cld�����f���l��}��X��]I<�D��G��Sr�}I!.�4�/�BRҚkC����7�lx�n�]_>�Iz�?}P��m9�g�(~���i���� M`��II}���ݸ;���(CM"������yO?:.@�B&D�����r�K���4�V��$�c=���$�죶b-2EǋBz���C�bhX2�j\����f��(/�V�j�`�-v%e�tb2�،S���£���}�:γ�S�E����5�Rϊ�{̛�,��|К�p���T(B� ��*�%?��[����" �����t�!h�?0.?��S ~����z��~5����N���F�$J�}��]_�+\RJ�l�á��>#
aw?��x�}ǎ0��:�}z�J|N��;�b�V�=�O`�v��o��2b]cC7�;  ����C��ԏy!9�Cy�n֍��P6=�K�)uL'�^�o}|O3^����/�\�%U�[�H*�J{�=�\l���ƭ�?���e��Le�~�D^�w�[�Ey�L�|	��i�w3m����b�q��G �G�V������J�����F���Q�yci���t��s��,�E0))�:g����A���{�;��x"h}�sn`�u���s�]�b�'�Q/��;�� u�Tܐ[wN���ȠK���n�S�'��o���3�5���_,Sb��M�O!G���u�*�MV����ʩ���t5ҷݨIL�fs��:r�rS׾�U|}h���p>r�}�:��E��qn ��5��;3�9��@��!آs��(`�>�=�`�q.;�v7)|�'�[9_<OҨ��Xq>S4O�d����5��k2����Ke���"'��NJ˔�G����g�y18|�YC��u��>-��)[;9�)v6�"?
Y��+s#b�S+p�t�?O�r y�����dj��d��A��`�e�L-��<��ڹv�`��J'�E�9<a�$��G�	�O��٤�9��� XU3o"j�*N�!`�R�}�[�8tqR�����&��j��D�����"�b�fO�שE���; !����¿��}$kp�	�(�� -��Ahe�Co:@�*��&0��9N?��$F�zG>#\�Sf��1�5J�I����^w�з�� �ĦuLs�&�pA��G�qq�`�8���~��!of���f��}��0g�IVLb�ݱ'dR�o��)l/��җ��%+��cN��=>A�n��l���rڨU�i/\����Pk!/�T"{WE�MU;�0;4�٬b_?���)*��DЎt�*�_�1�_#uv?�!ZPs��r@��5v6�d�SQ@׮����N��.��y��y@�F��,O�e���"�4���'9�b�u���X���D�̝�F�(�ג֢.Zb�+h�Ⱦ��NW�ͥD?��λ8��I�m��Z'�ɂ~CT����3��t�	��9�y��#���~r½�Zދ+,*Z�I�U����X�����}Ӹf���m�6W����j�(c���O$�e��H�O@�^�1�����N�<e�G�hk�8��|�� 6{�F��ɺ��,w�S�k �����s�����l��bx�~��l5_��z���E�b��XO��P*�k�ī�]]R__z��4C߰���B�h�4�7�h�=��Oca��j��ub]/�颼mu!i7�W:i��t�v.x�9�Z�(���(��x�	�9[���{,���;�23k��wo�$3"�M)?Wꌤ�S^�TٻD!���6L���ᝤW}�ͪ��]�ܻiL�KsQ��Ņ��L܆���#�T�}r��/�K7o�.ʛ��ZӰ��N�T4a&�#�cMWf\��~j�|���s���%� �(��#�5+,�z	�jނ�`'�jx�o��3�bnf�&�h�pyߢ���Lo%f"��p�y�^�}9J:���_�G50q��43ǆ[�؍np�Jz�Ǜ�s]����<��y�t���q4kH�v�n=�(q-�=CA}��(×ŢZ��h��ibjEej\=#0̴�0�����iAX���{��°�����m�+(�	�e�9=�:�St�+-���0p#�ͪi�\���ɭ�`�����;p?O�V�)X?y1 �K4���z��h���p:���s��_�zg��H��Rb��|�'{rS2{��������8�<�i�'8�#},�|D��,ec�ۭr4jo�Q��Pm������{�a��t�q&T��3�B�DG�$��6��a��t�I!���B���u�î�T��x��#mx#�-��i�F٬.�nc!*���u
�?�䛣��l �
�3"�?ܼL��H� �&��ޖ�oz��h;X������" ��u�;�ؙ��7�+Uͧ�d�nG��ӏë8�jɼz>S��k���}bY`�N3�Z�dI�P�n�ALP��Q��cSǞ��./���Ԅ���S�_�m��wdQ Lg1>�тZGoK�o��.�"��)��L�s���՟¸����I#L?��guZ
�U�-e.-��`Д�g]��݅"F���EG�|ڌӥ��E���c��L���-,�� 39��.V߾Qד5r�JM[��I���8��"���v~���Q���7�|�6~�fb���hEJk�&o�h�ɯ�	�3���L�����D�[�����B?U��':��*&�\d��m�t�3�I�	�$���c!�o��'��b�h���E��V�<4�/�y^��ꎒ�DI���qV�S9�K9�V�J�4��V�g���#��2�:o7H�p��'�a����х�`�t\�5뭌1^-���6[�l��vM�bsH�`��cHp3���O'��V�'�a�()�試�*y�̻� R��%��^ԓ��j���q�DQ	�l��RK��q�b�n�Z�sJ=��'�T�C�Pj��p�=�ﻱ�y\�ȎI�2I�$�/^�c>Va��fK�GO�Ԅ M2���.PS��(���R��vg��:�o��6�9�i��a~��_罹�Τ��F�A.�~�Z�jf$\�bˎ����e3��im1�Nn�:�z���?�5�9`vl�nJDT��$ʞ��_�|k����Fy%��Ⱁ�U��Y�Eܮ|���:�OYg�%�=��L�K��kh�O�9���x���� ��o{ZF�\�[�CNs	lǶ�c/�V�T@)#hᴕEZ��1ݒk�|��� �#�lS �Iz�BF��[]�0Ro�z�����f\Q5Eo����es: �PD�$�#m_م�A����~}[3�t�,9*����3�Յ�3c�Bc��%�W${W�'T$�� ]��Mj𳽤"��{l	���	��\,�]���0G{f��V�:6��0eP��c{���8��Z�]�VH� �*mߗv1�W�t����d�'q�.`s�9s����f�0[���w��å������$]x4� ѣ����h5���<fe�������][�%F^&R�j��� yr��aT�rL�������e0��z6��I־Զݦ�Wp�|2�@��ś�����Ԇ�9�(��ޢ<��9
�/V���[u�j�3�!��e����͍�&�;������M����x�%V`��t�-1&�\��RyU�^����P�C)({������I����u��6�`�(�h9���:��5��9VH�Z��E���I��*%B��[���|29#��O�(E��I�$�X�i��v���)7g���cރL��O�3�T�CK&x"S=G9��`7s�'8�w�P�cu�:���F 󜜦����}��px[�ֽ���4iJ"r�aqnٱ���|��q���K� =^)�
�\���kH�Ob��랼סiR*$�������L����J�ё9�S��s�'�2�����x,��nF�K�N䌊�U�Ϻ�t`9��z��,AUL�o�H���}8�:��$=yx� �I��R{�!|*W�h�UIU��l+�mS3D�[T��
�y�K�������&u%��c�����.��O�{�קw�k"����%�:<�yw:k��V�I�~�đ���rt�B�_�t��	���$'#�i]��O?��#ް�-h�[�b��gkM�u�=I��ڧ�κ*��O�W����:e]�I��h)j��ے�[���Ȁ V��a��e���'q�x%<~
^BIuE����'���T,��\I堊�6+��d�!SmA�=j:Ij�bwQ������N�Z����Ħ�`Y^�	���K�Xp`8�f�Zf�}ed#8;�|��}䬮�`Hj����M����;��I����Yn*�3L��#��7]�2��$|ߦY����?.E+��Ӓlf�tfUw�-"�x�2&(��1%o,���5�s
Nd.&V� ]d��\B��w�u�~(Q��ya�r���Ì-%�g�ډ��c��G���Cz�g{�	�ҭ\	@\�F�'�⯤&�8RT�G1���+���g�g����zZ���C�RH����)���h���������>���gm�'����4o*[��z@W=�u�Izhҥs�'�z
���ݬ7�����<�AOσ��)�<�y�6a�Q{��X�)	>��$L��-Ž`�z����R����	�1EO���y�� �G�F.���D6��d�g�qKxC�c<�m��ͰԻ�.��OzZ4ķ�����&^p]���>�:�u�����I�w;�zdD{�t�]T��(]c>�"�������(�/p ���e����*�s�psE�(�\l�+��:�6�[���q���®o�˓uW�p-�l��V�[��	�b��6���[��E�Ec�}���WL����)ܰT���^��x��;[�ߨu� ��5���x��q�o���$�1�Q�b#�b�V�M�������r*�(�b+Ϳx�� LLz��q!�x�͚��g\�"w���h�	%��sؙ��$��������c�ݴ�?�`��������+W#􈅗[K�ـ�p�,:�RN�c
nޏ�W��?���+k�x%k��3^2.��<_�m�3��P2�a�4�iyi���Yy�3d@�d�t�@,a�a-2�W籍�4���:�F������h�x��p�U,<
aK����|ph&���U�~H���x�0����*8.0�%����N���TI3��ZJ��R���2������ST����z�͸�}�@/�Q��w���vSQP]�f4�Q�}
�6�G�/����Prg��� h}P�%�L62���Xʝ����O1��M�r�-6�,���W�Z"�Y�� ��%^?�>��f@%����rڡFi�� L�89���V��=�3�����Z��ٚh��/)=z3\ʌ`)��F���spa����%�����$~�]�zQh^-�?�ՏqTp�<��+�\Iİ̳�ͭus����
��x	�����z��?5Nk}�?��m�����vہ���:�.p�ߦ��&p���#��)�z��Y���jŹ��I����?���卮˕��ی��^#�l��F�%�U���,�p����|r?o�Wԣt}c7(�x�K5��#]ع�@�ԕIW���46�L���p��ī�?P>O.d(�\̾�����pmĴ��q/T=��p�G4�?���{ ��
!��o���u)�Rx��_{��Hd�����8���vnR��[���r�C3v$|��H�Қ��Y����Ʌ���<��%%�/t���Y����mE������D��S�E@����σ�mj����k����9�B������[��F�fZ
��>�p_��{o��¤;g5����?�=���ƫg���O�$L=�c_�}���2.���Pi�	ii	��n�F:a@�KJ�J�A�AZZ��c����>�����ֵֺr��+W(���a���^�{A�'^.��z�ne.S���q�q@7>�����~,M��O;��L(����k���_,�f]�`�3@_�$�z�z^Z�_*�;do�Qq�j)'� ��A��E<!�_B���6C�U�xI��.�})׷<W�����%tN��8��I�hΎ���UyX������1^WԝE������b�S{C��A x�[zC�������8�
��g��}�]�0X�%��@�XܫZ^����>nk:�$�o�2'��J�C��B_���9~��4��`I��E]&��������[�7�a�;��a�Wo�E��j�W+6@��M�2I����{��D�H}����J�&N͛~��'y�#��1{����6ѥ�d���O:�o361�����v�A���y�d�R�yy7��Y��5�hm(۝�k��X�T	�C������]���l����R���<Ze9+�z@k��ԍQ��Aъ�	'����%��Õq��s�1�?�c#�E��{ϙ_~��#oWi��t��$w'q����q�{�=�쵽rwY2��	R\_���g.#z���X��Mz�§���"�b��%"�>���6�8\,Y�MO�]	зsಔ��%y���y5R�����*���>�o��UVpOzͨ�^�o��%�$�j��|�5���h޲��w8�2C�x��҈׺���eغ'�����æH��
z�	�x�tƚ�\j���?Kb�\%�FJp\脞@g������&��X#�A�|m�/��;[�e��Bj2'R��\Ěٸ&X��e�>�w����Qw�{}I�K�x����)=6_e��^L��_��y��ī��jc-
J���+ �wYR�1y�Ϥ�J�%�r�}�x��~�ڴ��Ip���-���fQ�Ϫ����G7�1�2��1��:��:�6\�6�v���F%���(t��(w�NuITY�����]��K�*���(*Oh�OO^'�J@X��4O#��Ċ?0}��9+���t3���kr��'9��J7�>0���r~f`�#09o�e9j���,�_P�p�z̝�����K��(��U�����4w���^T��(�;yG�U5��-S���F47�/�u����%�^�_���D��c �ak�Ik�nN�fmm
'�<J����n��}"������D���� J���meO��	���L�~���$vb�+��?,̙0��
�a�|���V�<8�O~��G"�;��[�&�_��t!�1M7��wD^v�M9𫵺�����^�do�V��;h��Z���pL���˜\:�?��AD�#�sab���ĹF�X!&�d�[�D9krK����Y�tŤX���HpH��5��g��,j��&���
B���� ȹ�r�����A\����~�|e���5f�������-�*:��/b'����$D��.Ã�yG�D�r��B#{��ԫ�eQ��{���B9_�	��A��,Ӽ��P�՗4���T"�3�W���.���G��Ki�^�&�e�<�C��D&��29���Cg�t��	Z
+��g��{�d�>Y�1w��?
��	�w��n5��7�Lg��_	�y��5	�*Gv�-�5�::�����V�9DF��s#^s�#��ַN�s��/�k�&�lɨ��a����5A�#���"RC.O+��F��'(��s�M���AY�@�x����1�.��*�f{��	v��R �Uk/��Qk�N4�
�����	�P�i��v��~�;x�`"��ă����,��`�MƳq�x�b���g�$o9:��w���)%U��2
�J�H"�%��,�XV�`�P!����w��kO|�U��ҪCw�i�Wt�"dB_렣hBt��n�y��ZH��d7=G��Vb:|�����5O֡G�6��{��Ey]���&�i?ЀgJƩ����wk��^�P�;���T�j����^yH�z�� �C��K�ul���$�P��V���s_ҀX�7�(�g	l ��bY<�<��$}cn��t3��GC���ߏ�>	�GM|����;K�s>�%QF�D�DP|�������AP��D�YUM�k�PRy�_��fB�S��@X�r4� ��=.��B��|�-1��D�)�[<N��i�r��P�[�>�Z�"���r������ơ��ʬ�6r!�G%��*���8<���2Yr:\yD�<n�R.q��V��ʺ��y�u�bCy�K�l�l0�?��@�7�1�X�5@�����eufkk���|V2�M�G5 '��#]�b\���i��48�^Ka	��8�Z�}���1D�*��"3�5Xl��F�b� q��yfD{'�M�;x��mu�t�x:�a���dƬ�Ȭ������'\ӎ�$ �����`Y�+��H�.�y�Sf��̀�vg��H�xE�m�X��3�$ >�y,��B9�aqUI���_-I����I�i������D�����b�������)z�g n��i��Z�h��<��n|]:*��	A~9��]��~�Q�Y*'+�Y��y"S�Ѻ�׵���q r0^�x��� �su"�H��aQg�gC��qԘ��=	@0F��7��S��|����� ��[, ��������H�cWE�)T��AC�e1;����d2�<�ǅ��Z�V����=U1�a����]A�Qx��V�1xB���Uy>�Љ?t�5�D{M��B*��*�V8����l�����!+�Q�k�H/s������4���y�{��LU*d�z��5U��@n��W������TN�Ǒ:�T{;��M�#M�T��4�QEp�5�i��v֋9���E�-
lV����-+������G�m�}/��v�L��迡iN�Q�CMB�7�!r7���ݤ
#c,��1V���Y~�7 ����?���F4o5R!y��PBB�qȎ%��O��f�{3�*��2F���{��X��o���@��K]�/r��w�I��~q�\��u�:��Z�7�#^y ��rƈ��iG���9Z��xٙd\��f3��t�P��#��u�\V�y2]����w.�/8�5O_�2)�B�p�JwT�%yS���褟�
�+_��`����[�����쓴�nP���1T�/M�]}��9���T؝y%9��k_����j0m�n��+��S�#���M�'��P�*\t�9���g�U�
{�+��9��nM��Lؒ�X?��	Q�i����N��>�n� �w����4h�!����c�.e���#-7e���U��<�Xm�7XR6��gU� �pF�ߟߥ!���$_z>	"�}+M���QGZ2k:�F�w���8=�7�
�������bp��nuLJ��y�߾��|A_9��L������
�X�s�x�1�]C�uΰ��d��L�9+�0*��l탄�7�=���벱-����ۛ��Z�"YM����L�h�{XȨ+�E�s�L������a��]IWDg�ygY �n%ɕc+w�+���sl/~�4QJ>�.�������bg���r�L�5�`ҏ+�ԑK����K���$�J�j���P�U� �0�W� {[SY�����ά�D�khV]�܇����{��U��V%3�lT�l�w%k���9�W�h�eA����w��� ø���#)jR%�0O�e5� w��x�&�SeY��9���r:�O\��j�>u��}� u�D|�r�
#7�� �ޕ)�D��SH'C����i�p�B��ƱB{Ǘ
+
�VokK�*���j?��ň��hLoX��Qe�'p��&���MuT�͡U�J�#!~�6��w�k����� �s������L���R�Φz��F��
��=8�*��E�T�Y���ܲZf�}ss)��JcZ�Ͼ&?]z��>��gZl�mK.P�@�����ƅ5��lC�0(O�z��q��?��|o@r�.U��$.�y��+��.]^fD�W���}�뾟�206/
�=/{#ANh~�C�"M��$�i��������57�����ͦ_���ڀ_&,�l9^�<�S���4�ֱ����r7��8-���B�NI��m��<?'I} ��#�|>�'j��w�;h����V��O��2�,$��ߚ��hzE�uz1��p�	L��L�D�� Uy��c?�LH k���F��o��׈
��] ס+�,���@KG��z|�l]E�u}��#g��@&��$�k�S����̓��H�������P�']��a/�z�T�^4lֻ�(,),�a�ߕ�w5����b�/�I=��m,�cS�;�6d��'}�8 �j��zb�:���@��2���S�7bh6F}�l��o^��vIz� \��cȕ1 �7�;�	U�:!OȆ�=[��x��u�x��� �T�넱����o��ސ�O4gb�*Xo~y�)/糘r؎���5�ᙒ�f��l�O�:��>��o�=���]�N������/]��|�ld�ểK5!���N���m��\P���;L���ca��L���@"!;�1`��X�z���'����p������%���L�m\����U6�I���4j(��w
z��eF#4���s�D�΋+�;�8�����x�`�'�-
r� ]t���:S0��#�zҁ�������H��IϡLԚ�-jϋ����:�,	8�Հ!T�,�s�Ѝ��V�1`Gq��dcǣ^!��m������kmA^vL�4�Q�d����C-�^��w�>A�J�=u�|\y�Wy6��/�4�V���F�d %�vL[00
���%�4�^�Tw�T��ϱ*�;�8I�p�`$�	����dH��������P��Gã�̾ �
FY��PHk����,AU��Ojx��y�M�2��O]V='�Rgyk���*�em:�����"�uj�뻶%�������l��N�	��|tӐ4���W��5wm����8@x�"E���� 8D�"3*7�th8�����ZW�����ed�\Gp\�}TR�nǈ Y��5��QK��;��κq�;�)2a~N��=<�q��ĝ'U_B�KQGtFu��m�y�>�K��Y ���6kcoT��3Cu}�V��=�-�g(�e�z�q�nĐuA@�ܼ���B��5��,V⡲I篧��ʱ�Jtn���|1AcN
��cK�*[���4�lMx[���%���]��x�����哩Ŧ��-
ϵ�p%V;<�g�͕߱��"T�A����8T�i�y��=��m6EŹ�K~i���}e9\^��4{��(f��m�o��k��7���>�w:���ݻ���1{=��iE��(*maY�?��U��3��g�x�UX{"0i»�������]!���C��K�^uaZ�L'W�Y�����3�&=s�}����ǡ�N�\��)�Fp�?p��g�*�9O�4�aQv��0y����|k�9�'9�QQ�f*�B�Lt���b�$��hb��T���$�<�	�X\����Q�W:Gk��h;�qu�tDLrX@]�wO����ɹ��&���B��i�����G����o��m��f��.��l���|�in����$틕QDG���D���>���%2�|e)�G�d|4��q�
���ʑ���4��\t�R���ŝ�w��7Y��C	��o�1��X��N�i̜��" ӄ��g�LwsD�� !�r��hhBH��XHdqIV��5�E�g�4r^]�W��q����$Lw6�A�>�1̯�OJ���eok�^D�J@W�u�*+^��cb�x?��uu�b)T����	�Q���^���f:����6�4�[M���aUeԎ���fZ���$yZa*��Q���݆/ױ5h`NZ��Y���Qjy#�(sU��9�K�t�#'sR`)��#��j�G0)�����C�b�!Ƥ��xM����8` 7\ϋ�ZM�Ђ���� !��uZ��O|9v ��LW`v�E��՗qi}���+<eYu����T��i�	kǕ5U]����1JFͲ�nV�/ڽ����sq>F�1�%��[ �$0pW�̮���3�	P��E���b�4�����`)*�
��˚pRtK�|c��w�d�u6��g���ټ=�oki��bm�.�{Qq��~�V�v��s1�b�'�D>��?���á\{��'��P�v<,*ą�2=����V��駔���o��vT^�DSQ�y2�ARa�����t��oG��w4�t��o��9K�(��#�����ߪ!�����/dw�����ۃ�+�G�8ǫ�3c�ׇ4.��� ��`�� �a\��J&wT_�-�z�2-� %M̌�1:���t5�5^��y��}�0C�^-4UQ�����0m�����m�@}�N��s*���1){�w� ����ӀM��N����c��N�G�A=�`BO�\�V~��{�[��@#7%�LW���Є�w��DR���H\�{p
ɴ@!�Pmf�2��7��kB��O.	Mc�{��tDC����O/@���� fo����Aa$7��
j0NRWvbm��{%�r�r��W6��[������E>�g���<��u��qm���=b�w� ����Ey |�Q8�2$�Q>O��ƅBÑp�Iy�����h݆����|�~�@���E�潃�j9S� ���.�3�Ej�ā%;��K�Y<Β�v��S��?* lq���
L���w2M�Ƣ��L��r�U{��l@�$�����k
�(X[34eC�|ag��켎i� �?	H2�Б�F��P�u�J�>��
�	l��,P��$HO$t>��]�uw����E����8�\l$_Ŏ�f�-�xQ�1��^�A$����x0�$�z��W��)P���)�35�5�ܮ�z�]��,F@����o�T�T\'{��z����܎�A:C�^/����G �Ԑߩ zͨ���iz�j�_�T�����3��{͏!�T�g_I#�?��}mO����t����M:nX�KC 2�.`���0y���ccR�g2b'�� �0��Y0����*䧘����{�7��,�!U
���\�L����t�w�x{��	�es������\�AA��6�yj i8̣^Wx�w5���nm��iW��D��v�ղgg�||��5$���<���T7Q��@����;��щ���m<�^}��̓,V~�L�B%�X�|�k��Fܿ#=�~ْ�ā��6,�b�d��*���#o���h�3�|��A��\\�}g�xF��sߕ?L�"vy��~�����[A�뇲p��4�`�
�F�_�1�E�k`���C�.��c�gK6�q��^R�N��d��d�0ͫ�Ψ��v��)h����F$?6G��>�C^d1�����{��,�jܕ_�!Xb�1�t~5��1�Ur�)��o�i���]���~�6mb��)�؂	ELj}����R����'�E����0�HB���V�zD d+*�[����3���^Go�׫u����[�+o�h���}���*¤b��A$<�&��]I���!z��SI���f��؈":E��7����\�|2�"�5tD�-{�1�y��ysA�h��:m�$�L���$i��:23={�'��T�N��/����.ǣ����y;LsZ�U��1m�( �Tb/��jQ��_�dȃ%�J�#���vfK��&�O �99�,oV����
q�J��O7��˗�Uk���B��֩���>I83�GI�%i[:��2F�2�-(���@�>����;��UiCɕ�W�x���7Ѥ�F�����q�S���~kϽS����ќ�C�}��#2ZȌ�rSD�	k+�����0�p�i���(N@�=s�o��f6	y�V��T:��<�#'��~����넑�|?'d��k�NK��LV�!��%�|l�c���f%B�
,�V� sO}NVv�\V��Hh���3x�1����?w���|}���e�Q�e�q�G�(,1�S>2�9o5�OC��ؖ�����TAL���a[�c(�	Y�]d@�L篅%0@�Ű�95���ɹ9���(��:#�Ϋ�Ź�V}x��=�3�;Ad��&�;��DZ콚����'y�F��-��E������@���pxΒ�t@�>TJ�g7.���]ZL�ǽǦ��j���=��C�������ck��)K3���W������
�]���q���#.1)�/�D�,��C��=�H-P�F�Q��l�k���-�	@"DS���@4 P���|�"]���Z����P�8+'
�^μ�i;\����=c�x�茩�NL>�O%:O�yy��5�[&���Z����&�T���(�
��Eǭh.�-� w�t?u	�j3#@����1��T|��gҲk��NgÀY��mQ4��*�##��k)!��^�ҁ�W�Ou�l�1�����aCx�������-R:������o&�^=&N!:�>��v=������k,5�{ך\jTߎ����s>�!l�S�G�X���5?��`yIO��-�Nߞ��Q�z/v�Ff ��Ц�	��wY�P�����K�_���� �:��m�5GM�� $�`+{j�j$�I�3Z�:A�.�qi��2�K��d$�ҙ0c�哦�a|>�s��X����,A�4��eR�k�Ć�`4���*륝�y�'p�f�y�E�X?bk�[]4}j7-'ˍ# W9]8��Z{r�f�{����*�${��蕲Ӭ�y|���!s��B"K���J�Ԧ�x���I�M5�����/<� ��;�d��­!7䥨�Bx�~������e����I�#,�zӣV5�8#N���?,ī�-A�d�����+�޽2-�KqM!Z��A�w�d͢R�[��BvbQ����s���Ĭ� �K�n ��D��hQ��J�6�{���9���n���k?�!��r���]O,��?�ʛ��]�����C��G��Y�p�#AP����=2Wi37�t�@�8�����V�Qط�./{c��A�ABi�$L#�h%�nh�� �/�BJ�����"RDvk*	�]刵w��w�a�%��M�[}O��<�.r����nO��#���ڟ\,��H|���g+�9�j��b������$v���}5^�[�-��hѓ�cLo5<���|�����"��[ �!���u��뷆R�*>eDn���*u`~i�;tY�kb]dɮ4���)y�H.&%�Ą�!�LB_O�]�{]�{񀺹����y�L�r-=R!�[��������G F����`$��ۀ�E�ש#���� ϽGfkC���	v�:$
��18�z(}�H+���8n��_�Ofh[�k
��@]�D���P]]{q��G�Z\��`|$�2�ѓ~琅K/i7�=i��"B����! bF���l�g��|���U�X&�K ��=|�w�l^&%?+��AGօ���Js�8�u�k1N����)ݿ`|t�	ky>N�����qۂ[>r��\�p�Y~~���lK�w��u����XV���	Q��[M(Z$���@�僧6�`��8ʢ]�5r=��t3�ڸ�L�Q��qL��I������tS��Ry\��(+k�:�g]�t4��i��rd�8��Tpd��q��m[�&��wp!��ĝv�Y�����tB˝s��g{/��ح�S�}���VE�Hj��4 t:�4hɅ�Eu�9V�ĩ�y�;�3�;S-��/Ë=d��BU�l] ��� ��*��y`}}ZSe���ǘ��3�$���$(����^x9r��j�a��@Q�"T
AK��:m��z��pyg2F�ߋ����m?����[�$\�i����^�a~Z�r��Y	d�ѳ���WU��	�V��ۜ#Uf�M����Z��cڊ��$~v�H^fq��8��l�@��ws�o/
臡�c�d�� ��ku���Iɨ����h�,a%�)���e�@���IRm�h�ȶ�JF��8����|��[fͧ��@�׬H����-W?;��I�p]�#�5$!cn)3��B^$�ߍ�������u����>��t��}�|�
�I�J��i=r��]ކ��@)�r{$z�L�ՓaAk��,PP�����H�S\FŦ��B�:�d����� ;�iz��}6(�ך針��kq�y���s��o��i܊n���}�)q@Tj��sā ��Q�ED8�(eb�����Q�W:1B�\/ �Pn���>�Z��>x;�۽�=Y�����	�h8I.�幢�D܍���6��E�4�Zb�<?������6��H7�yz�z�yMGA2�U<� ���)��h���JD`v��W�N�Y�x<��3���jMI��b���D�*�h�([1������Y�ͨ0�\ŨT���\�  tb��r���`*���fǀ����b(7��5���?۵� T��*ɕ��@�Z�Pp>=a�Ь�#��mW��B��J�@�|]%*����魊
G>M����J_�yF̞�Yֶ8�qZr�b	{~d��.�e`1��ǻK�<J��h��钫�S-�xF!�:L\�]���B��������41�	�o"e�Q���41������ҕ%$:��S�{�Ht�ʙI��J�m�km��/;��ݵ`�!�^��Ԥ��ҩ�}n.reF8S4���)p�a� _�m��c�9�z�뭖�eG�K��6xAziXS~���t�(�Z>�rP1-��V��n� ~�P�s���I��pO#kݓo�im�8���ӏ�\�9_9UrX�Hg2��퓅���8�5�����$�؈�C�ݲQ1(����/��?>��('[{"$:�*=���&���C*��f��.<fR���8���Vx�7B�g�q�0��b{n�c7��2ş��N������/�K��g���_�O}���R(������������w�����g�L�q��V¥�/?iƙ{m��~�Y�@J
��n:�c���!�\������o������¶ۡ�E-��,�R�|Y��paT���}��p�p��r��">�]�A������&5.��n���L�u�*�u�po�K)�{���#��s���gm��x5�5=����*s��Y��H��DT���7�YX���>fZS��#��g7��m�!l��4u�4_�C�]'�f����B��"Wk��s&��:gyB;��u�˛�h*��V>����O�.���uz��L���6ƫ���$=��	%����yh[���W�-I{�0v���k�����e>����6�ľ��ח�����^m`�ʅK�*��/����ݟ��y��
wF4�Γ>X\��9��8@�k�[z��3�Y�����AC���E67b�����ۅ[�����=���؇I��f�,����_E4��^nt��.>�|g/�h�Ǻ���tsi�7dB@����B�ޜ���>��H'�;r���9S0�b�`q�y&���km��ĮӼ�Dh�;�y�a�_f��A���d\�L�S��yR��/~��n	����R����'���L��-
��z��R>_
-�4:&p�Pg���?��w���Ws_��m�����zX��G����i)�n.t������U��իE�gn�PR�T���Yy������R���p�Hb��}#�p5�!=���z�0#�>A��?`�����,�OS)X�I+p�v)���'g�{v��<����rr�pTD�m���^�x��S���s��X	3oƽ�	�/��΃���dr7����V6�!�[��ƬS$���4�v�"�7�^\�����x�_���ۆ(Ÿ���qR� ��yg����ޓ������o�F_���i�F㸯n�}�_ծ��z=���� ���1�N��E���b|5)tC���#���~�k�xhi����恺���{"��sM��p����yۣ��������/��oʹ���F^�kt�H��]v��P�|� M?�l�����&)�E�>�i驛�;_}�^�[$�l��&k�݌�->:=�Z�!�SY��]�����ZT����D=2����&`�=E�w�|�my7~TP|E��ق_=+f񖢟~fga���(�&v��Ji��z	-Z@]-i6��S^0�s�����y����ʊz��r�xٶNA|�d�{N��!�[�ū����.�f�8�Z����F߱D��N�W�B�wq�(T�^2]���t�ɀX����Q��~j!M��K�f�!G<�4���֬y� ��M�w�$�Xۯ�Z1�����Q��aĦ��pp�2�v��u��{[ɼ#;�卋��p.��]��G��XmV
Z�|��7�v�p��,�̔��55�r\(�-��R�véB�ԭׅJ`���6����;�Xo_�ẽ�؝�?��L�|��V�|6�@�]�G�/�Tل(EΗ�8�w����g��k�i<P$�n1�:�A�'}0�������"��s���k���'�A���:H�N�,�@�n�,�����Rl�����E��s��?}�E,V�9�	����;������=^-T��5��tZ����WS�g����b�� *T�?|�9-6��h0 �4t/"vo��m�
-�_)���K�%�2�^0�Y���hupy|�\m-�⯩9n��:�y�_y:��ާ(�C�M����b����+� �T�ӈ�<Ϟ~��\6ek��i�}ǆq~�<�#� rr���P�:R���4jz�V��\g�bPe%m�0t�x�u.[������Eև����i~��	��կ6p|�3�=��Yӈ�����/�O��4�/J�o�P�r�`1<����(qo�/��5|jݰX��ѯt�`�o���Ŧ����
����,���`Ҽ{+��{�S�����0����� n�m��'@Q���:�����<Я7�DH^���WQx�ք`�M���Sfժ"8�	3K"	}���zk\���/vR��T�q�;��t�Q����;����!�K?5����$uuvf�׍�r7�e=���~�"�H���Y�L��T�������4V��,]ijM�#�2�s7�Q��O�b�6��{S�(w��mR��B������+>���%9�#�,�[})Y�(&
Z�ri�H���"����#G�{(.�Ü.��$���I)����Q?P�u1e�G�M�;]�`r���=[i��i}�������ҡ���i~�b+|O-��y� Uk©ѻ\��K���bY�W��q���"�'�v:�>�=٫��ۦ�/@�(w�DHL�OH?�j_����W�g�a�l�O������͟�-��U����а�t��A�)�r#��t��:���EX���㺇%�b�Z�N}D����w��q���$�G�T<k�5�_��24�&3�e}�9JB����0�F_ƅ�j��\W��Q(	1�-��%U�^�bOD���/J�%iT'1�G�^�.=��@�\��+$���2���,u�%�
L���msQω�yQ����V�[E+��?�8��Ur%��0�6�f�kX���(�k?c]��Z�U��aڋ��H�1g�©� ӕ擤�t
?�{���x�X�y3.H��yN�4�����3���5��w#�Kz�Zlz��k+�i����~���m+x �J(2��,j���0N�^�q�t�'%�ኙu�3�7u}/���Bu"F?V`�����؆�]?�	&:J��G�LC�`��T<UnlMA��b�L��?m%��+v��u�)�f_E�DF4�h��hw��
�'O]}�$o�4j_�TC�3a�d�2�,E01<�l���+�R��Wv���H-�@�(44q8�-RD�T����| O�+o�]d�_��覢��}f'i7�d������CX/x"T�o��Ko��6�B���a	���?L`0X��C���E!�<q�����c���&��'Tij�f�a�I�NKg���S����.?M���^��>�]�<_�7����J���Lu��L�~�P���4��a�)�@���aGggY�-�p��tf�t��`Glg���qmT)�Q��Ih���:�X̡췡xީ��C-:��C$4Ē%K�v��������ض�

�����޻�k��'�o�s��xC�9X���F	��	w9��pφ������nq���f���(��2`�	*��lu1^���\"���jy�L
DϬWںgBat�J������YA�����t�k�Wa������7ͺ$4�*���X�*`WH���	�&6�
�j�;ؐ�^˳�$R/�᥌�ő൸�:�v�ki�\O����t����"�x�[��K�:,�0�Y�z�"��\�/�w3_�9��O[����C��bz��!�al��؁����X��2!��TG�ߛ��a�z�B�������A��ߥ�[��=�s��/����1��_<�T���Aimx��R)��K|�j(�����ڌ����!�`�K���OC'�։�7ߝu)�~ht����0�.-?�3�k��A�S0��
V�ӫ�Y���j��W�z���a��r
���d*��w*�0S9x��P�N�� :�
�IvZf'��ccR��|Wj�N��Y/�z������O��8��`����xC�Ë.^�Ϳ#)'F�̗{(Y�>��+�7*~# �ڵ��n��q��ru�G�}�@��Plf�}!�awڂ����^#v b���d�W.��d5�ɬ`�	��z���zn�EI�7|�	�a;�a���o�1�R��t0��{+�Tړ�;j�z~bu=X_��6d���k�p�\��.�f�!<���A���
'�/���r��e0��:8�y9�+AM�S9�-�Gr�+�/��{�]��H���D���(^���<D��z���G�X���S	�����=Aj���?履uX�����J�ڐ�`d��5R;z�-��躻�58%{"��ۆ����R�r��y���+L�/�q�����m\��:�y���J�ӋV�t<W"��'�e��oRo\�3�:��C3(\1��d�&[����ս���*��'��m�ߗ���^��(������>̓Z�{)Z% S���}c��#�[~|�pM¯]�����u^��%�=��z�)�'��tO����N(a��<���M���ժ]�b�s�~��LCb���bd�X`������vi��N���п0AOih����+�!&3H��~`MI���t Z$x��s]e�� ��
�K|�3�Z�#�a�5ݜhq�I��k���~�T�%�ӖŪ�_���3�:���_7e00&szƪX�V�O�}i��:����d�H}p#Q;g�픉ہώ�W؎����zi��`X�kY� ^�*�ߩ����f�_q��tCx
�]��#��~	�?��_� n�ʿ��4�N�>k�5��0�����0�}���4w�/��"��_�]��1m��0�3���łX8Dm$c�4���|�����c1��׌��E�5�����&�JtDuk�bȼ}��BA � Yd�Ա�����	���U_�Y�G�v���\��͛
?��������)�+Z�Py�Wһ���j�$I��H% ���?��8�L�~1�u�������#?%M��^��c��:��ت�j����29?�����{��,��m��t'����G�����ey����G�x��/r��jR�_�����HU���Mp�;%˦|��+

Ճ�C�*����%�{��lJ��.��6��}I�[2�#2y�Lh9kC	�""��F�d�kA�x����I6^z�ޖ���U_���Z�>�tw!�A����)���	O��~��v!�����<-�'�]��$3��0�ɁHYn�����뇗��MI'�H^���NP������jOK�I5�ɸ��-
k0�'w?�ɺ&��/40��O����f�?6�]5`Xv}vJ.~U`~���:q�����7�B��.2���j�bZ�}��T���"b����K��p�32M�E�ϟ����(�Fܒgs^i6G����q<]�<1��[��v YQ������q�E�OM�M�RLM�؍�&�b/�Ǻ�JJw��W��k�,li��Y���AS ��߉����ʹ?Gס1:���㑉pB����U���G��q�����|C:N2�����[�pY��<��[�>ԥKޢ�iUtU���
G����
G�+f����Xy��i�[�VF��,C��\��bc����kO�bmQC� ��$��+�VӺ��:�*WL�*@��x�s�%/�a���AݕXi�>��lG������lQ>w��=�I���=.���-�LLʛy%V̄?���ų��B֮e�5�3��)P��Dy��Ǌa^C���U'�H4���>'�9�����ªf`�t�?Q���ߛ�z�#�@X�:�F����6�������ʕ�-tϣ�\�S\�w�e�>� �,V��f�&��{���W�ֱ��s�1�з��Exӕ3�W�,'�JEŮIa��٠]C�^�Z��i�4c@��m���$��H�9d:_��Je��U��K�z���z��ޔ�2u�# ���l�ڍV�۩�z��-�{c���0�PW8��k:*��͚-����<�E��mKk@��H�)�m�"������/�oDS�?ꋧ�<)g�O;0Lbڀ�L�!��ۑ����Tj�R����ЦO��L<n�XI̟F�F�I������2D�oK��i&���a���1�������9R�a}5.��z�zPT�*�煞�;NW�1�]e��D�G�Y�|������@k��~h/u��5z���z��|���z*~6�q���%9#��2U�7=Fܽ(#�߳R�5TI`�a��x�-��!���E�5߬)OT#�TT\3'�-w�����}�݉�-�@�W��q���N���cJ�5���(�Ŗ��|�0ήLY��uX5����XZ�\��n�� `'qv�ݝ̛%�..�7X���-o�5�s�h�Y޻�s�������K�1J7�v�}EsǮ���qN��iOQ;�������O�E|�9�8�q36�,հ��S�_�C~O����:I�۬�PX^�*۩O�M���v��ׂ�.|H��2�.���:�(�/�SJ�CJ� �]
�twK�tI#�� �H7�ݍt3�wP�������z�{�>��<�����ߩv8���\�U�Zsh��3)_�;��x�hR:�A5�V����}��[�&�����SE!u�w�s�j'Htxf��&G4�y��I�~��(1Vh��?���ѝ�U����E�frQ�~�OߛE2����?�+6�̻F��Xk��p�x��P_���:E-��4#	nX��{q��X_<8�d
�p�#MLZ�\�_�����]����F�5�w���%<��RD����cn�;uC{\7Z�>�i���S/��~C���܍|�?���U�~����-��ͦs�z�X5�%���l��z'���m�dЃ;7�=��tH�ָ)�ՠz�j�\�1��8"�t�"�b�Vq:�ߛ)2/P%����b��"U�ޚ�0���ݪ6�	Q6�&��6��;�­u�%>�H�Gk'�(7h��<oL-s�������-,�p�b�$��~ �1d7"�|ɖ5Ki>-�{^~H����ُ���V��\�щ��_��S"�t�K���_���١��1Nη�\�9$�Um&17jˆ�V���&v�6�1oTK,qŷʛ��%�*o��{Y�ENJA"s��4،J�z���+%��=̒�'���\3?�6��eH��:&�9�1H��=*��� ����|��lC㝹��(G���!8)<`�*��5L�1��6��R�R�!\E({>,)4��?�� �>�����;���u�2�]+SL7m����|"���+M��ل�e�����N.+��UQH��p��[qg}7���P88����ݤ|n��n\�.o�[A=Z$�^�i�G�y'��{(�ӭ�#ҵ�I����U��^R�^Ac[���bj�<K���V�J2H�q��㉻��:i�t�j,*N[�!�I��u�z�1�\�8d�С��`܂���bG�����q:h�a�����Ǖ�'��?,|��x�C�^,26����Q�^!��<ڗ�Y�A�}��l�)�xvc��:4�@եE�����/t�D(Xk�_�'��kYu�Z#����IsE~����l����m�qT �w0�O�`�Epxާ���O�2I?4�R���&y��f���EoY��<\��;]s"�ce s->�����?ռ�c�$�����02�Hkk85꿆wKR���+/	T�$�kd��V dsmr<<	�$��EG���׺H�� �$�})�oѧc�J�|T�D�|����>��պ2�	�M���`�b�ԇMr�(�$���e��<6��U�[H��|?"�^vp.@
�����l3D���7x�tc�^�H�0;,���kT���}�W	�:"X5��%/���N�o�/qQ���p	aJ;e��-떇`9i�rx�L(9�Տ�w�i��{�1K��W��.��:���	��'|]̬�� I������(��S%�}��5��W�UN��QX���:�EսM12 �mpJ�3���23�L�z}ſ;�*�8n���7pB�^:~([(����;\�b����~fp�c�-%�2Q��!`��t���=�]��s��z����\�wn����E)�Ȏ?@��nI�+Dp��V�ƷR\�1�f1�j��c���6���Z��hr�.DOKK�,�NY� �p��,���a��B܄���{�������}%���݋����Mu�:l�!<�����	WŃ q{�P��6�&��D���|��غ��S�|�c�m�ęn��gx �Ǘ+��o���t.�*��e��p��$.f^�v���\�.5L�B�:{��eh�1����`�3)|�/���%��	��[��)�n�g_3�l8#�$�ZX�9;&JY�=D_!��J[��`��36ml[1� ���/!�ڱ�*�3)��Gt[SDv�]
 ��k� X�I2<:�������:�}��޲����ݮY`Q�2���skh*�a��+���H�6i�:���c[�G8_7�O���~�O1f���bį~�A�H*U*�o�`�$��0A�k�g���5׾�.KD�R�|�$��R��X�W��&�$����(<'�<9ч�$�0/dd�s�'%#����I���B�sv�J��9q�?�����,�O�E��)�J��,k� ���iπ��؁7�j݉(U�̽Z�e�8��Y������+��l�,c�o̌�,p�=�X�����x�v����TB�g�P)t�2�U/l�+"���|�1����Q��	 X�2�nB���}U��{Z�J�V�_-�$��p�d��,�f�՜�S���z��g����,���,�yd��@�Lx��:����o��2!�ڸi�ɏ��--�^����aoD�,�k���M�vU��c��"	�/*�0���ԕ H��~g��v�ح������Q~ǒb���2��Nc�D{H�V%.� ����IV��У�W���ͩUP-�w�|���:*p�L��z�DzЦz�
��E��;��T��EC��@���W\�����vz�%�ї�f�_���*�()���Y��E(g,�wɯ�s�d���p���^b����xM����;lŻ�BlIs4i�?7K�N^8�o�:��ǜ���Sy��B�	F؋f�4��0�W�2�j�Q���]��hv�[�3�㖝��1x*�I��MD8��;�G�m��C���+�2�W�v�+T�U����R����6=�Q7�z؏�d��y=j��R�����l��Z��*d.k�	�Q�!t�S�� 4
����f9wS#WE
�2�X�����=۱����A��	%JP�E X:�Jcˊ�6_��.�l������D[���sr�KF������솢����X]	�|'�5���T���|��6�(����a�Zb:|]��Q�"3�0�J0UV5��.����3n �Bq�+vG���CD�s|^��\��$ t�ؕ�s��D���s3݃�2�ץ�sSrs���(�L���Ê*����ϭ���z-�o��`��J�����b�bs�q���U&�_�S��,8Lg� 5Ȉ��r,������۝e�c�s�e@hq����	���6��n��Xq���Əû�#�����#ϳ�ώ�M��T�ˉ���^�UvV�xzn����Av�#��_2�┢��*���nl�����(g��$X`>C��I��f��E�:N��Qn!�i�.Q��B��I9w ����/�A���j��%!-�LY�$�E�����.�������w];S��T���{�wS�WiZ�/�?oǈ�:����gʬ{*��D�:M���9G^)������ܛ7}�_q�.����:&��AjO��_ĸ;�OVR���&LTaַ�)$fg݌$K�z�~�
*k7��t��W������O
_��3�M�q�S���r�G�L�fNHJߜ�R�$�Ut��K�����<��Y�V�ʠ���H�8��v���O�{����:���{���N`*+%�*���7M��ܕګ����l�
6D��}X��R�_��V����%"���7�'��qjL� J�ShX����7��,!v���_o��| Vy�B=�m�ptZ���ө�~sF��H�B��L;�8��uҢ<4y���Hi��̅�8D��+��l"9�Z�6N%TO��w��y�cWR��,%��
jE�Qx��WR�����f!ϸ<���U ��q)�jش��I�=�X�ֶm�l{{��N9������7=���8
E>�O��=XX��l�X�$�Z�?�T�U�������`(2`+|����fs�n������E��%u�ّ��.��Z�>C��ӤP��m�{>��[t��ĉ�A�<�g��ҍy���8�v�_&B���p������^�.0[a�p�Ͽ�<Ю! �N� ^oֽ�iwp�./ex��+Z�֬d`�>���o(��C���*�.�L���Lx8i�r�ǂ.�
'o%.�k?���k��&�u�a5��kh�d���j]1NLH��)��5&K|�<\�{%�u���T��&�b�����5��~�)����9�w��!��dG��&k�Y���Y*���y����"��Vύ�졥L[AB���=�%~�}�:u�si��&�f�9�I�UI�B�W�C=� vY��'�u̕�¸ߦ
N�A���G��*����H�j��v��0��&7����n5�Wg������V@}�R�JsC\L̷~�r�G�7n����jn��=�I��G����v�"kЭm�գ����j�����L�^���ɩ�gq;"=.�����O2Ϻ�	U�c�RE��,����U=�SZ�߯@�b���X~�ܙ��{��]�<=����p��7�������]�B�/��H�O����,��Yց6��sX��c�G���[x�?��k�J�]T�j���n�l�[% ��V f�Nt2]a��ď"�X-&v�c�Den�z��8��UWq�[��kh����_ۂ����vXOo'-�È���U|�:�y������ѭYMUR2f<��|[fͤ��G�����M��揜;P<��).�(r�,Nˣ�BUU��$�w�䘣t���=s&�8"4e��e��3�?�~ h������F����v&R��` #�kL�p|�X�k!{[-�a"|����x�Ȓ?�1��H�P[%#d"��NҀo;�_t�uY��;�e1��<�����S��YHb�93��%՚o	��H7>Ί����M�n]��*��J�u^���6�7��Fy��V}$c*C��x:t܇?�ME��o���>���{b��jc-�Ro���b���\��1s�&
�yA\�]G��֓T������՝+I��>Q	(�:�&E������������H,A?����׆�y���1p��F^�`�ᰕ�Z�%�={b9�ԓn�뗸���0��xo�~eS��j!`@���yP֬�,>���bݤ�y��;��J-w2���9���h��k\1W?Z�	Q)�jGy:��T�Q.楌��.�M�E!�r,�av��{���,_1��9�$,�F�+l%�!銩�A|����\q�Oɲ4��D����L�WiW+����g�8�R��>��e��u��94�@X�gڄф�K�����<���M��N�e��nA@Ε%����$��?���<�"1���7A:?
�B�q*��Wu�'�ΡU+o��s|�PC�,��3uJh:Vl�;j1��d���2�=���b0�<Hl�%o�J�-W�{8=��4"M;͉UgQ�i ���U		a�W߼��brҥ\) 
�Q	� +��zа& �T��w}�b���uHB��nL��B�j�ּ�����^0��o�[���R����mL_eO�{P�5"��Q����6 O.%�r����ժ~�݂�}�R;��N+w��b�x靖�gA&0z%�s9�%ٕF���MUtՇW��Z��~�x?����/c�&V���k�;��2�@2�A�����J�Ɖ�E�G�ˤ��Ϩ��e�*� ��a	�X�ͦ�d�q/�E�C�ܰ���=| r�'�lp9~�js+��>�ڠ
b�<F��,'������
���q�jԪ�bA ���� >��3ɊS��8���0�b��"D���G�b����Z��X9׃���)�[�,�T���ܝ 2�M������O�zm�&y�صﱾ�E���}�����Ё�>,1r����O�̗�ٰ��զK�'��M��xT���!.�5n��!��q�pt����O}lL�@������pD�da�g}�HCsw�(B��i�~U�1�@J��$WƫzAB�9��I��ި�B���G���)m�Ś���z+�D����ϗʤ絢!���t|�)E~���-.��xu�1mZ��W�9�	�W��K��'$ׅ�s]�v������yN[i_qh�R��l���!��[*��q�'�"�5���!��u9Pq�b_��e���*lzpAPnf�*�<���z�b�x(�e����W��ٲx�,���}֦�^�_�ç�I=kS}jܢ�xI%��w�������
o�m>��n��n�{����%4�i�4�Æ���}�
 �X�z��z�ԍ
ZX:2�}��֠l�EzxA�H��-����/CI��<�QY�̵����>�J�>�H�}�ģU6I��`���]h[����+���|C\���Vk��Ct���Jw}/�=?�
>�� Uԃ�]^�0�)E&☴��3�b�#+k����`���F�]u�r��J4Y�/;�(�o�D��3���A���{��Ό]ߡ�q�K!��F�(��p�*�O�!b�n��\�rh�t^D�i�����%�byE�q@ofigCq��5���6�ͱw����I�^Sj.�z�!6t҄cH���0�p���f`�Q|}f�|��R�T���B�����I�<\��1�M⫮��B���5[t>DUo�V���b�4��%��!��ys#�Oɲ�d{]��΂��y��䖀D�],�����>���9��Z`1*T�`����r =��������n_ 4b2tE\]�y+@��|�BBWi�?/>k���4ŧ�$���Y����vve�Ҩ��{�����J�����jk+3]������^x���Ofm��A�����_�Y}��#J�����K=po���=1����r��x��S���3��.}7\��Zr�☧�Ԛ���H�6����}+w#Z��i�I!��-�^�+�"�b�rް��	9����V��9��A�^�^���kC����Ĕ��Ѳ�n?�hR[��'�ֶ��قhэO��Z��(]FہدR�	=M���4���7�#>n�4b;iK��/����2!�9���m������`���VD77q���p烔s*�lrs��Va�?,�|��rN��?x��7�͢V�4�����oN��N�E��$�K�}s<En<�T��?��=q�+�nJ6���������.����C��TiV��7a�Qǔ�9�4�^�%��Tg;Q1�F�5�y��`~h�[xF�ų�ҷ�'ي�!�x�`�Q=J�"�-RF�릫/���̝�+H�<����Ÿ�g]��DG�9}��4#�Z�%��L����N�q#t73�筢�vv�؏��`�?H��}�5�d8ג��m�8���$+K�Vsӓ��^�lc�V�S�|�+�����p�l�e���2�LVK�sH\�r�r/���O��%��;@m�R�!��=3�E��ko �WҐb��o��__���G��N�:��Uj�tG�'ƙ���__I=�U帔w"*I���h�������`.�uB�ė�B:%ɴ� �xƅܯ�xN�X�k	.�	G��A5
�DA�l#�C��,�m1ǭ�k�wK����k
e�RQ��e^�_�0F���+^�b��#���kq�|�� ��I�=�9�H8Ir��Z�wI*fݖ(����o��v�hZ#�=�:���:=�
�E���o�����g�K�G-BZ`Å��IW��g�H!"$��X�͵�������7s�֯#��T�D��Q^�ԫχ���oa�R	����_�p�I��/���1~hJ�����c(lCrm�i�I9C �j7� ݳ��{�`~0�ʣ��.�KRA����U[�l��[��V��Q�)�J��"ui�_"[*}ٲ���K�̣ҙ�u�'�S�PeZ��۪������P)!nI�=��=����C�cBss6�IiJ�#��MJn~�[L��ܞM��h+���;����{y�K�Oo�*��Ok�����H�~��`iU.���~�}M!�Pn����0�$���'�a��)���<v�KQqU���"΢�/��ݳg��5�n�|����|!����ns���RRytl4�Y�:ߥ��9���+���� �ą����fᑻ�:�J̸	�慯���C0Ι�����~L�:�"E�'PC��Si_$#�[�ijn�E�-~H����EDD"�4~S�w?�<[�J���.r��G�X�8̻��$�S#�ͤ��.����񡓠HȘ
�D[�����+�ޛh.q�i���`��V}�L��o���@�o��ƹ����,�j~�i�Y�,���$u�՛/����Oyo:(ܗ��'�-���{<��6�G�E���m��tc��+��qM��������8���G��VyBYtr��M��ȋ}�8�h�����H)�e��$����5-���7u��z%��Qy�EB��L�Cd-Q\���4D��<K��C���6`�7ka4��ٻ>���"�:
��N�Ӂ"�����C��1[e"��y����W%ᔜ��x�ͻ�.�}c0p5���[��a��qg\Vf�v��8�wDb�9��v.�V޵Qjܳ�
ү�+W��x�&y(����ڸ���*v�\�D����&�d5��Z�%��Z��5ʭ7�:�s�t���	9wZ����+{C�ߐ�Zh�3SZk�X��./T�����"Uc�;|PuX�?jS��>rOm��٫׮3�,%��OO�W���̶�Ry�ֲ䄍��v�!�F������I.K�m�X�QĦ���I�OG��̀�//j|�̱���I���?)c���L���l�gCJF�^��c
��c��<��[6��M������ܴ��QM5z��R�9H�|��Ǿܵ��Y�Y�E���Na���*�3���.,b6o����r��D���OÄ�7��� V��Z��)��b0�kX���Q�e�#��x�� (�m}�	ћ;�-�a2/JT�&#�{�E	���sz�zE|���^	/�1�dJ.W�{��L G�������=~\�Y��J�k��W��F�%�JR�g^&`I����t�5�}�����#����:�����jsٓ�}
�{�$3zC��s75We��S��j�	sI�	���7(uAx�Ui~�唥�H�K����c]�Az��J�O���Q՝^
�S�Z�#�Lk(�d�҃|�b5Z�QL��\�-u.��~|k��_��~�U�9��E �C�r�����t��r@4sRN�IPѰ���0�A捚�����	���.wq�kV/��i����8̒��&�׿���Sх:�$�}����n&6&�<+�Ȟ9�m��<�/��h�Ҙ�§¯^/���a惟�_뢵�s�$�!cv� ��7;\�2�7}T ���;�C���cED�I�� ڒ����&h���.%b����g�6�?����@TA{��&�`HeJ�"�f!���bJ-��K�?�%�0�U��oe��
�����w���B6Fo\��������;j��y6=��t���]��<&S������q�C�'�P�1����j+�[���ܼ�#q�ƅ��3���Ҁ����d�%E���� ;UWB+�c�x$���Ϡ�I��"f�N���HX���0�7-���WY����37$�ʐ�zގ�VЍ���S5	H}����	��8�N\�.*E5,�
$����i7=;
*u����,���ˎsxd�E�/=�,=5�/`6o2ծ ��Uʔ,��s@�$zd�'2g�cu��0��A�/V�]AO��h˹UH���	����"sfnw�h�X�$\%�ܾ]�5ǿ����1777�F�-������M���R�aB�ESglЩX����@I��w��(W�|ơ`����؜	�Vkz�L���kX�"�N`Q���R3J9�*��7g�s��fy ��ZT��n�ǘ4d����Q��*��rkW�>���WR߱�<(M5����̉S�| �=�a�{�(�^�q�� �w/���(��������)ԵZxϮ%-؃gN-�x<�g�����է�^o0q����@.L���V�R\;�
yW�G��ݷ��[��jY �?W���O���L^�ƍ�%� �aS^�]��Ғ�M�:�̻i:>2T
WK���:(�(.,O�
9�W�w'���sn~�T�bF�I	�{uS�M�ͯ�C['=-�p3P���?�U�{�N#�q��_����o�6܄�g�.
�&�H�;��d���ی�7u������N�꜈�7����"a����N,o��XE�����;��j�މ���jL\�?��Z8��j�v���o@`*d���8�m���Y����_Zd��Lq��*+��L��%Q�ZOx^1���%���4��1��0��|�zܟa��Zv�]��
5�ʊ��亨B��:g�]����<|_O]��[��Eсjz+Q+GW�K�z���ܢ#���C<��3��f���Q�m��i�׳ɚ���(���D��A��C��<_��:Kϕ�>;>/�1�3�ޒq���1bso��&�jY�|��u$Ɇ����%6�Ki,�`��ɖ	p�*bQ��OԞnD����?��nARږڪ
8f�C��/�4opmy����R�<�f�aJF���ɿm�������'Ϝ��2����~1t�A�ED������%O����6k���IAV�UB�:���`,�X�(��"���t]L"�J�@!�m��!�G��L��Ā��`O���֑�؍W�����^)/�̘|��%T����~F�\�f2�n� �c�u����B/�ÿ�#J>��4%���������t9y��r������R�A9�?λk������Px�Z�Ku��+�<�|f�UʨP-.�ؐH��VLkM��>�w�ީ��j3�y��ȑ�֌�l�dD-~�I�[�xmb�6!^k�b�\K�;LH�ƫ�2��Q�ˊ�g
����ʇ:�a`&���dzD�*����)��߂N�z	2�g#Z����C(������8e�d�-z6,�v�@W�W�������l�uoY�[��{�V��Vr�D>7o_��6��Fq���(X�A������.P���E���8�'��:��D�F��J���<�%0���o�$���]�5��g�(2�s�|�Ge����ZhM�;N~n %�$ٷD���Cd\�X����qr+JCJ�~q	^}�)VR������[@���~Fm����(��$xt�\���g�^�t���cx��I9��ZG���&�&�[в��zo�u�_�ΐ^ԍ�������Q�VLd���ilq�ǂ�^�/Hb���z��u0���8>L�~�3�^|�ҀHMj����qG��=@v�j������Ȳ))F9�F���J��__��1���Z���;�Q$?�&����an ��#t'�Si:�ZyX�;o���)Y��8!���+2�Xs��{IsZB���#���u��^�)d�Z�Z�+��~&��ǃI���73�'=��Z�� K�	��W��k������u�:G7�\�V�E�d½Ӄ�E����Д�Î�S��/09�������n3)�)�c����V��m=
�YÃ��f���P)�RtF����{-,9��\�49���o,�_�p,����Ke���ۋ�֏}�(�����+��V��`8���E�M@�+�K�0���+��&�{ڟ+rؼ��,nPܫ8��ֺ�dNfHz\e�Elo���xi�a��/c��#��1���Ϫ�F��������N��@���I��`���<O��);��݊��=��;^gz@��:6�$r؛�Z���땯�-�n+O��c<o7l�̋���S3� ��k�$}�D�W��o�U�����a���09��<�!p�n ��xu�qz��K�qU�j�S���9sտ.���e��;so������V�c6k
1���D�S�]DqA�7'�[��eݷ�N���{���L��MUKA���1&��q����n�q��*��0qVVV�c�>USNx���B��n��9XW�Q�o7M�V��4�O����M]�Z�Iܝ?
�����H�>��#������:��m�6���K����B�T6�K�j��;���@�Um~)֏�0?f�T���s���Y��g7�M���ѣn�s�b^��m!cAK�������1�1�[�wgL�;�C(�4�7#9]]8"��ʹWu[a>��Jl��u�g��#i��U�&��}�5����Q�O؏�������e�o#�k��Q'wfY��!J-'~NcY��3�j�~��ڪ�b4�N�%'d������.~p(�y�w� �����*��� ]���0`O�J<9����'���+�=�u��*7N�Bh�:�i�?�[��X���JCaN�g��s�>a���a_��.x��Є�,f��F`H��'S���.���t?6}�d�W*�U����ypK�9k���ˣ�j\����e�jO�kˢ�t���2\�Ȣ2^OR1�E�=�!���v0@s���٠��G�w�	�ww�:	c|�j��}����oF��"̢�o>�`�B�.�)�Cz�CM�I�.�2Ce�����]��x��}L/Or��W6�dď�? HWe����P�}�8�����G�� f�Ԙ�D�$Nʃ�@�N�>�PM&���i�l��L���$�[���PD	���Z�Vqx�,��$�y�{�o���������|�|��|I�:t��]=�z�N�������B��4������a�f_B�}�a�|��}S�Ѝ�JruMK�,_X��������~� ��{P-��Ik;��<�t��#���pIlH��ٛ�,
�1@h�k�G s��Z���r�r�-{ޞV�ｓ�A���r;>�(xUǎf`�ι`�:��l��̷��OD02{�f[箘*}îb����'� �ԍ��N�e
��Ѓ[�����+�!ͯHЭT�8p�R�+��-�A�V��< ������>j�f��:"���!�΁�b�A��~ٌ���ǵ����aq?[ܧ�G,����yh83���}��
5�{�/\!o?�g�9���D[hr�o"Z��􉻓~I!?�d�Gt��Hk7���$�'7��~Me��6�X澥�s�}�<f�o�BE ��5Qq�% g�����p�;Q@�� %������v������;Э8Rr�z8�B~�̱�J:��}5��\ 6�p������=C~G5]l�۶xt"P�FӚ����wjT�l���2,�mǮ<9����#Q�`=�88nGi�^bdʖʦ�H[������وW��vϝ_e� z-��k�<������]ƥ�y����V�ϒ�_sR�� �6ٟ�����@[�"��ױ����܇{�.�M�FԃB�#V\ɷNMw5�W8���密�D�(U�]'�"��H*�*HŻ�p~�O#%-������t'˳uH�6T�]��|��-7)�ֶ>i/x�$��o��'D�lC��7���A��z�ė��{�RSb�ona�#���7{�Qߚ񋹁O�A��Є�> �J�JEs+�&B(��g��M�����o���K-f/�J<�`A.S�Pe��UDl��h��U��݉Td�Jx�E�r��e��ս��O�]G�էG�fq]ZQ:�/�z��O�{ɜ�$ �4����x���쥷��!�E��ڃ`I����8w�PQS!~h1W�P}�k6���M�f����6
�5��hē�������0�p�l;�%Q���9��'q�Yセ�2�s�|{�������ђ�j1�����oz�������i�m��/�E�t+���a�*�`:��3-0�3J8��|�K�s� ]��w�ښ��!Փ��3�f��8n�t���K���Ҹ�sBA����K�wJ�C�A^o�dl�C�S���(>�A/��ln�=u���B��Z�A�k�'Z�>wca����X�k: 0ݹ�5��Vd�4m�"��{+��w��i�Bk�,~��y���7��ˑ�I��Z�`)�}K�2&�����NE~�<)9��ܡ����oU�^	��Q�5jr�H��R�n���N�D�<���G�T�*�g�����;�I��r��m
�t=�У��q���8�g�C�v����y�b�vД:�S���6�t��\��y�;�5�l��b&N�^E��\�^���^y��Q��.�5L��K�ylG�w]��M����*(3��^��R$<�%�%)�>��9����Ϡc?�M��z}Y����A��_�.��=N�+�CQ��PŮL�=0*���W ߻5b�@���0�o��Z?�b��Uu������0������돌����~�b/j`�᙮*U��!v���f�"W��Y����.�/�LΠ�7/�o}�X1��K�D���c۠�>E)���eч�L�����~�Mt�fcv�n�>�6!��>rZ���>��+�j�ow2�F����H��n*-?�JCuի{���F���~;%���MsN��`6l��Uܧ�?6�#�)I0+�[���$:�ؿ��_1^� �CW�_���N<O��|�+D
T�*BcL�-f �1�q��-�U87L���[yB]i,eO�2w�	_hk.�]2�U���L��? ����s�����q����	*��sO������b^M�Tc�~%��r�;?:α9�U-Kt}͌�^퐹�$�������?Vo��hM�f{�yitj?���@�&���@��BT��\R�yG��_1�A�SDu?C����C[oE�ׅ7� �
��ه�0�;�%�B".��H��a������!i8I��\�
��Rg�;.���Nl �}z�������� \�� ݭ�0[��W)��-E2�M���/ڸVH���)Q�f@-��\0i���3!C(����Bt�/�c�2�����H��G\/�C6���X	��o�8��.w�w�>H��tF���h?�����_/L��sTFrO ��=�j�;*���#�M��#P�Q���BO>s�ĨRI���ٴz��� ��4��{��!Ŗ>���b�\��B�hr��`����1$^�}�'��/X�.��~�@^�Xok��ߎ�:��c�&8�K��
"��=C���i��@6��?�D?w.Y�/JXQ��'���=���kj�|�%��%-�|N���8r/�̷Az�"Bs,�������Ő��1a���+>YF�٢���m�$bw��ho~�BU�2��J�g1v�g��(����d���/��4�z�����e��� �X�[����������������7���k*S�_�ꃪ\%�6�Z��y�6kw͟hy��n�`]�K�?�t�{[��\F8*�N�h�ƅ���ieF<��%#ʩ��7o����e~�-� �S��,��C"87��$��N[5~O�eF�J&�4Z�a���-"4����8*O�B��Ӹ^,����Zr�Ж���@I��R���p�x�����A��/��4=y˗5"�b�ߊ�v��:Ʉ�❠Zk&|��v�)��a�1�p\�.9��
�z����L�?���D4g� 45Dq{�{�ږ�u
�m���(���EV=��^���a���O�/ˊm3\ڜt���}���� �J�D�f7���6��5�F�6JSo,�l�#Ā��ͽ�R��o��s%|�H�$��˜�p���,Sء6i7���Gc�h��%zV�)4oG�K�b�
\x��z"��Խ�i�K�R���y;�\;�i�O�{.oC�P�b���6E���0��
�.Fp,
��QJm��!g��
�C�����b+�B�(1~ݙ:D��3��&�trton�����P�%�����%8@��pp$OKf��u�a'��i�)�J8F�s�dؚ�p�$v�x�e�*��.X�Tsn$j�_찘2�����:�&��V�q^a�����X�AW��nΚo+&�R,T��aR���`�3IGn�v�H��C)s`�0�]�����N6I�����/^2��kGe�M���8S�{ۈDP�.�[�
��}Fh��1�W��Wn�R�_��p~T�pY�LvP��R�O�-�'x�AI�[\�~u�p�;3f,oJ��KXb����KuQ��~sDh��<eV��\q/��M{7�d?!]t��aUPv��22`M�蹾sL���s��Ȑ��3[r�4n52s��ԥ^+�6Jv��#Xp�f�:˔��8 �ן�O���sn���u�j��a��6Ü�.X���A�����)�!�EHT
�jj_$��-����Z5[LG�g�3���C��v�M�`C�U[޶�u��I0�N��}ݩHrH������X�*�f%�f�N2|��AUu2'z�"C,)�Ph�������]QA��Q��q{Q����-٧����o��cY9�1<�K��o��a��0i�eZ�I��nA�,���,�F�OR��%��^y���g�+�cDj:%������ӓ�N�٭Sb#6�ʘ�t~��+��e��Vmt�rS��2{E��~M�� e�N�84���+��&���\�i%�1��8W�{Ba�X�Y�N��c�����AS�)��N�jM��U���Q��+�i���r��'%4ˈ�����:��pγ�z���3�1�b�[�I=�g�[ؗe"�g���'m��G�c���/���H��R�� ��W����|^�.[���7N����B�e���\s�62����n�n��JԚ���9e��
�
�PȂ��#�����T	�����d|��gdj�eZNϹV�,�*,�H-�7�]cܩ�<�@4M�(5~�ӓ�Xn#��=�머���U�+RWV�5a�Ϝx���3�@���l�`�^�72H�ȣ�,<���5��MjɁ߸Ȁ��E���q�r�o�t͂�V?�R����i�ʀ���f7��?%������f&�{߹Ѧ�%*�ǯu��r��� ;��'�!��
s~��dC�7��#�Ț�����ZN򘗕,}>�]�����-�·�Ks��GMtI���8ɓk�_����������FEApI�YbDi�Kr���EP��k��fU@�K��{w�v��;���|0�00�{��{�s��i�G�,�����RA:�T�Kck�Z���ݤ}���k}��q�f�黧��"���Pk��M�B���̝�@�ʅ|z��/�`֓,�KD��R�*5�?��N��[��TV�����06廄�4�8������'���5)q�=8��x&����lE�7B�sCo���yʾ��^���A�s*����Ei/Y�Pη�ÆqZ�TPzǍƥ�EE��Ճ>5��R9O�b�N�ǶkF��C��+>��f(����N]yy��y�1l8�������x9ʫ=J*ȸ|𣃐��7��8���lH��7�y���"�6V�e���U�t����w��LM{�B�y}܎��\T3� `�(]Л��*�����~?Vt���In�*o�����NV�	<���q��l��UD`�WsH��=��0{l�֊�VX)��&�7.��ho�
����rl����OxWb�F>A,)))s'���˳��Ki	��7@đZ,a�|4ɖ7k�t�qa�u��#�|B{�Ӂ�-�S����8��P�9�YBeU�nY�d�܉���������ܤ��"ٺ�tb?M��e��U�[L��n��'��Fr��0)��%��J��!:x�zq��#�����>�6,�Ը6Ze�Nz?�ey�`�(�~[Ȓu���L$m���.٢YVAЃY�
��N�Ň~ή��Z�_��v�p����n�}@O�#�f�+���tt�\zTݝӭ��e�[�QZALS�7c1�wj�	�>�x�5�C]�ͧ&eo����O���v�r�%2�Ig�x��F��>�?�S��%,J����6`��A视�5�@��,C�7e�<�u�����C�����ȍ/'�@�e��J��Í7�V���s�B�%R<m4�4�,���\q��iz�V<������U+�TCs_+I��l�48`b��.G�b0��n�b�*n��Tw	��Dw#�i���{��cL�_5y��½_Y��w;8��2ȴ��܃�|En�)��_n���@��5{��W������K]�#��L��F���
�� ��_�C�^�~�r~��xlh��X:貒������W1f�R2'�f����ƙ�@p��AƇ�a��=�yH�ז�"�g��e�-SR�^�}�X��4�P��"{oS�N@�g�����;BU���V���.�ďABw�$DakvA�k^����s{D�k�?5X�C�0m����v>��|d�m����=�ڏ����0h�@�8�Q�Z�)���zt��t��� �/�5l'!�붆we*��﯌���W�H:�Q.����w$���Xn{J��jlv[�^Ȋ�\o����<�B$[t�_�����u��<y�m{�?��*�I�8a�,u%J7D�2r�q�N�sQ�:�"��,��fH�{!�ъ�ʁ�?��������������*�~����z�ū���|�{���d4��ܲoڥ�̟+�>����|A��T S�f�����G��z�>Y"��]"e9:��0�����5������h���42�u��v�L��{�p�G<r�|[��?F��xŗ	ᤅ�r�qV}�
�m�C��C��p5D�*���uЛ(��\���Y���qg��T$�$ ӘS����>\��.C���Ĵ�#�ٺ_��ETx�4nr_�^2~[�)a���6 tUP��'2P)z�Y��F��[LXf�xUvH2�λ kg�����i���6T4�7�퐔+��M�W�R1�+�m�$ˬˎ�| A^�)��pAM���0,����1�+������р.}�mux��n޾�=�Ҵ���_��'�~^�W�4��NF�!�z���D5��U�fT����z�Ne����u�z9s�O���%���ɓ4�Z�t�X��:���Ҩi�O�\y����+_��f�`��Q}@w�@A �џ5ܖw�H��|�
��KKpx�K#��QWX%�q9�(�e�o����*����Μ���p�v2P��U,B�>�,��Ts�V��1�j��
�}�M��O*���P]�j��χ�3�[�Ο��F"]GF�����F�^�
d_J�q	>�K�2���?E<���Tn���=�D:!�izO��`hl��x���}�i@i��	r�>�z���.��Q#]�z�l1�`ي��h�C�I��ye?v�?���
�%�ns֫����L�t��xw)2\f"Z$ ��ωQ����
����-����E�1�Lwgd~:���h�.�k�uM[���バ3U6͵3��ǜzż]3�p5/�q<�K��I�|ډPW�4%g\��.x(2q���QϮ2��D�X�W�N��Â�$�EE��Y@j�g�w��>��hDGKtv�'��ɯr��_)�̯V�S�����K��U�8���ir�/�]F4��]�~�d��K�H+��`��h�!D��s
S�U�I�I��7�����A�#<�����ƃ�nZ>�Y��&�S�)��G��oz%�$��%���-�)l����y!�#N���R��wH��T<	7��_�y_�I?�����{3�U_%%�9ޅ�J\i@�(v� n�ձο�\>�����E#�Θ�Y�I\\N�~D�`����s,�����G��*	�ٖ��t ��BWy��be�o;sO��n��)j���V�����s/����x�d���s<��m�#����Qj��1��P4�P$�֙���<+�bY�:)���l�ϡ���*��*��lp['�65%�T�$�jwt�IѤ��*&
�C�S�V��SG�zSq���.<���W;�S(�J�=vj������0�9i#���6g����gca� ]��I�}O���k�)YO��j/�,:ճ��XD�X�=����-�~�f�"$	�C��H���T��N
�Z��K{��9��W����ɥ�.<yޯȖ�#�k'D$-xm��������k'�(٨#<�rB�yd���+��k]��đ������Y7���|�TK���vLG�&�m���fL!�G�P^g�$S_�Y�"�~�Ih7w�@y���R���Rj���6�+E�T��k�bF�U��$^��.Õ@�X�����UH�zz>7�l���׌h`B��X)����V>&|ݍ	�����[C�ި���n�����X�
����]�y��hd�D����_�={t9�H�䃀|ư��g�N#��J0�3������"L"1�~K�e�y�tkr4�����sՓ�r8����(\]a�m�"C�E�i�%�������B�~���,o1���ݎ�O7Sx�G�IsP�~��hM�Qf>�Y���ǘ�L�b0q{c����ml^����"X$�ҽr��J����K�ng��]*7���A�L	b�a�le�B�Ȋ�U\�q�UG��*�L4e+馟#�B����ɽ��5G"m�Q����=��}o�j�h���'Nx�GsU��MjWz������{�)HۯE�*�ޓ���=���")ٷ|�
8�I{����.t�ś�&���C��M���py�>�qá�r�V���/�*���<o7L���7��m��y��V�]U��Qҽ���d���l�T/�(��N9��O�y[Kf�\�z�w�tcx�v���Nt^H7��.�E�P���?��7��TH9�j��ͬ���Iq����Ϲ�,�$�'��B��*��:��c�(_|�;�˪>�.A�ìK��#L��\�%�������<�����닑v���������L���A&�:��΍�dP���Nk�Uj�DG���Z��.�F��s�.�V*F�r������W�a�/7�8��s���(G���8H5?��~64�1�Q��d7��"���	�D�	������hUte�p+m�h��
~%qu
*̄RQ���V!�筍u\֯}糤1����Må��RV���3���f���ƃ�нNN��i�#Jו���G	�hph�>���+��VȦ��H(���}��X�a��9�ѓ��O��������E��]� � ~�7�lK�7W�zu�7N�f�}v\8׌����������F�`����&T�2&�p_c�x�Ѱ�(i�)��ax^���,����g���iٿ}M�Y�$�p�{���f���̏�Cyn$�SG�&EAvɚ\��4P�Ҹ����&K'��v�9����~<��z��>�/[4OeF��T� ϗײ��6��L9�M[0Li9��d{7Zٷ���z%.�N�Z>E�;�]<O/�j���mf{�� gM�y9J私R�hc7�71C�>��m�q���x~�}��[d���Af@!��9��Ra1�Y�i��N"��b���	��1BېJ���״gp��"�ăQGe-�{��U��"��.KuEV�2�J�}]jV��	d�9T�v��R�����{��C9C?4�J���3�UHߕ�L�9�w�{�1̥&щ�.g���w���,�3���\�&0�H5�JY��"�d�H�n�w��sI��Ky4D��cE�Hys~�q$����7��y�ˌRx��~�i�`L5	U��{�xx����<]yi���Q��-�'y����4���_��K�t���[|X7������|5:�>�����Wz��BOݛ�4J�6S��)�ƈ+������
��N��I��D��O�ֵ��r��+���|����#����=�� ��6��Tb�"�?�����A �� �� #�A�Z�;�(�&ц����h���6�m~��l�!��I�m#,B������Č�Kg�*/���?!J��0%��<�	l8��c�_8Ǟ�xr�4
�j�t<��^_+i���6_�Y�$���:y�������B���7���`Sj8�@E1���k�KA�����絥���B)����k���iʷ��?&�\pȚ	ȧ�t���S0���,.�p)�O���� O٘Q��5�`Ҡ�'m8,)�σ��f��=�.�r���J_���?4��8) �,r�Oۀh<�+Qy��f�]���g̚�HOW�6�r���؟ �v��}�����v��T��꺋.G������:l3Pĥ	�4��OSBކ��c$A���7��@</�Ѥ�S�#Ď���}�-�W�m�B��Ro�������\�i�{�eC'��J��Qγ7��᳿%��?? �x.���y�����'��F�2�Zt)���|+�R"�
����eR�<p�i��=@�B�s��2l�$ip��s�0��.`��>0J�pq����9�O��}FQAÈ*&�R��}��gCZ�]�`�}�4l������5�R�v�t��}?^ta�2�	:՟������Pm�'�:��<!_�qͯ�M�E�0&g��!v`���Q{�p��[š����~it�L��r��k	8�5��H�����B�)����
��W����o;
��RV�|�S1͘h�$��5Fg`�]kv&�6�>,�G�������}�ͷ���	
!������Ȁ�g��K� ��(��:U	�֕qV0�А]k�-c���� Oa]� ��G�&����6�Cha����$z�L����G(���Q�x����\�V��]]�g��6����I��8��Ef�u2��=�[�!r��7���EX#�9����:��C]J7��9�)%��;���n�M�#*�	�Y���_��Yk��+J��#��ͽ<�"�5���U����ph'!*;P迗���C)����6�{ �����"�H&_V?[�/{@Y���# ;�O+Y�_l��9�DX	���c��G�ׄ�oڀ =�UI���� ��>x[K@Z��B�����#�ML�\4���E�Ň�s�OZ����Y��Ҳ���iF�}E>�
�E
���Hh��|��7�_h����B2�;?��/�dX�e�`���V�?�|���V�qe\�����Z�Tq��Q����h��� �`�%�W�9��J��#"h!�I�bF�͘�U��DK�j�5�1�0Rh,�7��F�^�r#F)�]T��5�9@��b5�̫{a�E�7'<�[Se�}�����^��u�M��%����v�*o�@̶��"ZN����.S#�r)�ј�'��"�J��.���
x ����A���*=L®gDQ���������p��i��|��_�c�M6~�������@�Ǜ�i#�)��nQ@*w������T詁Y;�K�	�/\�&�
f^g���~�����j��ݒ�$�R�|zPKY��6@�T��mBǐaY�}����}���#�.{ʦ����U�ͅ{n�4����5�>��Zu�ؚ����ah����@x"蘾2���M)�3�j06�^c7J���h�����NW^G4.��px���mZ`��4��/���e���: �W[���5^-��&����.�i[�Vq��>;��X����a��(3��0�x%���slW�U���+��)�ۀ)xA�#�9�z�!+����%@��𹠹��@����2H��v4](ò�1����)��Se�E?{|
�ꥹ��f���ۘo���o�%Z����T�9a�����է��/�i�R�1�|�x��J��t*�B#���:��*�?�vy�����|KUV�{�c� ᕩݳf���ҔU-2����Mj���ڳ�\��9�$���,�i�m<d<����C�����5����Ї����=���6�j>z˖���̺�FYN�@B*����#u��G��mƕ��P�C!aY��m.� ���h�)*
��wp/���
��q=�,�1���6���*$��Ya_�X|��H����$S�|!��<pJ�x~���@�i���N�ٳL*x��Dm	���2.��o
C4����$	���?<�h��K�8�WW1�w'�zd�"w5_��yI�-��e+���<˯��1QC@6���(S��>�I�O�r1lu`%'B I�����d��<ݴ�s��,�7{��شvϹ�o���N�J��5�{̗y�ڋ�,ާ����=��e��nll�~�b^u�����Q�1�ʳ�欋|��b�w��dB&�����Q�0u"���(]�/�j�nO����D:��|� ���c0ߙ��]�4&���)��E_�d#u݉�J`j���c�&��8���gʭ��Z���wEqp�'&���i̮	�E�D�OE/�O֧���=܃��TW��=��qML���bk-���ڼ
 u�7�-�x$Sbe$�v0�=�-�%�Zy�b��6�
�^H�Q�@�2��,�����Ҫ�؁��-�<D�ua/>�ҁ����&6���= �D�����0	��\.S�Z��[�/ϼ�V�_H��r��������< M��0D� �(�.���@��,&��������"��n�N1$oK�>1x#��?+Yy����e~�����Ǌ��(��4s�Sr���͜��Ӫ��=�Ȭ��Hќuy����*j����;���.���P�`pv`M��뚈t��(F�ٍJgUqGU��$򬏮�uvGVW��ή5�Jk��'���"�����un�^}����Jc将�yƵ�K���]E�4�֭��dP��O�s}Պwyq���D ��?�T� >q�/��tѶ3/�d-5y���j��$MO������W�����ϼ�8��|Z��"���a���aL�l,��0h<���Y���S�r���n��Pu#^����pJ��͂N�LK���W��TcBX"����gA�����ڍ~z�PE�_�w�]��|��ĿƇ�<�EVWImH�R��^U)���#ba�O�a4�Z������[�Lꌛ�Ä�"�.
7��Jޕ!M0������v���_�1��`��%�.�tsь����JD���Ki鴔#|�e�`F�N�� �_`ɇ<�KC�b��x�]6Y�Ҏ﵂�7XL���&�%~j�bh�%��z^I�k�����/�R�r�G�2�/dO�˻�)'0�ї�M/zM0g�c%��*db�ݮ��xz/����T0Ͱ:�5�o<jID�:)��s��Q�9Жw�iG]Y�#��������V?�7�G�QISwYN�fw�^��vM���2͉M"����W���n��4��]�i_.L�0e��)���x+������Z�k�4����︘��F��q�Y�D��|�jU�ܙ��}�en��-�SUT�~�E��8�|��ê�a�IL)�V�G�롴��h�oo4V�,�mr}Lˡߕ�^��r���ѭ�[L2�l����>N(I7�:�%���T�,��<?b5�b�Z£x5?�]�7����'8�U�V�XY󔥰��y�U��r�~9�pޙ�� ��m>�{BJ�e�g�R�F����.Q�P�R�ѧ�p{,��Be_�����Z$>b�;Q^�>�|���EV�el�kn���u&@P�l�q�z��I�<��˰$4�C%�(�M�ȣ��|M~۬�Q#�۩oHTc����'����p�}�?DxRW0�/H>�rO��"�Ns��(��4�C���&y,���yb��\����#I.����+5=���[�&H�9��6�0�V(�p��k�Q�ӌ����x��Q-��q۴�a	`�/�?Ӱ��\^#����B܍�H|�Z�H��;>���@.k_ͧe$<�&�@^�[���-��v=�����b	Q$!���|ֿ�^��|�zy�o-_�>Nׂw'�����<2%�]�1���0���/%sa�I��i��1��a��V���Hy�U�:�?�I�n(.7M�DuX��
'�匱y���H�d�fţ�!�f�gz[7����OP6Z������j�V��o�ax�s{�'`�����,��#����z���K��np�Y<�otc�����o�Y���X45*��5�i*?x�?r\,$D���� jݗ>��L������k)л���`��:���Z�/�<��w�i<�]���o��ç����݋�n������W�0�7���J��a�r��֎\Ƽ�t.��]�&o����~�_Wv���ǹ��3k�u���'���[+1��/8�5����;f���3��rצ��t墯�e�M���0=���^��g��,]��|R^�_��- Kn��<�p�J��w��~��)���J�p9��;����ͰNò[qc#�f��ݶ���r�E�"[��8�s�ݡ�GߝmS4=r�7͎�_�D��߂��5�0ʒ3����1߶�8ƕ��j�]{�XJ��4�Až%��.�p����l\ؔ([WɄ���{��K���D�S���ˎ��+�-��L��B��g��������#��9�F9C!����L��H��f=���Q���_)ݫ��Ej�������|\�/1���gg�S����F��{C$��8���X�)��GVZi�8{��G�.�?9V��Sh~��,��=��X�y��	��p����>MIS�-��f���)��k'v��&RH��b�H�n�3�wH�ؘ�����2��?̛]r��}M�+��W��A�B�����c���*e~/]�j�Χ��j#N� W�xY��j�z=�����$`�u��?1:^b��XŻa�Y8����U�㛹|�uqu64��/�����@�D(�V)���Lm�:]�%�=���	ʚ��Wɡ�~��O�r���$_��g��g�O�dab�m!Vx�-	��<�R�
}9@��ٮP�JN����p����}K��ߎ6<�:=�SrH_�_~(B�ԩ��P�yOd�:pn؋�X��]�Pk2���H��8�d������i2y�h^__��Q�[�L��������t���CA�8� �����
��L�ت�)9��������yW���?>/��AD�$��Hjڋhm�L���P��x�i4
2Z��Mz�/'��;4)[�XH�7wz�믮�Zk�����KF�g�VARfv�&�jB������]�z[�'V?�@�Q���v	��d~�K��T���M�PE�xX`����f�w�|�4˾G�ڮٙ:>���b�rؙ&*ܱ�U�-�}�/�������J�"��T&/�_��U@�6羑�菅��S�%ʝ`Fl����&ս䪇.���+垷M}7 �\�jlT�O'áM�[T�OW�}Y���?��)��"d���0�~sҷ˱�����D����rq�y��	BP�=��V�Ջ�p���#��ҤuMQi����?aV�5���$�{���Ԏ|�L�#^�Ӆ�7����ﾹ'5{��/�V��"r�c�'MRF{�Q�D_���
L�6{�R���Xy"��>��4���`<�F�������"�<ǰs�LyOkT��ʹ<�h�~�VA/�O!y5���ONɜ�T):-���ڟ�.ᾐ�&`�NP�7V�0p��<�5�$��Ĺ1S�G#3l�z�'����;�D�Q���[Y"\�w��R�b�b�:�Gh��{�V��Q��N�bV��ȉ�3 d�h��s�ڭ)g>DS�.2_�uQ��F�_��������'�A����@�o����"o�qى͊�'�7��?�nuz����������_��-�G���'���\l.��J�稿�:�ΰ�m�f�z�1� �[��g�-o�r���B�U�q� �؉�nߢ��r���B��u~ُs�����(ܛ6��-*y�q��Ӽ\��Vp}G�!��L������eO�`_��i�&I�	��/��\�8���)�s���">�'ɂ}�W���h2ɣ����O������^9n$R���R��jkL��h��a�۬,�y�?�J�E�0��y�k�Z��gfb��ͮ����꘿>"T��ԯj���Y����8&kt��J�2�T��ttyD�PQ_��)�*�\�?�G1+��V ��{n�N_�6����)�+�b?�p_��)��1�z�蓰����3�)b��Qe������0V��@����o.4�6ȥ��u�"w��f%��jPP�RO9~?} 7g����ym�^�
ѼSVE��b�y���^;�e:�S�������B���W����U��[�_(b��ܔ��o/�3:��]W�u�PZ���5�Qk�lz{�t���J�!�-6�� ��ڂ���׸Fѐ9r`�����x�1�s�Q2"B�l� r��Z�u�����P!3}�M��ܧXʜF�	��=�-����X(c�v�|^�2�_YtH�)�Q���uib��|)*�Q�c�fS�⠀Z��'�Ȱ�Åc�֦�f�p�� {!��xŎ��-Hq��c1nR�����#_�����p�� �pt�k���o�஑���(a\%1��Q������,ǁ��_��Կ$�Ȕ���(g��1f�R�B�J��3т�R'����0s�p[���{�A���|}����ւe !�������w[�k��f�6r���|�VV;�#R�^��r5�;�2�T�P�F��{,^+��\;��7�%MG�66�Y����N�eu����I���O��>/;�e�8ࢯs$(v��l�/�\��w��J�����Y�F�n�D�&��[4��2W��|��j�k���&���/=�,	��LH���GVY�i�w_���ӌ��_�ik�Gxd9�|�т���Dc���d��W�\�Pg_��wCq��NRj7��w'$���}׸#�iC鵳z�h#�Z0ĶZ�׺؅�f2��#9�1�T���j�`Fw~cz?��ʋ�R�͹�p�؆��c"j:벞���I��o�1�3�k����;�Vt�=����~�����ɤ��iS���Uυ�m��?iX�OL�Ba�H��J�ee���U�1���Qt�K��� ��������^��Q�^���q3XD��ܥK��Mu��*	��FkL�0��e���X��i`*Z�>���c`1nc8�;�(怾e��U���+aR�Hzۺ!�VA��|�C�c����G��1�R}�<2wUb̮�9��=-9�]W�7QIVv~��<�Iv���⏹�y�	�X��d�QY�!��mׯ�x(�k�{t��\��|�����nz[�V�12�QH����s7,ͬ�G���#��cҰ��F΄�=J��G�� �k �HaY"@�8��\���@�^���%<@|�ºkf@9��,C}$��?�l3��������~���bgOu�r�iTk\�"�,��W�;T��Q�Bde�Q,����%J��e2q5W���kးr�
�v=,�����DV�}�~��� ��n�ST�*O�u9.�썌p<�2�9���ҹ��-އ�r����Dr9}�p'k�͚S�\N�~��4q{�Š���G�a�9��k������y�y+k�MɆ�`�~���-̹�'p6b�6��j�_<�s ��H+Z�6"p&7&���_V�>y�I��R)�*�&X���u�b|��� �����ċJIH�}Yx $N`_r��\Vb#'+���el� ���<��4DA��.i󰮍���?41���㒟�.ƕ�{TG�1�8^R���J@[v����Ð�3�����6��^q�el�q��!FåC�f�÷h���%Thr�����Z�aÑ3xӚ<���s�oP0�bmr\�A�Gx�O+؜�U;����f���Mg��z2+:9;�E�#���ڑuwޞ364q����T#-����Q?�i��Tۈ��v��^�����C�I���!%>{�.�WD~�6zTi`!�)��]������ _`'C�7���Q����/9���|q��y�X'�V���k�������"�� ��-5�G�~��X�(:�M�<�O�:�x\#Z�T�!%#��guy�� >S�^5d�3ʅbSH��v��~\�C��8�	?gA���y�:��OKuï1����@��i��!`c�=�޿ѩ����T������F���G��_>���0�^�
��q���]2���(��O0�����$2@^�"� p�6�R��ߺ���u
��B9�.�%�k`�
�V��J�ak�U�3_h�����S��f�K�;���Fq�&��jo�8�dY�$9Dbk��=)���m����5�0j:S��t]�$�`�\�-�۬GGwpcW��x���O;ET��>�����ޥL��dLO�8|��U������/t�zL�_� �^�;Y�݉i�=-[q|TJ:!l��,�]�#��#0J/0���x�t�#:����mUꥈ	��K���X�i7�oj������I�C��� ��$?�۷�z8+� ~!��;ZcA7�����3�>h'�M���^�Ҙ�MVn@�TYɞP�䀒��]�a	�7=���e�����Z�W���+A�þ�d����V=���a�T������/l_GS\�g.�`
��;Y�eMy�#��+�<`�$
�f&M_X��Y�<��=��x��	�ܓ�-H��A���}�l�~�&��:H������[w��9�������(;�"���v� h`t��g��9�E������s���,��(#I����CbߡWw����{�v��`V_�9
����2��������i��,�]�)�=:'E�V*ݬ��N��d��	$̓9��=��J<{�}�����[H�E���
#�ǉo6��B���E���[���������7#sɥ1\2߮�Ϣ���l��(�v�/�J�B�]��:��v�g~砋Z�O�2>	7��nz�!�"��V_�P6`3y�֫�+Zqf֖m�_d�I�z<h���x7��	�(b?�_b�?���
?���� �CMv��"��S����y���X-�a��-hۧ�db��}�������}@���[bNm��nf�;R�\��Z��V�5��yr�=�v��R�ʲ�W�V�����0K��l�00�Oh4=��Т�i�����NRUZ;�t��{��٨ݚ�?߁����m��
ľ��9�J���g�ɟa��vXABƔ+��.Es �����A�+���{6ԃg}{t�;�5>�tƃ_����Qj�,t�8�U�ϫ�d#�)պ��Ҭ���"�ñ�5�ouDm�CqR��,I�_�
̪2]h�Awg�	X�1p�p�̖n�:�OǷ��>r�����]�]2�ג���V)�g�$�,m��Ͳ���o �EJ�FU;�dn������Q`&��9�b��g��3�k	G���hqE��v���,��=\���v4^<�Qd�����h�RP�|�aH�T��ݖī�h�9H�PAwqC�����|Y<�HH���X��W`>FZW�?]��g����Z���M�`�Be�O�|nR�&����v�`l�����<�{|�(���:�c9Vƶ-T��M%Q����ʳ];R��3����R	�����{��F��.����P������AX��[�
}A3E �ś�'ب���-\;�+��;�z�)�|_�p�����y��Q)�=���G�d��#�k��]!�M��O�,�Zұx��^-|��%���㩢���/<��+���~���-��)U�;%r��� �.Ox����"�s�"�C4	�"���L0����q�"��t�7�$��WZ��a��X�Kv�Nν��z������W¯��X����lX:&2j���]h���m`5��r��L���Ny��gLg��7 ��V
��J���C�v�_&xYA�I@����M"5����z�ʳ�,)�j��mP��zeI����|��y�v�~�9�Wt�MClk��MҘ	I��/���8!�����Tmk9K�5{ނ�6!����c�g�7��%���Oȑ`���U����L%�ja��� �	nd:t[�y ]��u��!��l��4� �m&	�B6c��$q��h� F����������\k�V(R���'�*Ç?v������g-,\o!��Am��O�xkx��aCc���O���W���_�S8� Ŵ���/�۫>jh�9���8W���QQ�{~�|s��f�k��L\oLչ�.8�@�L|�E�X�H(A���#�"'mYf�t`�"y���E�/��{�ޘ}fb�3y?(55s�o�Fs3�G��}�Ӎ���w�+����[� �?�וWg	��WS�n�v�FF�N�ө{)����`
Z���u���1 ��`�3+��^qH遺g���}\ u���6���`�Z�������T��>>�݇7WЯk�ި�z��(ӂl�M�u���\�,�0���m�a%/�=�Տ��4�ϣN9�8���l����M�Pʷ�0��:� kw�o")82gnQ �Y�(}���G��5������dټ,��R��-Ņ�U��C��!�N�m�s�����n��i��v�*ڄ�O����E�ca�l�m��cE�l�<���I�z
���O�뺥u=m;� 35N-3�����h�Z�!�6��}z�͌,M�º�_(�h�w�'7��b�����;�<��9��g�<�3Ӟvk�÷"I��6Y�*���r��OEE��]���G<:���|F�z�!��Fd�A��顸�t��W�hxxKM�h�\4���Ek�1/���: �^�.���G�-A{b�0;��z@d��lǣ�{�������UhZ�*딖�"��'����|$�c��ٝ��n�-�) De�e�����E�Ćj�^����Ey��.#R��d�����Y%��h?�	�gc0x��>�pCe��+&@1&z�s�1��h�:�d����Db��r&_Ä�x)Jd�U��Z"fj�~�%'��w��?%If��x����)t2���t�=t��ͳ�Ӹ��8��b�1���F��ᏞEf���ۛ/��tj"o�?�K
�_�f�	D�v�F�X���g�Jw�lu�������e���=\�n����i�'�ͯZZ��<�\��[	�[�p9���ERv��u�'��<���85f�_~��T��Ԑqy�<�l�u�t�)!��g0��v�aI^���k��:*�� =���e���ujR$H�s���J	��PЦ���-h�	J�%��?
�r�`�\�G�0�x��&c����F�1�uE���u�q�Һe���)r�`�v/�0=�Ѩk�t����8n�7��\TSHI��s�qH�~h�+�ׁ���{Ƭ��d��3c�1:F2.A��曫��2�&F�קx
��7(���|Վ_���n;	�Ƚ#q�wF���/�+��T=n�ٳ�hf����4��O��x�bݫ�&�<M�c�[��<���_��;-�qI�,i�`H\������v[oyo�f�� �(�d��|�t�q�i������I�R��M��iW�]jI0�o�(�W�֞��9� ��`�LG+��[h�EC�����f��3��4BZ?$�K�HVk^fDIN��h��#��e�Zs�.|���5����9��_º>�˒���y���>����:���`ɀB('�V{�˲�����[]�B�;���$���U�rL��Rl��65c�h����k��>@IݛMR;����]��0"���=���m��~`W��pH�R[��QP�`QɢJM�U�]l�Db!4v��-����Wr�S��m�$�u�}2���
�ş~F�(k�IH���yO�����@�6��>M��o����k1�]��`�9��_RBB��@��[A�"����B��G�����,���ѥY�Ƣ��WTAmeq@E,��]����J��U�a�7�7��YM��%� ka6X�:cQxoÃ}?�wk���U���1׼6�TH�X���{�8]�}��!�6��f���$6�b�S��l��X}�|��Y����;�G�B��LB����/�(��?ݣ�)� �7]S���Px7*�zĞ�[�OeOS��	|A2����S��Ϙ���
e���Ƴn+�l�rAE>@޻V�Q�V��b��=��QQz����Gt�%	L����C�v`z����piy��{"C���+�+��c��Y�x�'���3����4.[:X�W g�=ӴΑ�v�?L}eT���6"��t�Jw#�ݍ�ݍ�t�t#�t�4Hw��0t�������2�k1��g�+�)�W��D����"N"�<��7MP��:�k��o�=�Di��걫����e����4��(.K�xQS�&|�
.wý�� ��7>��/�S����)�c�G��}ɹ�����堆��Ai�����u�˰6sPQ�G2�Q������c)��<����B��p0�.~�?䑿jޞ���6ܠh��}��a�Wz���w�<^{�q|�A���E���S��B����]ޮl�F'ގ�+��>mR��?����Y��S�m��X��sr��̲ؚyL�\c�\@�L������;P��dE�#Ā;{�QMg�[�JV�B��^{_���u���1�����P��C6)?���E����2�.�:�='q����#�a�a���X���������[�r���R9	�"n��nk9�!���$��U�7j9�l�)�5���.]Wj�G]��C�q�ӕk<�`\�lU���砵N�$���ͺ2ck˴�꘨�@��<��1�,[��oF�o����m��'�x]�
�"��q�O��p����h}�B��j�w!��#=ii�0���-}�Rr�����5�;hL��p�ξ�N����S�0}.��:��<�c�r~Z��5���d����	��l��i��u��J=�{;ͷ[Q�/��U��Yt<������
���v[�f.�U�������5ςR>倭-\�xi�:̻�����*6�TEpj�0�ǽ��C�ݷ�i�Rr%��cv,����L¦��d��Ee�E�֫��4/.��N�1�u���kM}М|v8�aqF��I^r]:@�kv�EO�}��.g�����`u=͐G[gzV�=�-2J�Pr��$<��)U���զ+9�~��D��ܤ�l����="�__�\�3�8BG���п�ld�i��#� }nF)ʦ-�[�A�=KcY4�S������V]�D�?�!�͊��K�ܭ�͂�z0����sy26�W~����+[�(W&mjw W�"N;�m���x�{��]D2���_\w՗ Az�rwr���I}Vu�w�/	��q����]��N��P�b
7~[aĕ~^z�q �EA�N����3�]QC��p��fW�LwT�g�Iղ��8�}��8�(<<�Be�^�I2�M�>pg�L
CA�+�G��<r���=h��V�q�9� ~$_N�֝IV��
Q/!�*��[o �l/[��_P������Y�oHUkm?��5��ک��g�*]h��N�-�B\ �L)�Afn�e/������?2: $otG?y7u�	#\��>y�j/�0FX��yP)�<ΪaCt��n��7��+Bꎹ%]�� |esM��i��P��`�kE3�\J��Z��������j/���֠�|�-q+�g�Z��A�˒U%}㴇��t����O^>�+�W�(�olu��F^I/�~����i>b�X�
t�N��\��E^�+h��<+tg��K2o`��l`��O��pb��!W�nZ���"��8Oi�a~�y�gT�6m����@��<qQ	���O�R�f�j�ϔ4;n�S0F�Q1i����Z��m�����d��P���-��[�l�F[��!0n=ݳ(�_����8��l��$9�vo���*1�G�ׁ�E^ׂQ�B�-��ca"o)��<�H�:\�����$��ꖖH!��:�(2�9i>�<k>�n,A�#��]�(՛����8��q#˓�(d���|�;�|m�������kYF5m��m��t�F����~RS{��ţ�M��!�5*��L~$�w����F�gZ����̢P��ܪj
���,������}��9r�f(mM�1��~>rZ�6~M�����S7��ѭ4L�x�14�Wp�9�h�B�Q�ICS�>C~f��橔1���b�ܿF��3m-������jMGF[WE��N�Cs|��i�j�Rc��D$��sĦ���x)�PJGT�^ ��~�1.�Jj�~Wѳp$P����s�z�m�+m^�o�����T�&�����#0fE	�`lTJR��g��oK�u^�.檟�g̰�-b�V��}Xɤ��.��+���iQI ��x>�mz.z<�B�i�R	�+�i�f�}�����E�
�%��C�����oѧ�';W�.!«*�퓨?�?4��%� ��:M�C�m�FGg�M�S`x�����am�]���_��Qh|oZ�3 C|��!v:��y��߾?nP�}��-G`�W|����v��֙F��8����1�W��%lv���>���Wr��Y�x�͖�?t迕�y�A�z��ڌ�v�@9K��N���z^&��B�Q^�ڧy�(������K��z���i�ѯ/R�b�H�����<���,�W�����c��:���Sp0�ꋯ��/�
�}�X�03�@ۚ��*�Av�>�ᕉ�>Nͭ���h[���� ���lK]lQ� �?�VcE���MM�����/��fL��i��&���ga%	^Zp�0�g�00���|��(���҉�50�8[+鈆� /�?�0�5�����|1 g�,���av?��a>�W�"�$���:�!D��'˦��rI�'��UE�*T�ǿ�F�bn,�����!�� Y����]�y
�$YN@U��Ǭ�$ZqS�
n�%�%�80?��1=Ò_�����-j�G-ܟe��Ļ��$�W�ܧP��PE���!נ���Z��=,�-TIs��#��ˠ�CS���TP����>�~#s�c�iYk3^³G�TV>�]�3�[7�b�����P�9(�ۺO�U�t?�` a�mtB`��s��[�Z���>�� ۻ�&�Ay�(�Aﲡׯ��C��f{�%��~<0�(";V��*t����Ocb$f
'=����0 ���,��#��>����l�_�4�>^��h]���yC9X��d�m�6.� q�N�K�\E�r�t/�s�j�.��������Kg�����/a��앉fRʫ���u����ds�k.
0���y�T����ܹ�a:��'�|b���g��*�*i�r�xI�UyH|�S��S	����݆��V���YT��)k�����sᵙ3��|`��M����;�ss����)���[�(��&�7(����b�J�49�݆	I��Q��^	���<�{/�ȓ�vC�za�3��1��|<;�]�ؓUv�����[�g��RX�(8����^��P�w���f�����'z|��u�tͅZ%:��w	R����`.O�|ך/vb��
�^'�o�W{�;5�͟�Zk��f�%mr�}�T�F�2��wA(�k���=�����O}@����񇣩�";�<�����^S%_O�*�Kʿ��f�g���CY�p�\�y\�'*�1�"UȉkU�(��a3�=��y��#���l�@_��@�Q�FL	.�C�����a7���ϙ��_s��`�LU��\��Z�YZSV@����E�cNHRR�UXKJ~���}',�ۊeg��z,��71-�%����s�[N;?ݦ�FX��-�_-џ�[97m�`��nx��m�8�}.~��)�3����U2]�h�%j�oW�<,-�Q�W��,���.N�9!�v�74v����~>�������痢�Ip)��L�ͮgc���[��B�PR�fG��z�̆�)�K�"�����#�d���7h�`��:��[>P��w[~���%}�1;��F�'�7���ظ��
,�.>u�٧J��K��]]\B��-*-����6���%o�v��FL>d�����$4 �"l�|!��1����G�Cg�÷�	���^�v��Gc�0�S˔_m1��yZ:=5���:�!Z}ޞ��v}�̈��G�"���7-P�o!)(F�V�/����y��tj���P��P������M�����-���ٳTK{��'2G`��&��M�V�/�<���
����sK�J9Tmև���5�S,���N�� �Ϣ�O♼a�S5�"�-�!��"���;^�u��O|4;���u]\L�Y}�,�w�as�������0��OQ�
���C!W���}M�z@ֽ�]:U��ޔ�ʷ��"$u�+�;X�1ko��z9�Y�o
�F
��9V���7��?��՞�-O�I��'�'k�h�R'n��?�DU+�(�!m�N��3�=i��l��:�"��sj�l�*�K�ٺF������Ҥ��X���鹐�I�l�7����9�_�3�1�'i��(��N�m������-���6Z2���sB4 �b��X�N��~�k,��Ϝ�z����D��<*W����/���wO�����t9[�5��	��y=�q)F2���V�w �����:�&�}:�Q��a�N̷�@�#i��.���]�d:�/��y��ǐ�ۊ��`��\�'��a��?�<LG�2��oc��?�Aۍ/S��ЭdҠ�+t@ض{�k�r�*�F��j5��3��;$;�r�&ƃ���q9ʁ	y�%D'�#޸���SO1�8��K�vS�Nm9�*�,��K'��`�_=�3Q�Ay o�v���=�y��T\��<e'O<��M��m� ��u�;ݭ�O���h�GGjzT��]��4YTw~¶��s��)�g�L�/.���;����e���G��6��F���8�Y,��U��nC���R۠�iR2���W�Q�&�M�O[�EsJt�Q�m��
�.K l��5gF�ì�V(���rJrL�����2l�ԥꂄ-6j�P�v+�Rj���R7~���{��;<�AP��qS�۩~C�Y]Qd�J��\o|ԫ�Z�l��y�������Nc�~���*��r���#G��-���\B��(�G��V�\m[�
����V#�v-Ao�]梹��b`߯�c��ѣ��i9�N!/�p���n���^U����� 	�e\o�
��.SX�,
Pm=��&�I ��LO�tn����9-�$����x�q�-���|��O^���D�����C4���Bf�È��72�1���F����S.r,	N'����*^�gۛ�nP�o֪��3���D���sgaT��I���"q����R���J��6vh�R����;�� ��4�`���D�L2�o
&��xa�s�]��M[��*O,��	'�G6Vv�CAڞr�Ï�xms��n�>|��|r��Oe�ߣ��ݹ��:�z�N$}�z���\�ҏ7��
�I�N�~�Q����9��>�� ��F��F��m��O�: W(�ˬ����T2x��z`='VeRNh��d�CSO(�E�D�6i6����>	�m��w8���"�@�s�xe�?��������;�fü�Cy�Ps��R(���D��~�#S	�|����+�����jO-'�ئQ��߫$=v�E��;��������ZW�?ލ���n���OY�?�i��}�n������E�'��n��~�\=��k�l�2wP��f�l�1���--����y�4�,4������K���y�}�eAL�1n�8Ʉ���]%��I����	������>��o���U��fGIU�_�aݐ ��4�F6{��iҚ$��F��� w��_���6����l�������1.�S�\��D�z�[�H@LB�Ҝ�ٴ�4���h��)�Co�˫7/@���SFV�]cNb�$}ca�H���~|h�e��e�����-<x0F�K�2���Q�G���պ��p�+�k�X]��G�1x3��q�`�_������uĕ�c�Z"����8`�� �"=S�6�iKn��P5Vp�4e{��Iɨ�ڬ��Ek_�ф/\o9���>��YI@"�����'eIy�EW��/��kys��x]��V���"�������7�U�6k�A�I�e��W������h��Zd(���y��1�������ԬH��A���+��?�p p�r	���w�)/���au�&%k�ݝ��u{ځ|��ѻ&_~��"Wp�F 9CoJ6��݁�J�^+�)��\3��;��g3��:��e��C$bғ�d����b`��	E��A�ēo��
�ww��é���g^kw��@\%�.gl�)�H�EuۍB�%*����BI�_"|�Q�>��t�`bkXN���{,�Y�Fޞ�b�L�#`ɬ�FyB1{/F��[��դ��|)�+�IA��� &�a�Ӧb;⧯L�"�x�{�~g,e�G�u��ײ�ck@��� tBy)_hrj����L&�gS:�����"��aP9�JC�C��y������Qİ��H��q��&��Լ�@	�9]��v����S�O��eq�C�R�f��3���i��=f���~:hEkJ^� �E(��I��'���¥���QD�v ��E{	!UD�㫝�n��Hg�fB��� � �[��W��&�f^�i1�	��Q���$ʷ1��pm�rS�;%����p����o��㽶,5*��Ë��*M(�N<ϪC�eN���f߳�M�w-���S�'Y��X����B��޸�Z�M���<P����c���Fq�hj�����q�����l��	���e/B�c�lg�������k���;ƜG�3��oT�r�����F�V�_"BN�	�O��h�T����*c������b����ފ��DRUܭ����4x�;����mEa��4�����Έ�	�B�G����.>k���f����RS���L0�ʔ}�&?�~kurN6����b���09�0>_�X�F�u���
���T^5��
Gݙ�xq���|I*@F"^���[������n�^NnO�|�����}���uԦ?mr��F�����0|wt��n^s)vO�o�E�)�>l<;���m/��ȷ��.�����l��|�:|x�7ٖS+i�*�؂2+�d,2K`�5����$e�!Ƿv��֥5�?�6J��̯[���I��Sɜ���t��������b�;5�oLK��	R��ګ&��oc�h`l��Q�J���H�D�"S�J�ǻ=�E��-�SGJ�n�E�B�aA
���F��̕�%����>�\�����U��B
|KQM��IH��hn��c��+ESd}�5Z��G���I2FH��E@��Ӭ�͐�TK�߫fA��y�D-2g����g��6'g˕Я�!2�ddE�E%�KZ�ږ��D2w��V�B��7��צ쓯�d��ݛq���Joz�RN��� 0�7�OG�kP��s��ĵ��b�H#,���B	k;$�R��Z��F�L�%Z�ExP>�~G�[�K�7�%%���5	ɧWՋL�!Au��.��4�J	db��aS۵�秹�����e�TgӮJ0�5��d�* �[����^��t� U'�`��eA�Ux�e9Њ��	[s��!�/���%y?���7u���5��Z�~�����O|�P7B�JF�T�'��Sc�թ՝3�2��<�܈.WfĲ���)��+ %��ϣ��*���t %��fr��^��Q�o��ɱO�N��O%^��hdZ{��f��@�S�&���oٻ2��p�n%�"D�r{>9��#x�׷�Di�����l�^���JK5�+W�Ey��'�����z�bo��5�Чݧ��r��O�H',���������Q���S�>|�A�f�ι�U}r�56��'j��R��#�FϞC Q&�����h�`{�y/S��D�N�4���$�7��%��߿tիQO�A^�����g�޲�\}B5n0)��D&�>��ų�G� ��/����^�����W��z��k]í"��1gKܿB�ڿ�~/�7��0)�0�XT#0�f�󳈱�q�B4��]�e2�A��S:�Y:�m<O'��<8�Qb���P'����3mD3���Z�&� V�y^אָ[��A�o�A�2����9��FȦܘK���is�R�39G��/���j8؀gu�:.h�6�/���<�u�x�XSu��QZ.��� VF3�w
1
/Y����W������8Vv2�.-�{��\�������tG�i�I�/�`U'x¢�M�熇�ɇ�ʕ)K����,\\�n�MM�i/�s8_��@h�VZDt'�5*����SI�4Rh(��������4_��q��������O�jd�y�K�|@��V�I1��=��N�kh%[���9I��'��V)�)W�����¡���7^�9�P�t"1�e#F3�2��[��v�]ޏT�_7% ��5"���ws�{a%La�	�.6���9;F��6ib<]��Lܮ�YK��ڊ*��u?�� ֕P\�=������p��I��pI?^Գ<��O�*�u?�?�kB������&�f���nf�b�6ΰΘP�"f��v�GQUqޤ��Y||��s��2|)���b�x�8W��t^�3��5S4���N�ԩ��/�T�mK�[��U
��P����5���_��c2�eDHtOȪ��O9S'���Պs��^&��N7�M/�P�5���]��s��\��~v��q�j�$�tVUM|F}E�b<Z��OSX0�:`g�G3��ct�H�f�V�դ�@�������C>��[����Ê*�b�E=���Vu���R��l�V��[���$��3�X�3���8NE6�5bLNP�m^cl橥X8�3�_P��ס���`�b��|?7(�.�_��@y�8(�@y</�*.�R����j�����sY���ƳF��k�WNJ&��B��ע�p��O�������nDko�7�����46N�a���*�f����������ZjȈ�Α#{��Ğ�%�A�gh�Pc_��`�R�(�hC�������x_PkQ·���a�	�U)T�9�|$BI@��#9���3}���Lf�̦{����d���O3��ؘz;dZ�w �f�inm��j*���>^n(��k8Sa��%t��|�4����U�?��� @|�	�*+r.X˭I�ֺ*v�^��)��|�|�t��]5�4o�do�����@��'��㜫Z�h$�{��ؾ��[�q}�7:s��d6�yh=ļ�F��0H�u������:����ɋ���N��ٌ�ڜ*��M�(���RW��� �׿��1���������tlwa�.O�?�W�;���/�ݶ��،��68\���j�b�7C�)�܊�u���Q0ߠ9�rk���i��c����}R?t��zY�G9>�!�����ׂ�$N�R��������[�y�t�3>ᇀ��
q\Lw��%�x�Ϡ�ٸ��K@m��H9][s�����n�vZCF{U~���Q#E%�X��]�Q��d���P��a�tP���JER��Ӯ��U�̙H�j��+�� �<J�DHH=�����G>`��a��>��9��Kȥ��>�R"�O�����=]��b�E��sW-�^G��ݕ���ɅG	��`X{=O��=�}�ml�7{���?(2K�'i�_~$W��w{Br�}�r�q3�2�EG�)�;���}���P��(s�)����7�d��>F֤�i:���6�4�]�=n��#Y���u+���a�̧���t�a��l2�N|r��k�rbl���WϹ��O&7.o�j��G�?�kh�{�J�0G�@���P&u|�Y)�	Duom�7;��cv|��o�C	���Qk�L�t�V��21�r�}6	OQ [+~Yd����'��K��`��C��Jn�ښ�띣���u'B�,��N��/_�-3���8����|�&�33�W2�vY"v:q$��&_|��N��-�"s��I�<
�B���	��I����1�waA��f��`�)�Q���2n�p�j^����-����Ȋe�$.�ʝj�!#d4(���a�ޗ���.-�=�g����ZNO�F����r#{x�̧8�����	�}Q�2`�f��&;�eL?"�A���T��ܼ���BV����y	d}{�0��I��oڇNO4�^�[5�ĝ������#�k��m��Be��V���0�I���N����Mm��8�-Y�;۹��M>�g��2�v��A��*�+$�)���E�|��K�g�&S��v7�K_,���˘���#�V��(���a�jg���#Z�? �sb$�w�B�MG~����چE}z�H��,A�p��Z)�}�l��m�`F26��,
D�M��K�^����\���$�c������F���8�G�g�`yS�s�����m����y_��9 3���E�+�A�[�Z��WS�D� �{��u�n�b>��'G�'�gN�M���섇'� �3_�:�m�= <�X�_��7�^�^����������J�	���x(�|��a��|��ր����ň���V�O��|a,Ob�j�+�T�-��J��;_���,ۯ�؞zvҘ���/Γ��w~������������xȐܳ���h��o�~%��v�B ^�T4f�����y��,��LuҮ��@�]�ܮ�xfF�ח�;S���=&W����zr�-���O&;w���z��%���Ū)�� O��7�������vlJa���EJ]�Ni����"���F�j>��_�R�ּ��6�� ?RK�AK��%���.�~@b���ꪅ��i=�O���rgS_X��A���/mH�H�f�,��]SG2�J{�	�I��+��B,�[<���>��ɔX�?�#�.f�\�Ҡ�&uZ6g�G�A�J��6F�����j�I'�7i����f��v���?P�tP��r�MQ��9'$PX P�t!l�l�o�rɳD��vh[�Xa����j�o��j�0�Q�D��E��}ʿ)�<P1;x���53?�Dإ�\$��*����I輞�sVD�GT/�O3!]-����lT�$��w�jY�S�.Q�m��5.4�=;��>;��+�(�z��-D<���V�ʩ�FX*^
�}��*����\$6�!t���u(g�Y,��i_2��HvW�~�TJЁ����T���TE{o3sY���s�3o�jݡ�ljq�2t����������}5��|:�5@� ����������c&����^�
��uͨ�tR��@�"���ۅn��<��t�����k��
���2��՚�b���i��
}�R�|���L������9-�0H��9e�g�	�0������4�^AJ�,�*�����2#�аJ�DDKs���*�/?��:Vb.u�劦�,�Z"9��w�_����]+5�z����g-d�Ĕʙ��^������_� �w��`v�O�<M�;��s�u����N?�׷�FDxo�)���L�0;l�@����,�-���gR�gd����F�ʏ��@�s�Npg�<���A�a��������P�������
�CKDk�I��L�����sS�K���L=�}����U�?��ѹq��\��zߜF|����͈W֡�F�U�3)�&��x��c���>�u�0q���o\�*�i��/�B�0}�Z��e���+L����ٜ��&`q��hǴ�ƃ�i_��Y����}�;T�-j�-<2�q���*���=3j�7I�va��m:Ů�g�w�eϓD��⠐���Z<���S�i�
��8��^��qH0�Ι���Q<�(Y�Bzq���Bn{���|����L�՛��噆��]|׊0�>{Hҵӭ�������[,mi��"Vj���B5n-��\+|�\�.���?%��jG^j�ZD��r�#J��2$�<r	-���M��P�g.����ٱ}��t�����"5���W��zȆ�MwoII~dGMH�6�3ޮb�4.�m�뵏W�z��BB�~[���kA���.䐼�~���r#�I�R
�����"WA&�@��69��ڛ�)_�Rۏ�L>��B��H���L������N$Wd&�_?NP��m�Q�'�DW�D�z��7������@pa{+0���y��F����;\���u+L勑)��jV������S(p�|O�<���9����(OPY��	;4=<�ؙ�I����z����ʶ�>L���C�V?:�n��T2�j%.�.��/ؔ��r��M���8۠�*���>�|��r`��@��P��
�ൌg�E�3��٦,#�������,�2��b��z��0��yw�Q%S,�����W�DT���
Sx�؜��Ջ�8������Rd�6�>�a_y�RJ�����r%�eHFE�ЭA�
��u��
z�jzJ���B�/�٨�r�qO���s}�;�R�1���Kz6z�>TC���؞{i�3�=:� :��]c[��-@O�yr�TI"����T٫���[��	���u"�D�`���y, �����
��O��'Y�K�x��h���K��Cn�ov�ĉ��������b</I�r��@�%ɖ���&� ��pDij&BAl�
��8Z�b��.ޏ�F������R�@�#��O'�#�U�b��VX(��rZ��,w�G|(k�^���	��:�BS����{_@�̣����`���͹�\	g���gq���b����*m;T18lt�dU�9��y�o�(;Ue����x"��.��R�r���D��y)/�V�X��=k� ���_�M���3d��9�{M�P��8�od�,�j���iKo¦oĆ*�P��v�T��M��b	���BE�_قy�i�Dj\������g%��4�es\���!$��G|�Kw�
�dPt�(m���оα!I���5�?�ў&��0��jE�V�D����W�<񱤱��%Y��M˕�_N%5���g�hf��d���d��k>܁�gܸD��N��Y<,5����]2���W����-}.� SD�?�Ѡ�ƉP�qF1�A.�z}�[1���xg{������R����֏ 0y��|���2=\��
�|f_��ll�D徥U|������(`D��5H��	j�Nnj�1À��-�}<����|M�&~R�H��-��u�p "��.�Y�_�ޡ�&�$��x��6������mD)-���L��_���ₓw/�X�}x�YC�'���4��,�(خ������͑��X��"�>�ҵ4Pq{(����i���$7<���8�������qfr��uP�<��@B����Ei8�0�����~1���,�QC*���������vO-�Xd��fS7cq ���ly{.���bkF�g!�<��(Y�fW�=256�j����U�	�'��G�x�J�FJ{?�| �0��u��>Z�"S��AJ��TT�ｎX��_&����"���g@:�.X��B��`q��`��
~H9_��f������~(rDC��s%ĩ�{{w��U��$��J��L�o�#���m�{���鵘	��@�گT��ތ���W����'rPp�u.�L-�'A*�6�|l�翃��H�\ߗ�r77E�AE�W}w�'uJk��I��p�B-��ө3�xC(pӂ뿠F���D�nJ��Z��Л.�dߞ�*9�߿�����yo�.��\�~c�k�7B���9��UACm�'X�9=��i��ߛ�0��g�P���0��)q�k.�D�=�����`��؁�Wو�|}�癦�DO܆
S2��~i��v8a�-�?�.���ٛe`"~�GU�(O�b�k�P��k+N	2�����{�%�Fb]��b'��;�A�'MVJ��⻻8�?:��x7��G۳���T�;��K=Õ��q��$�?3�q�?�a��x�b)��9���(��̦~���!����c��u�:q��&�j:�0�|q����5L�B�G�<jx^ĭ!�ݙVZ�����e�BZ�K�$�A���ŵ�u�_)��J�_s��4��!�P����n/қ]*Nq��̺��P�ݧ��Qq�5�M�W�Y�Jq�fS��~6#~ Xf
����pZ��+��,�t������k�UkY�G���d�Sj��ofz�E� ��kn ��r]��]V�����L�k�n�"̪�!S��%�3M�\w�s�9���.w�ü ^�;��L��$��$������3A����J�G�����1�S���N�AQ+WiRTi-i&�em2�4����N��c���"����:h���s�?�d'¿w�U�o��
�����/�[���@(5Ta�~v����`3b`�~��KbX�~�l�(�
(Z��ō6
�$���P��Ę�JI���*4�3���Lt{f9�������4T���?�=��S�y�z
}Y!��YS�פ��Vs��OFe��o��i��jr��ܿX�I�l�;��{�&Mqy\�A�'y�AjI�Q���7��{,���m#5���\/1�����,~
	o�I��f5o�_&�#���^����~��|�,J����7��c�C���o���|(��P�I�@�4Ȇ�z��d�+3gq��N\��D�hDvc�]�6Ԑ�db�&�P^��\���q;�+���[�F$���'f�-gb���
����
�(��6�x�h��<9�.�:F�EAO�xŧ���v�Y��ְ�=o-h��	�Pu�fL+�J��(�I
1�?ҝe>@�Px ��IL*p�=s�:��:\��7����QV~�"ʰ�9��T_
Y�N�ڙ������<˳�b'<�i�̀���NF��H��_H��8�ހ�p:h� �Z���:vFB��l7�6��[<��E���0Lʪ���]�iRTE�^���ʂ��Ol��Q���,��&��g<"'ᵍ�{:���1���3��
-iW���T7g@=h���hmW�	)?#���Xz��m�ja]X��8�L��^PP�F�L��ҙv��dTp'�'b�Y9��F�'�FJBGB����r�"���J����8'Iu�B�iN ���L~R���_Jʡ'#��p�����V>�1-�{1�{%q�I5��k>�F�(������3a�u{dW�檁���b��+6靐����Z���w�E�� 	.�������ʵ�)|t��7?VX��Mi�5�g�+P���cT�S� ��j}�M�����G��E��LI�%mvs�	,w�?}����?������� }b��s��p���3S+B�,��-����B��Y�&�T����[���G�֡0z��MiN��N�m�#��پfJ���.�E�y�~O-E3���$�%*�!}����N���p��N'Kz4�N{^��4L7��-�ŭ�N߮��c�ؘ]�&��2�tPv��׉-�%� +H�����៼~�S�4�RK!^_���P��2�>�Q{f&2;��rwF����L���SPK�8�&=�w����zX�'[�w׬���7�X�L����2f>���|X�x���f��~W�8�ۓ�A7�"7�A��r$A����,��r5l1�!�)�ȍL�SF��g�x��S�\[�$�t�?a�}�)^�׏��)�f�m�[��~Ň�ӄE�lE����
7c��WI23Q#C���/
G2@؟/ka�|�>y��.�?x<W����,
���a6�%�6��C��EU�kc�)����p�~��dRT��b��=y�p�U�3��.
��o�l������QVCLFH��F����]�� %�����XT<�X%�~������:	ߴ|�9t��1��g������$}�� ʵ8��'���J�;1QO�4�^[�x�a�(	>���%+��J���8ͱʐm�e�����ªqҺ���f����L�� ɔ��l�f7��"��J�dަ��j��,�d�ko�	i�X%�}��ĕ�,}��,V��\�E�)�Ew�rM֭�~I�晘�-:7��9E�:����!�t0� �zl�0�qdx���/�3˹Қ�-+�7QH&��a��aD7(�_�-�����)Q�/��JB�氩7�2ؾ0�bg�p����"	��W�G�އ�jo�g���b:�0Q�VO�aL�i4�WU�6���(� �]��3K���S��S��w�$E��<��i�y�P���G�G�#������������r�����E�-s�_�Y8��y} 'AL��*����NG�v*����7[�C��~����v��:��<�b�������Nư�7�Zaھ��'������u]��~�_�3o�;H���^�J��}�C�)J-@�O&r��صL��$i�6V�Ҫ����%�R��5#�5��<�9�������,m���ـ XW���(���[�,�OoO��,���u\9�����E�P�����ig����eho{/�	��UiHK�jP�G����^#��"�*��l�Ga��X��������|ti�:C��[:�!�:V��M�)E��׶gѢ���Q򈻦��&��]	m������O0�'(��={m�r���Ed2���������I�����tUG2n3��wq#{�PX��@%�n�j"���X�+�Һ�����d������]⳯��g�f#f��fg*��n^�8�~|�9�K+�Q��-���&G��O��.�����V(���u~Ga�T���'�(8���ߊ;�/<]pQFI��0�d�P.%��n�����j����� C�twH����  ]2��HIK� ����C�{��?�s�=����Z��o�yb~�9��{[<��k����6�E�RA���?�����J�F�Y46��Z��&��F8����uY0VÇ�ɶ�����w sh� ��L����^��|zl��3�^o��dM�r�o�е�~�ŕJ�B��W�:��/����N��IX�s���W��n��H���\��QAY�"{N�a�K���tLptֺ=����"�AZ${I��ߐ���#��g}��5�]TΤ�x������k��#���] �[�v��2
Y9���|�}8O�� 6�ú��Tz�jε�L^�b>���U���*3��"@Ч������Hdx��s]fD+f�o��6�����({�:W
̄
]�e��u�{V��\����~�Ι���!�\�M�:�~yX���=e�$E�p��u�0��	�r�B�b;��5��f��*R����	�]�埰֧Y䪯_ݦ����'5l�ɩ�s/�̭F���,}�/3կg�Xu����W*�?�=�����W�����/�߫C=ɜ��U{K���O1���:c�^�D���Hm98T4��
X��|�mO�O��:T	�p�C���p5�B�y�<_��-�8��Z�o(�6�2Zb�I��m��[�55�/��#Ъ�y'��!|�r�^��P��P�Q)��j$��;c�^�E�r8z(F=� 7����M��s�<X���f`�P/��!Sm����/�y��'Z�(���U)IL���m�K9�Zb�(|���2��õ��]P�Km�N��� �D�@���QA\w��-;�f��^�y3b7rXx�a����dW��]��[��uT���НC������6*Z��S��k��v;6]Z36ŞJ��� "�b�D��>Y5N�6HI.5|f�#�!p�� I�y�%܈���"7F�ߞ�IO�u�
 �J����O(���̻�@���i�)�:-����9��&i3�	b�����*M��U�ͻcV�}BlM_n��u���H&�U���B#��H%U���_#'�Lo:vż��>���,xg ���/q�??��c�ꀱy~��e��0���2����H�[���'e�ϓ�X>��D��`n���sŴa�Nx�49�@�g`���[ ��/�����t�c�Vn7����阮6z`�)�/^6[�5�vE��BHA�.܃5L;,j����⇂ݻ�>��}1�2p��������R� b�H�
v/���лᲗkȨh����ἇ�}��Az�cS�$�t��k�˩�kUSխ�F��U�P��>fT��K9/P�k�Y����F��_CH�#���?v���w�SfC�hQ(|T5�;�v\�P�#��@mfl�Kl�4��z(�)�i�а���-=�hW�0U �d��� %$!�X"	��|\�r���ϋ�@�7n4*z�d
-�����x<ߨT�s������ךS�?��d?\�ͼ�S:�'�vv[��9q}7Q��[�����+��qk̆�`)�Z^��<�;�����Xi�]��~Y�Ha+�w��P1������xl��bg��;عp�kO�)�|�dܳ��;t"��\_�nt�}џA��.�c|�xd%�g`�V�#䒼o�}2A3|������:�,���d��y!�����2��&Y���D��j�$�.�;�t~X7�eQ�ɂ���~[�ab�+ 嫞H�hq���#Y��6G5w���rr;�ل�[��O��#9��l�;��q^7#�tl`�X��V����rc�cD
a���L?��:S����J��?�T#����%���J���V(�&�q{8���$�ձ�g�s��y���{�A9���	{b�I�����(^;�7Wlz.
���T��h�_���3|m�^Q�n����z0��uG�H�};��y_���FTc���w[H͆'��@C���p�,��;�3��d&M�bW��w�'S��'g?��1$���Ұc���4iHүr}���{<����@��3r��6���T��?�ꏧ�`ާy�5:Vv��>HX������w���f�Ic�%��[e$�Ҳ�wR��WWjC[��y���׸Ks�$W.� T=#ud~a�*B��Y����w���e����2������o�ݟt�stG�d+�H+$o߶g��:����hCӆ(3t���Ҕ���L��u�G��'�׻�j��%��gfr���K�`�$D�t7EG�X�pΉ~��cյeCq�4Q��I̱!���_w����-#��m��Dp�c�K ��v���ҦVia7�ǭ��ۼ�p�(��H��G!�Yq5N�_�����M4�hEj�G~�0-М��Kq�*����}��?����x��7t�6���B���:kFDr�gGCη.-����S����
g���uq�W�T>����";��������?*/)MO_�:�$o@���D�3J���%��O�:�Nc�᤬��x�:`A}#=��`)U/�/K���ӟ[��ۮC_�'�G���D]�|�m�PSx$��c��典_:DY�%�:�Ҏ\�Mʡ�0�"��J�rX��
D������o��d�SCj@wF*���8G���eњM ����3��{w������!�Su�2��/��R -��� &��R�Hִb��z��s��V��N�JŔCt\w8�P���l*hͿ�4���R�Ss�����ѺY���q�4���u�7�j?/��=��߆&�,�v�訴�Y砅mr?�)4l��~�p��L��XՎ�ɜ(w�&��$��	_���l���O6@�<�̦O��|C��F�rӷ��F7�Q�~�+N��?�V3*��Nl%���I�x�,ɍ����_�x�x�w�&�&���I��\02��y�ir��
����޳�]n0����TAr��K�Fr[6�{9�/����`"�e�3�ber�=�zΩ���.�)i��:�w~p�� ���H�UcS�ŷ7{�SSw$h���V��FN����k}9�	��&~����\�-�l��YG6�d��hL|�I;V�t��cƳ��fR&��P�:�U� !D��37K��7+]^*�"v������������GR2�~���
n��#b�OBe�]VY��Y�5s���r���tv��9��/^���K�k��n�OT�U�.�a�EJ��7�;+=;���	 S&X�3���A��*QTٞ�I� �0��+Kv߱>&sV^ˇ=�o������ ̜�:����@7]�N�X�VG�G���%cqK*t���B1m�u��1a:Q����sHe�������q���?wÕ|7��IwN�~h`˚���h�������ۄ�Ar�Q�rw�7E<u�r��ݦ\�_��<�
N�u�	��ͻ�I�*_��9�O�60O��	�!����9ɍ������g�}�dK���W�E�mdd��hk�=Kx��fa�I7ien��=p��թ��� ��~E|��w6���Ş�X���؃C4����A�&�1��6R����L#y4���K����ǰ^���2 �\8���h,9GI4چ�����w��'��>/^2��.�:�O?0+�Z[(Ѯ�a Q���F�c��↬$���)���F\I�2^��|�k�j�C��aܷK� >�BH��p�r'S"�Gm�'�y�q�lr2�-#֊>���B떐�"�B�Y��! ���$Ӻ�f����0?(��p#��wk�0�q���)�B�>�r`����	�/J�'�Q�PEb��;���@ HV@����:��-/�����d��!>���v2GI^���͇uH�$��g�.{6{���1ظE�"��2}��Cs�������#��ł���L�T�C���U6�m�.i��1>�P�ld�2\���f�#�#�9y<�K�0G�e��ew-������N3�#~ɧ�����UѾQ�l0�� ��*��1V�ݪtP�U�c��F���u|3��)����0.�%�՗���q� '�D��V�?ĉ��)����T�5w��ͮjr��a'���-GP��ǣ�G�����g�+�9����mԨ�{�&��2�CI���5#  Mѕ+ڿ����@��F�ϲ�VMj8,X:#�Ь�O��M�["@��HT}�����u�X+���_)p�j� �E!�X�nY���[`.B��,Oo�Re�QB��}�կi�;�6�dFE]���ܽ2�q�Uޔ*��M��#߉�8��@��|:^�@�T��ξd�Uh�!WJ\����<����
'@��Z��L��V��pR8N3vWL�F<��9�5l�+�m@�F��e�A�v�D�v�%_5���V�S�������4?XzV�n�S��̀����Ul�Uu۬�$�����>���n��{E�u���EB�rv��tLu�k;}�QV�.]1�G8!�u��5(���[Ϧ`��Jn�@[��T
�!%3�Q���r�ߊ�vQA;�tfC����o�'�'��.V,Q��>b�����hڀK5缾C��i�	F�J���4�yv�K<��$�ק{�S�Xԛ�͗Q|t�آ?��!]��骢ӊB�*N%9@L췈�3���������T\����t��wu�,���Rc�;���'\C{l�t_y���t?YD�(�P.��R�p��l�~V7ň���LQqPK�F�6Uj�^�3?�6M��&n����/�ɵ"?�|$�ܻ~��p�뢋!�kQ�������ј�����ê5x��]C	G��v�5Y����oDNrd6�]�E����y��X��B�0qRx�
zgC��GSV=����������� ���$k7@��\����c������X��Z��i	l�0��y�%&��:��82�E�����ԃ{�ԏ�y�78$�E�F���Lơ�Цw�؍ Q<]�p'��ҝ�2F��t���f��~��L��*ϢW�����x�_�vD&$kP��M740f̣�ԿS�ޖ���I�g��;�^*��~T����f��_ČW.���C������͖��ڱa�Ʈ��*��.�����"T�8�.�M���>�#���ĵb"��}ݯZ񆇴�y�^� �`��(*��4��U�Ɛ��O�w�n���n�qVU/-��_���[�c������.O�}p��pkz��hx�4Q�#�BT�;��n����B�,�������b���7H��*/N,��E>�hۏސ$ܠD-�\zඇ!��S�t������~�ԢrL��zFۣ��/�R-�S����#�fb�JY�O����ƅ`��).6��U %5:�{ʟz��N �h��Uצ�?�	p��_���d.�8>�"��Ȉ` 9vZD�Mc~�{��DI�u֚V�@��8�nBbK���h�4��E\��s�9��R�h�|�AX!טއ�\jM�Z�Zu�ب2�M7_Gy�ܕj���H�kV �����uϊ�n�0OS�r�G�U|�U�+���$&T]���8n�0�"�O[-8wy;Z23����ܻ��8`'�2����M��錍-~��0h���w{7U�9q����n*��[�޼��hhq^ltν皻N�����)�Y�I1���Q����|�t�������!�P�u��*��a������0?�q��$
E���k*��nb�	�&1�s��>����=��U�k�eO�}�,�4t�xq����ƭ�A���IM���p��:��
ױ�ri�_�����"��'د�t��_�[�1e������#�S �a��v536{A�hi$���F>c�����>�����������{Һ���Ax��V8���kA��I�t�Y���
w��?x�������7�tZW��'+?���5I��l��e��e�`D.��o� ���A�	۲�Q�Gy)$�^��k��cl�_�(�Y����_]U��h�2G�L{�o4S���'��<�g�:����Y�`>F�������̙�7���G�sj	8m��;F�3C�nHe�6�mOZ����H�ׯ�����h��~L��0�TY>A� �R��m��U1�n�[�E��E&,��N:K����i;��3��<����(�#��)gR�@t����[f!�猂���r�����>����u*�dD���P& ����dٝ�GN $�|��ܾsdԞS�$J�E4�pxi�S�"���j��\��6[�6O˱�M�����7T�c�e�ʍ�Ez���/q��~XT����p��/�ڢ���uU[�˓t��X��qS����R�d��ٸ�H�kF'ʁ̌G���jL}����}�#����
v'��T~���$R�k(��Tz�h.����O[;�����f�K�$B+�m��S�G�vSjV��i�y�=O�x+1A��᫞eF��.uK�k��+#��G�9��I�$��0F���Ņ����HF<cU�e�/�1ʵ��<�.n���|-j���U���8	z1��p!�����f>��W��5���8�4o����j�nR������B�h\��b�	�������'�c�7��^��5ٛ(����dF)��<���W���ts"*�)�T���k~�2%&�U��=n��Y˺�����!�9�ecϸ!�a�x��J���U;׳�M�~��m~q2뒿�* ��$K�KI���l��Q<����q�<��L��<e��.�i���,����|��N�}�6e�������)���~�-���,�4a)&u�ī����uɅ.����=��o���y�!���Z��;7��o_�
�*��l+0�JA�YV�}}��|�n�x/����N�����OhY.��C�"peÂψg_({~����e��%}&@�W��N~�/�E�O�Qe� ���u?��ܳ���3��b�+�݇�ყ�,���_�nx�]�n�-�8�&�
(�3���E��-�&Y��waI,����BoF^ĊM݀��F<.<ac6c8�]X~�|E�-��/�̻�[�aLrw�S��7�����@!q$ʼQ�F�Z�5�k.G��T=�#6���]PJw��@����2غbu�obN�<:��F��2�ۯ��ڪ�>B��(x�z2BJǑ?)���7+������(d�v�s�i'��XӋ��R��q�GG���K�
B��s�%_k˸��փ�J�	rы�8g#T$w���gW��j�4��S"W��Ǯ^��hќ��2���\�Cbv��D����y?���;�	��]Ҋ����>���JDؠ�
��JOZ��|��.����j�p9j����!3�X��~ɱ����]:�x�;�Y�V��쵟d�����QW�|��d���4Z���0���|����� ���<D_�t�l�}y�Љ�;���<'A�hDZ�>�d��(�<�usuF���*I��;�>���yzSx��an�2�D�,��[�O�(�/��-x���"J��8�P	ռ>�N�O�j!���T�<�^����i�����@r���hF2�=-�ۣY�l�S��0�Iy�eF���*�ଆ��k�Μ�9\>��jC+� 9�Kh�\����G��6��#o����NT���q��b�un4d��ha�l��\�$0*.�Ƀ&�Br���ĞA3��ڋh�o��MxJ��C�z��Mu\H5�F�0���`���ˠm�;��[�����)��jÎ�,��D�kX�X#�U����-\%�Z��AS�q�f�CW����A�g!�_b�r����'�OK��+��Q��ѝ�����[]�}39�Z���wv��ً�'?4[b�G�Q�^g�s��Z��~�5��i������$ӊ8@.w#�P�g���9��Ql�Y9%n,��U-��eU�Or�7�S�5N��d�yP*��5q@�9��"�Y���Y��8բ1����5��.A,P��LY��}�R{�w!�[���)�F$�k���7s�v�H�2�r��0�x��S|Cr���E�i�O����tTb-�Ӵw�pJ��Ŭ����������(�K�F���;P��i��?��N'h˾�ה���ɣ��C���r�H��(8Kĳ���G�Y�K�<�J�O�jd�%�@T���a�6��c�>1��}G�o�asS��dhţ%�Q�[�c�]F�_ŵ��l�x����{0����p-P�y⍼�\���c�xP��\���ʍ�;���$��/v�U��LGv�SL����9P�]u9��̔S=���L�.��l�?u�)���Ԥ1bű��V��mK�i�(��3;R^%�E-se+ރͣ>l׻��Qv��=>0�����7�����<$�*R!�����%�d0��%��4;�����.�|���"�L�i~P��B��Aa����&���D`��&���r`����i5/v"R����Z_��V�f������Qf�f�S3�Hs�׻����#' z��8�V�7��M �*�+�RN�.H#�
��03�c�~-�Z#U�����^������l��C���΂S=��Y2U������v��3�R�jJ��Fm���?z(	您�������X��y�[�-
�dM��b�_B����UgK�6"Tc�A'Z�"�W�,���	6 ��(ɣ���P�+ʴ���.�&b��VD
iU��?� ��mt���|.���{�0��`�	�x��ca4"�(�s>'�G�9F!/���S�����{2��wI�/|�N C7_@���@��:g�L竔8ᴞ�V�a��>��O+y���� $_%�����9J4DX��Jt=���~��~:�>��S�Z5��֐�����^h����{�������ipkQ~�H��p+����d�W=�����9�M�8L�w6�����ێqŏu&"���2�Ș�1����)��ߋ��VĄM�|�O�e������Rm��$%6��*yxHx���O�y�i<}uO�*�mQ׃�a 	�7>�*�P��FmR���~�d�+�Ots���e��6qݺ��f�,քϐ��fl\�JΙ=G�؏.�R�'4NW���b�e�j��ŝ��X3-��|-����]l��ow�\�$�B*�w�7�ާ��1[�r8*��)9���h.�^�}�ZQ���_u��_�]IeH4)�L�K�3X�=�F����q�� �d���T ����.��u��Cf���,��U`�b������_��I
hW����2S�Z�;��);<�0��+o1q��w���=��l�j���	�ܫ�;�� �|a<��G33V5�`�z������{�wm����aʫ�5?�f�&q���_�V�(.Fټ� c�� ���}�dy�����ц�����B�uݵ�%v�)�L�aS��J�2c2ꌧ,�Z��f�-�j����$l���^�T��s�p��og#�漉�*Om��?���.��Cl)��}[���-<�̎t�0��W6�����ś^`'E��͐ N���}�(���)�A���-����'/��-�j�{^2դ��vs	�.ы	R���X3D�F�*J�ň-Rb��\0E�c����r����	дޭ�5��������/�i��!�Z)Bh�L;Y�<��(����Ih7I�v)2�Y�V�2����U���!��q����ְWV:0�/sЫ�7�^���>�d��vYH�[��U2���f�����}b���sP�p��V����F��(�:̶&�:=���E�/H����\�=4���[�}$1:�j�D1.��B0�*�D#�+��f�͛X�:���!��M�@L�Ѷ�'F���+CD�Y�����AsP����
��&�a[�rv�u�%�b΂X[Nh����+��E,,��g;@�C�������(�#��H�������He�~���l�J课�}�T�23U�[�u�rq�E\�g�}V����6� &;ʌF���?����.�s���u��Ex���N&��,�mŁ/�h��/ǆ�P?؟����p7�OC����r�H���x����FF����+�p���5��9�P�*�,���&�K���"2��M���&m����W[��(�j�=���h	��q!'����>~�n�#X�$����P1����1,��ڰDZ�QKm�%���:���{�����iY3�j�3;!�"J5Rb��ZQ�K<c�̨�i��Ř�cS_�W+��Q1h����
�\����I^w\�;H�}�%X:�~�/�����A��L�G���B�f���1�FA�LG΂���R�:U`�Mz��� r��U&���-n\���u�@�B2��XAYA�W3X���|�i�P�.j(A��Me�������ð��ƍs�����Dp��tہݏ��oV����]AG�0�s��nH� x�X����v�\q��6��&�ɧ3����Xn8��*��06ߘ/�B�����o��n�|X�J��)���v���sMR�E��Khefؕ1�g�ViHC����[���p�������TES)S����/�i$��C�J�\!m������s���$�̆ף��p�F��"���Ef�2�'~�τ��<��i�OO,�_W��d�Z�?�^;CxD)��%gߎh0��&=�5z�q"�7$�t8��������C��Ң����NJWvd)�ȩׅ�|�ݨ�&L���4�w��~��Z呄�4S��:B��r+pK� �;�N�yg��v@���)d �ˁ�N������Ǘ2q��;Z4�qJ#��F���8Ql�w7��O+$�5*���Gb����r4�F��2I��$���<1�șYr�&o��1��E��j����v2П�Ik��&w
�r�`*�~�"h���F>2���5΄7u{��;���d�q���g՚,m�]Xx=��\w��㖹�b�z>����l^�+ӈA��ۘ�`$T�PR�mñ���~mA 8�9~�o�#d�OVl�Vp~>����7��5��%Y�������~��"��78!�v6�+���Q��T�q�K�J�n�.�
���f�7�dתġRN��+J ���sI�m3Za�6�A2*`�_�ɱ;�-\KAOX?����F�r0Q%��cT�=W\���1�����:��俦�Ӑ����v`Q:�E���3�q霶jU�w�~]�%�3�N �x�>h�=�I�@�z��t����k��J,��L�, ���eZi�{a��\#6v��wGz�rе�D��|�����\0����X"��ǁsb�t��}Q�7��]�«35xt�b�=牯W����vߔ���`%�(��b��.��^g�6Y�팔~u�]&���TA{�>
�&l�T��7�?I�$�*^;v6�Ř��/>~7��J�A|�m�^Z9�e�vU��K
���e�،�l2!'6H�n׌돣����9R3�@K67�r�딙;��&��c�rF��$�C k�r��0���D(��+J3`��߯3� J�)��a�A����&�2���Ǝ#��_ej>:!A1D���L��\C�=��(�PU��OfV���*'v.U�qQ��T?~�������}:mʝ~��H[�3rU}呃h87ʱ�����ŏͽ�i�Y�H�A����T���S���/���_
��w���-��ԑ�4-�ѯ|�����ӆ�~��dsh�υwY�!�=³;� �T������X��:P�J=���j��Bw"�[.
:���w4�Ufd>��xLET׵�8.��-_��VS2��now0��V{���S0����#���Z���?�;x�<L �LBP'��}�N�5Kf�v"SR_$h�)<whnX����H�$��I�N=�C[g~6����aT+Y����i(Ek22ã��������8��/��g��8aD�(������/�����ż�z�"��f#=CO\f��Q�lb�-���B��ե��Ԏ�;�H�43n���/��J6Vg&	��at�k?#�w:� ����D�B��IMr�e�J4^�3��̊1����PxN��&��ǻT�G�Ex�ԄBX1���Y q�-y�� �x�=�A5�\g#F�)�X<d����8��>�� �e�WR.���%!�����;o��Y�$!���n3���'ǓhO2��_e���~�d�$��EK��7�<`x<���e���ݧ��+��
QUq��[v�-���M��h3qҹ$�us�����XLH���\s�����Fڄ"��BE��'_�I�נ$�Q���ۭ)�t���h*�%��2p�Q=���寿ǒL����*�#����UÕ,������a��_Ѻ�+��"ˍ�@6v?���a2�Q�c��2�����,�i+ʏxJ���W��d�l�J�r����,��mzL5��R��E������1����H�.Kz�*��LU�+��H/ D�}��lV�_b]�.;� �?�kYǎe�����;.8ؾ���c��5*W��ϼK�u���Y@�`��S	�u������*{�ǌ����O�j�L�;�M�&=���F{/�-�|�:v�p~f�s���8��d��Ȣ��T���h6�&h�� or+�GZ���n��S"!��U��Vf4w��>�����c�o�ݙ��׆��*��s���G�1V
�Oi�|T����VaQ��~���S*����� � �|��׻����!�i�{�y�ba��q�w�������N��~�#�Z-W�S�����%9�%7�/Q=�^V����&�6$�x�8P�ek�޹�|A�=�$qNe㱭P!O$�&�Rtnpm�5P��e��Q��htij?9�<��Q�5�~#\ٷގ[f��B�ѽ�q(HB�Us�%�]l�x�8�&�;d��;b3��[(�L�s�ڻ[<�媪�B�1��ru��v�� ��.�@5���Wꦣ�|��Uj���d�ezKy�}�}^o��Z�h?��s~�n����Mɝ�}�F��!�b�<�i��ڄ�oR��u�GS�!������5N
��
hW&�����|.�� v�g������Lq��8)!�j9?����'�v*�y�G�$n �ꈲ�5��۵��x�,���ד��p��2q#��U}	��{M� ?z�H�������n�&��u�&�UM�*�*kS7�����Fl�������]��o�:����î��q�(Ӧ)���l����Km�|��Ry~��`˩E��k��Q��M\�O��e�>ʠ��p��eN�7F쬵l*������!���Z�Ϟ�n��O���8���t�E��r�ⰸ�6\ݤ/G|�1�:��XEoʐ��]��%�}�K��ԂrU	�b��7�H��ܣY���{�|7���N�&�Δ���*!�����)Gf�H�Г�Dc�|viZ��p=rd�A�*eO��@�}�S�/��N��sN.\C*D�}4�U�"OȠ�y�dMY��������g/�]�0lC���7�.��D0�fd�*���1�����ggt*>�����k��������a��Cm;3|��7ޣ��f�B��}Ga�Ts���Fqs����1�q#�W�u�����wvq��xa�?�'�39�'�?�j���e�0��\����*��/�)��;���-��\&�?�^|N�~���aq˟[A�&O�
��Wd=v�=��]�����7��
<�~E�A�ı�t-���{������oPSf^g~����~ �	�g�*��@Tٵ+5n̆���c��̌���K6k�Wa������#z��5�n�D�4v�6��5ohe��%V[G����Wx�� ��s��L�tv�c�%�O�QTq��V���6m��
1Aq��Ĥ����gZ=`o�(O�4��Q]�Ƹs�0�F�I>UJ?.����kJl<����c�4� ��-d\����y]~4��R�(�9=��`�YeI+�}���!ڨ�mn����K�8	��>�{�
Q��xĹp��S�c�6�E̞�ؤ�;���ջ��#� �=���i 2��Z�0A��bP��&����Z���Лu�[H��Bs��*/b�1@(��O�ZF�0�s�=\�j��nʼi�St^�'��q�IR&�!H�h��[�����3~��J���R��!���n��#�A+M�-����^~��|^󈌬I{T���m� ���xJ[e�w�/����.�?�M �-��-"<��P�*^Y.B�>�@�/s������UbRϝ�5����<Q��:
�W*��M1�f��w�du)R���!n�I>�gR/�p�s_a��쯴'����7!\�B�\��@���_�6 �stJ,�5�K'�	�Уȝ1��3�;Q̑�h�����&Jp�PE\7��G�Tp������JS�F�b�����N���d�]fNeS�z=��޸wDSH~��l�����y���d-��?��$?��O�����(�'����\�}��e�~Jr�-<t���6?�Ȍ3Q~0�l�6��e���ޛ�2>��*gU<�0����Q�K����s8@��o����[o趣qHD�,����0���%|o�������%\�gu����񌱁�s���N���R������1Ɵ�����2�B-M'F���T����ߙ䳒~s^n��[~�j�kQ�#�,�u�|L� O]#�j�\H�Ş�K'UQ�c�w���2n�S5�嘤�Z��r��K*U��՟24�$�gMA�����ʆT1G~��=+^?wr{�ܓ	S~��/����$�2@k����_�hd!����{����QQ��u�������n�BK�ϸ�Iqzo���<�gt���S��΁��~�+T2s�~NLW���C��q]1��[oS����<���D�dR�6�N&�z�ُ����J�$X���R-���p��~cC��bSz��-XM��O�1:�3�<894��(�_��Hkb��s3P�:lnc5-�\�����GC��'q����B22�J��}4��0T}
J�Q-��'|�����R�z���yU�����v�����m�CJy�U���bgi���7�^�H,����'�]�G(����P�6&N�s��~n3���Ej���,m���J�&�9��*�$i~4ߺ�w������`d���j��3��),�k��چ]�o��}���L�u %i�;e�^酼l��ͫ�<���7��p��x���Z�N�jn$/��B�����4��j�\t�%�c�;�,`�o'�F�^=�yR�5�0��?H|C|���R�wg~�,� �q�9��2�Ǝ�������GY�}r���{X��¼���ѷ�nG�?;��g���%�@��������HF���Il�
�&/��M��{� �?y�����\��FH|<���T���"'���L�+�
�g��?���!���r�A��Ȓ��u��HQJ��4�fR�w����W۞��c"�ׄ���.�ز�����9Whq ��/K9����M��Y�������A)��=���<��,f�{ʨ?��H4VN��w�X\�
�������m2���L�1��h���s�=��0�i��+x�V!��^���&//
���Z�C_��� ��0��g�1�:�E�K�}缸_�ߡ6W�Px�R|hխ,��)$.|�Y=)F���U����B&|�7/��?n������n3���J���U��P������0�
C&�GW4��+�ۡź�~�ZG���j���AAvE�-����:�;*���������w��Y��'5Ma���[��6�dO|��IUu��~�M�U�vZ���Ҋ���V��Y��Ń��M����6K�~i��!7%�������~�o���!	ý;�mi�W���������k�&Il�cC�3F῭�6~-��dj�ɩ{�Me��G����!ve����u���&]9׵,,��r}H�����қ�Kh��,�2z�c���3�#
R-�+��`�����X��?��c�Y�Hlb��o+\�3X4ܟ����e�1%��\X8wz5��k�os։?�[�jC��I��	F56ȗJW���S�zk�3���ro����3����o�&�asL/�N�
���[[�၆�J�Z�A~�z��%]�*��S���M�����������;[Fߚ�ԣ��֋���%w&�T�_X��B��,����TA��WjQ��8)-�MY��?ǿsm9'¦�a�|����|��{#{�@�Y�/�PU�.ԩ]��\n�$��W�a���p~dt*���-�d8��gLs!i�p�C��	��њ��{���=����<4��`:�+yo}.ʈ�$dX?D�'����j�Oa��y�T/��*��k�`�}��ۣ���f��ū������υ:�����3&\-��6n[���Ԥb1���UE�`rm���d�N7�L���nR�q��Kg�G�۞�j #�;���U�Y���������>jr���H�M2�S�c�	���Z3� X��J�W�ˑT'O�>]w�)/��wD�iۻ>���gJY����������As[��,�I&�'�~E�7F��I��F�rBRf�����[݄�m��"PB���>�^ͼqHLr/���@?������H8O��Da�ߗ	>>3&��l�ꤷ?7���L�OIIi�����LK5q��v��i���}6G��戞���ɇ��|�A!)�H%�R4E��8��م�4"�4���HK���w�����k��F�" (H���@�M��[ D �z�*HoJ�ID��P҄�Q��w_�o}����u~�g��ʕ���{�9�k�5��VB�3W��Q�I���{���nW� sk=��=�#gGGjy�~GE�sv�Y��$�����t����0�����Z$���V�)�Ŋ��GJV�4;��G�����\���;����-4
��w_QY7�<B}�|l���(�։´��>#�xϹ��罯E��g?d�lႆ���;h�Ӧ����;�a_�nM�e�ݛ
�5��0޽��$!\��� V�C���mY�1���ߊ$#���Dj����u�4�U��T��r\����K�~�1QH�U��ԇ�J���.[�XP��wz���fI�2`�zϧ<V�z�����u�� �Q[�X�6��+������ƚ�x���߰y���ϿXoؑ�u
#�NGl��u��|���0�@�[I{.2�K�l0�B.Y�}�"�{��&wO&�>����~��Ҵ&��&{`�N|�N��+p�_������h/j�1�R�#HN@�o�fئ�]�o�nq�O~��{���xvp�$��x�Z ���q��:��c�oًB4;G�sm���7X!�-�sY����FS�h�=g^�j�U��zB �$�#h_�q4�O�~o���Q�73j�@#��^��T�C��h=�4#P۹9�����kH�н=�q�n���'��v�/'�JP�eA�0�v�(�����GU��m��D̫xʘ"l����Y9��iK� ���e4���{mO���q������#��/�觀:�n���i˾�R�v��ϯӵё�6m53\����{���i�1�����y_tI}��o�;3�RQ��c�y�+T��s����m)?*�+���7?���Z��S2*�adpK^�=]BUu�x|�d���@L���sOm/�h'|�c�L���N[�q�ܾ��, �	�K6��3� 0��o�2;
�?�ý{��8�淹7I{�uf�#�y�rwV�z{����\�$l
#C.3���� ��r���%�#?6m��$� ��D�b���'�J�L�8?j%�&����K�L���ؓ�N���������<
rb���Þ�+K��g=&���5�M��0c�}g�{���"2K&�SQp��τNm���aB�)�[�'� �D�k�yi���Ee�)�P�?{�zU�+�S)@R�=��|Q����o �ЖG����aB�L��?
�̦i�O�؇����A/���RßX8=��D���~Cnî}o�<����z�������[}��
�{C���}M�� f=*�_�1<�OCJJ���$��@�hIQ��$�d�R�g���Z�f�<��N1��Ӝ��
�`�Q��ί���}�bv,_,n�~㺗�]�<��8�$���í�Y��������^���ʚ��Z���6��������@ͺ�\~�5�ĵ��3Е���/d�iϥBh�l���(��S|
t�vC����5ST �R��w���Z�9��&
���z�w�R��y�~�>���"	��K���:�!g���Y|��ں �����w��	���HK	�>��gL,�����&�tL�QIw��a{�N���C��rҠ-k���-�_���R����-���x�c3g=��5�&^S{��e[ps�OSh��>��W�s�a�z�{�����f[�IN }�+���� on¿���9$�JR�8��V�ˠ��O�D��tY�����Z���n�.GQ�=V�A?
;#9�fq�����
q3ф��:����%�iZo�-U�����|�N*��e��� *a��II��{��OǢT�b1���2%W� �x[SO
Cj�G�>���EnY6�5$�1�a=n�Xx��~$��G�jJ�y+3l�f6w�j��Xs�E�v����M���඿��:���9�����ש�ӛ�)`�yS�ݻUP&����9����}T�0L�� ����ǣғ��	Le����仆�,��j��F�_��NFއZ�tE�iyǐ�_�"���@�a�E�(��AU�=�&�e�/��7�_�Qj4& W�DUB��(��ss�����0�bH��������ܐ5?��-VlN�2���Sv�0}cX��jZh�D~�ߊT��z}����~y���)]�;Ѡ���%�e��Wj�7'��5eP�MV�B����}Պ�h
������K�	�(%�f���6<*[�oI�D����!-%��׹hU^�c�4L�t��?��xI����a��~䮩'�� ۑ&l��b��[u�T��	�g
4�(B}%۬���ۚ;�įY���:��Y/����Irr�lL�>�o�7����WE�p旬eؼ"6�PPn��Dܧ�W�����_�������6�&���������<q�F!jc�P��	ˌ%k�Zu� +�X�z�c��@͝����֯Z� %�-�2�
cF5�9�`�-'���re��@��)sʖ��1��?��`������a����ܛ[���>KC�C��2y��H�E�>"��o.V� D�#̕���W��� �I�ی�Y��':ꪆ�_5���nYDQ�W��L�N6۟Hb�o;}~V��GS6�=�*P�������OƁ��ռ�÷G�,��35�ѐ�0���Ư6�ж�+�k�yY)X?��j2����N���Dkr.����,t�
��M���,4d��b8���v����]֢�M���o��Լ�l�;���8| o��x3?� �V>圏G")��n�GF�N;nVE�I_'�JW0Ӽn��gp�5���痋���3��dC�|v�l�1P	Z9�q~|�{U���2We������40��_-�,\�OV[=�7���O�^���?�( ��z���3���Xw3�(�\���-�s����M}zJ;�oqi;�3�NITc�*��q��0>�vuR�sZX����Gp����eE��	�+����d�Ün�d_�N��kuz����
���͍K��J��8o��o2��%#C���G�9�� #��gX3wZ������kS�G��mf�ڌ˂	{<O �z�����RO	�)�� _��&$��E�QZ�+��Dp`@ˀǌ��9)�%_�7e�!b��77��2H�|`����:̸�U5b�lf>�������d 4m�Y:�@Q��gQJ������R�n�5}�>"|Jl/�/}U����`��L���w�X���S��� ��{���t�7�ݯ���woU�m���+N/��8��e)�ؕ�nx�^�§�I��a{D0�>�k��Zc�אDU�-���q���R�p��~I8�Er�b5���̹���R޸�:[�����D�El�U�DǸ��=��A���$��L�OC:�)����Ԩ`�Ŏ��	�JK��x��d�4����Ӟ愦u��;�|�;��P��k������udo�U۝&g&����:��o�l"�	$�:H�D�����m�1���:ow��0e�>(◖8[L9�/M�C�V�v)kz����=GĤ띍OG��xs�]���9@oW�k	[�{�滾u�����jL�Ds����)*S����N���p��ĵ�uI���a�m��K
�_��Y5A��t��c��0�bY�G�&7��:Ȣ$M2�������&
E����+דg5�ܐ(p+R�=ͻ�<e2���\���t G�	Am��k��H[`T��h4W_�g��)p|
�Q�9���3΃���~ʐ7�ӏ�3�zY
�e�&���T3���h�h�z�s��ZD�9�0|At��w�Z�*9�����=�'��-=[��z��XV�%=yk��*Oߝ?Ð�"����Jjܾ�{��w��%�$�}�,{��w:=2�rR�Ē\��ڶ�ӝ��Z�L�����dv�c�T��Xi�=�&��޽ �O؁�=5��� \���dPs"Y��8���U�ǡ_���A;>�<�#�I�b��� ФZ��k�uB�������j�Qn�a����/1/,0�^P.�g�<��$;PM[?^�������R�eKCN�Rp��r���o�o����k�;��r;�4����n)�oiσʩ��OO5�w�y;q{��PU�B:��&�%�=�_�}�<�Ѵ����ǩmr���q�,;�91�]�9/��j ���"�&o�L&���ǥ&|���xN9?
=ڇe�HL�.˧�eB�D�kn���O��*�n1�5�{�Z��̅#��)���qɠ��,���"����u�ϛ;��ӵ�.�����Vk�^��{qI�_�Z.��ô��+j����m� T����e�Q��9�q�T�?����<8�ڂ�u����A����F�Ŕv� �I*X��z�вX��w�4����:��գ�	b�[F��^�4H���/��b���@I��;ᵥ������V�^c�	;oY36��:��f
U�u�#����pO��
�S�z�Z��u`J�A�yKأ�o+�w����s�>�'��n �5W����n�� Kam"���6�=�˧M�<�<'/x6(b�����t���D�$A��Ư]�q���8�ŷ�͊U�K�i%m��;���!��ݞK������])W��)?^��^S����6F���'�3�߸б5æ�'䱌?�8,�_WM� �z{vm���O��x�����e�s���p"���8���L=+G>xuȸyǖ@	����5;�w���aj��I��[-����>x����W�\���&[J�>ypRɇ�D�&�Zf=�T�s�Og�cl�z�(�De�g���^��B��_)x�j����=#�j/����찚�Rʄ�b�f-�l~��L��D��<�������;��(ϵ��q�z�tC�������'>c��QH���^�6�z � r>����#�%�{h�+?R
jB�nq|�����j�{��1��Y5����հ�bN�q�5+��G�a����C�E���cDD���f���)��DB	2��Gs�<Qͻ>{3�5��'g����׹�9uM�М�"\xM�=w�BF��+����L
^5u��I�3��������Z7�n���#��'�W�N�Nd�b׀X�a�51r
��B��O�A/(�)�o��)����dQ�oݶ!����p�ɺx�;h�}V�t��R^R��L�ke�/�iw|eq�k�c��.tѻ���V�9��"���7��t�z<���/���dc�������߻���D�b�Z��M=��USUM]���m.30�Y�$T�r��.��g�Z��I�gAN��~h�3q�Pi�]����:�0ŇPA��!�!W�Q���D��$��I�H�m����,B��'o-B�;���[�����.�� I*���s�P�u��,`:'�,���PS�چp���]�s��+,����_8�9�6tj���#D��Sڲ�|��2��ӾO��n�_&@��Ny����:/u6�Dz&�]�wBaIf����Q}�f}�{y�e8�h�cq�j�����;3�����؝�v�q6➁�,a��&k��i�Qę�uc�2	*12�	}^\�Kޠ�~��پJ^��o��3	5��k��Pr_��;���yU*�<�$��$�k�7�X�0;�G������w���U�� �6����ǖ��u&���M����ip�Ǝ�-�{�5|�=Oo}Y_7���v���4堢aփ��-G칤����������A�;f�ڮ}G-7�L�>�����������٦���o�*�UU����ЇE�#�8Af�$�ev	����E��Z�x`t�!�Z/mI�}�kH��k]w{���v�my�����/��I��;J���R�{�$�(8J�ݢ���o/����|�K�n�>mk���v���ú@���-Tَ�/�'�����R��7g��;�1a#0�N{Ի�� ��_��T�O��We��q��.T���M���{S__�0*Z���ޗ���k���.�.�)1[�M���oK5����ιi��8�8>��L>����{����V��^�R"���`�{I�|�� � I�S���6��c���Wo!��>	]��K$��_pz1j�ʹ�=b�s�������n羧^��s���+L��]C�^c�o\C|�{X��d��� �����}�x���ur
\��"
(Q�qe��2� "��8�ka�n���@A�*I������䒚ϧ�JP�	�ȊM+�ťmy���X����F&�����j��4xq���[���Ô�͂�����&�ϊlp�Q,�2h�e<���e�-�6h3~4��e�&*�o

G�ӑ�6���Wn��j�p��}�es��Ӓ0�8¼�z��Jb-u�M=��5(3�~�9<@0��f��/��u��u'��*�W)DFI�o���F-ai�N����J�ɑ��75֜�rua������n�T�����#�O�� u׮�bl�쯕�
�'$��t�vk�@�DZ����zʅ֠6��=���{֧G}�M�7�$eW��e��O\FX&O�;
���E��:L���,*�8�4��gK,��g���3��{>�hQ}���
B���{�B����"��ӗ��~���)|-&�Y=��cmﶪ����#����F��ݠN�O�-P�C.Q ���T�	a��G &қx/K���@nϴ~��}B�؜[@� ��KL��4�rY}��}����h�I��A7�gi����|���3�����]'�M���}r��^X\��F�[�#3�;h���^t��7�*g���&�A_��=�ƩERv��w�>������X�R���)�����N�αoY�YZ�O��\�8��:W��%s@Xf��s�?@*��9V���JN�i�>
W6&�,?���%Wq�/s%�<B� �tG�Ƈ������8V�a�I�ymym��&C�u[ITE&{�0�}z�DW��]�y��Am&��J���|8�tƴ���M�oH��;�W���)ճ䬄#I�%�eF�?�S�ր���,�`�*�h��k�ah�i]N~����ݫ'^�FG�N���b���R>��p3�1�*�/h���Ovy0��v�5
mf��E�a/��Q����|��1�4#칶+C��u���J�s���"8r�
��/7$Wu�%��~�)�3\��:���29�Co�щ���S�5�Fn�Bn�g7�#o���)CB?ߎ�q�n� �1��`�R�x��R�I�+�\A�:5�}�^h|x��A�R����2#��{�7���'�f�4V~�(��ލx�k�SB���E[��W{�H.g����?PR{&�x�!O"M��!�n�{�U_��%#��j��]>�$V$�3����K�p ��.]�7I �[�"�^����_�$��� �3�$|Kt��K���L��F.y����9ذ�P�#�ĕ+���q[��_��J�ʊQ���< G��!��߲S�U0����Ƞ��˺fM��~;3���.�r�
��w��|"mL�7�,�ؘ�<Ӯ�2J��$���q����*M}V�c##
BMޓ�{��3aQQU/�n�c����Ӕ�ܱ[�::k�.���+�5����� �Z��8%HWo�Lnfm���uUF_.KJ+��޵���35�߾��?j.5�����Jbϼ'_KCV
Y<�dz��� SI���L���v�~�p����~���->��>��oX����(ȨH��쳭MW�Ķ������t�?�.���[��V��6�C[�?be�K!F J�F�DL^��fD��Y�Y���'ͦ�Iȋ X�;I%�����rݮ��Gq6��K��f#�(X�B�8+u�mS�O7�F	�4�/2�=�ON�{�\7�l��ySr�!e���MUp��#�E�����88�)U��f�(�ҳ~$���o�0�H�8� �џ�$�-����.~]ϧ�?��>w�6&�b5ޛ~BGl��4\Ǒ�q��g����$mqW�Y�2��x����������O�:��;A���˹߲��m�S�}PWZ%>���	���O�k�R`�J�ƒ�S�0T%�8v��L��÷�2u��#��*Ü۾����>�R��+����$1�_�ȁ�Fz=oC��,�����^t�C�n�s��u&X��"���;��%��x���/vLS7�b�S'�tu���1GRaϱbs������/�����w[ĜƖ��ANRL���kK���YuK���90E
1�G�^O)d�v����g��:�/�����Z�{��C%�]���?��ނq�$��Bg �@7~żϦ+jC��.�J�x��ݬ�~Wkx�T��4;e��� ��\Ns��t���`dpu��!�w��vSVD�k=P��-YlX�2�T���b����H��z�S,��Z`U�-��\�^�g���w��������P�~�Å�����u_��sH���}w�r���ӎ���1eB��7��u(�{[n�6��Ys�Z���44Id�iA�d��E����^�#x̪V���`���G�5۟ɒ��mW�$#������:K)��KMW;7w���?Nf7�i�s�D���T�=�p?6ʻϓn+l~�X��" ��i�r,�O*�j�)�w�O��������H�w~ڸ�_H���\�@c��,B˃3;��;���^h�;7�t���4��*w�Ag��&�q���=G��cLX���/�%��H�I�O�{���%��3��x�+M�8Y�+�cn𶾩�����̬�u�f�BEdM��۱�ճ���<q <��~Z�`�޼fyչy��㓃/�.�1�����J*��&vk<�7(�W��ee��2aÑ�@ka�~DB%"ޝ�yZ�~}5w�{oېa=�Ec�iUXK�	�ӆE\�iN� ��&��Wwwe��t�M�	�I��7 X����~�[#���]�O��P���Rb�v���S���
�
����FO��'�^Z�r��O���D�(�H1A$ �x��ar�Al����u�R���fՅ2K�K��
��{[O����
Izy�}�<��v�c2�������x�i���L�<�<�q6����;�Sj�ߎ��.r���x�p��!PX`Z�P��:�t����1m��a���)^�g;g'/�{��p�=�;v�a(V(j�`6��m��Z��/F��5<
L� �#�v�3#0Ԝ���ZGxL�����W�'�-:n)�2u��)����O!����Q��H6��}X��G�zp�HU'�D�O-B�X������N�X��Ƴ����4D�C�,�֠P�1i��P���I*
½�,!��3��Yܓ�Q5��V�p���з֫��Vn�<�o<L�k���{��qgy�gۻ���#����x��/��NY%:.E�`E�j[.��7�����F_NFu1l����`_��d��L�IX9���M���dڕ���8R�H0�mK��3itH��	����wc��w�(!�(�n�ל��t�~�`��C+����TJ����W�,_}�s��	��ȸU�q�������-	�����DT�*�#8\PAyِSͭ�z��+B�=�ǟ>��qbj����_�d���/~ >�=i�Z���V�|Q�&�v�P�G�	[aq��Yi���?J]�x�>�},��̟�b���tO����	fr.	�F=Fi6~Ao�ffM����z�H���zl�G���jJi�v��0�}�SB�%5��$Zi�1}ݍ��E��E�l���G��WQ��0��6��9��CJ�D�a(U˿�|�����ׂ§tv�~E����"��4ƀ|��<߶�.!h�'��t/{��h�EY�B�a�0��y-�i�@�*D�?��^��:3�EZ}X���Fa{�:G,�h·��r�z�7m(��sx'�H�Q�)�~]�.0���sZ`�%��Vi0)� � e3weY���]0*f>*�UQPޫ�m���|5ц.b�!O}3�y~�֓�mG�K�r���:��l�D��w�׆��tr���a2eŎߠ+��R�?��4��->�s@�c��ceeV��o]�P�GZs/xK瞽՛Λ��sG�X�2�=�3��r��u��Q��^�If%��BԓF�o�F����z�\;^��sꆻ8�٣�ǝ��J�x1���	m>86�Z���;]0}R�YzBlN^V�X��0��?�9����ѴN:X�����.&#��¶6�EEh7��X�5�W��x P�����҉�;W��`�9�?�i�Yr�=b��	������R#�KEV{G�ܿ��p�e@��2�c1O�޺'����[�?3���)P�Y�c!U�4����z���n�;����?�`C�6l���>���Ծ�Q�Y�Z�x�ϖYI,+C�J|JT"�\���{��E�U�tɬ�&����;�d����{�SD,���X��t�I2y��ʹ���7����g��m7Ìᑝ���o���8^5<#?L����;��jnݶ&Vs�f?1���S�'ɢ���7���tN�c�z�!��*42����B�R�?���=IV���F"vFػ��L��o���ԫ>s���$�^��d�I��˻7d}�})<mN2I2;�`\�7��bH��[�[ cvp���iXS ��r(�ﻜIt�	{�Q����qr��4q�?�י1��f���y>:)�֍δL��o�����f���^]����E��5h�,0�Vw!����3	Z��E�sR�q9VF��;'�vKf�/���_g��^�J�,��@���7�Yw��9Z��G.ʻd��s�v��"2ϋ-r"����I�Xm�\��0���1
z$����ꁺ4$���+�G��+¯H��d?�SJ��R-=�
I��V�C9	�nA9�}ɝ�B&���O l��=�I�R��}����(Z�zAo� L�IԍB&���r�[�ܶgo����Z+Z�l��~kc�\��-�s�R�4���
��3��:��ў�Jb�L*��{��f�1�,+���?���B1Aagutb���F���V�����-e6�w�d��p�s�2���]6 ��+j�R��u����d����"͗K�/�/�"p�i�(��&�	b/6��XƿS��0?���@Ù��؂%�A�z�I���ta��d�I �6u� �=ir��+������v'�%�}W�+�k��m��)$�*�wN���q���t�v+n��V��.<~n����K�j�굅��9��kފ�W�!O��Ԡ�j���E��Ky��|�:i"o9�=|F�ݦ�\Z�"e�vmj���nu�G�?��g�t�y�נ�V~���%9���pO�!���z@&
WMp1���	Cm������0�.Zl��1Ʃ���dݟ���GRI�-�g�N'7%'�3���B�H��+0�i[�Y���P"eW��wo�$SN@4��<a ��RRbN���2�s؞���,�L���4THt����������,�snN���Ur����=�b�F/6���ow�k��nJ���ߕ~���Ͼ��&=�!�ax%�`7l���'PSX���WzZC&!,���g�{��*�kG��^K~���Mg��I/�j��Ƚ0OR��¦�G2O��{6ʍ���A���Z��G�w�{ai�VT�JTd1Qz��_%�P�Ԃ�N<v�P��Bi�ח |��~��i�a4"r�)$^4)K�$>�I�)��5�Y]�;t�v{���]=ز#�5'����7㪘�=!C{)�#�'���i��6���M���z;s�\����{Y�����֕�؈���<�.'�xV±dZ�q%�Hi����7�N��]�����!��&��{�ǿ\��aYWW�S�ҭ�	71k��I�=��$W���1�FKE�Lz�7m�ܞ�ʜ�=�'��* 􈳿*�#������-`^���J>�4FQq}ҹ�����"�z��hp��N�QS�{�`E�Gq��A�}��+���t�O�ߜ����1������>��������3)��X���{��2�Ou�_�¢��z`S�T;�u�G!���kj�1ar������$�h������\��i��Rh��?����=?G\�d����6N?>���diU��ދ!!e8��y��5��9r�t��{���H�m���V��bJՌ߻<�7�G�J�}JL�#.$H�[k����� Y')���s��:З�i	A�=9��EZ�ė#�����+�y%i��ZI�u���UBa+�zbU�ݦ�D����e=ĳ<����}��� s9�
�Ğ�qP��U05�R��1l�n+��x��8%.�o��K�t�u
*#,���{&��:��������z;��sp�4�wZ��-�1|�i�g�O���X�'A�S;��2��׹����f��QKA�2����M���D��j�T��}B W `��w��M"�e����X��㿱7�7I;���*E�����>�6�Q���/q>-K���Rm2(S�eQ:��f;"V9�_�\7+����Q;ŋn4,{�������k7/�����b�E�D�SF���Z-�磗�>�;��˗=`09���0������7�©Q1��}��/u���{'��vo�U����&��WX��˳��[���r�����m�g�Ǐ�Ͼ�/����<7�(D�ok#R#���+�x��U7/)��{4�=jK��(J*�ۿ�{��͢PwP7�ꮼ����(�{ ��zi0�O�9ǥ�p�6"�sm�PcP��W����$�%ɟ_��~������A��XHc�46��T˺W\=�.��.�
���:w(	���H����?�,�X�{�F��;9#�wRJt_�JJi
4���H��V��������)� ��������x��	�Klk��{�BP�����s~AF� )A�o��·5j�����5c�G5�K�W)�C:��;݌�4�����W�`���͠�p����̢n1�&-�zw!?�bzm -`�y��hxy��),Swb7��g��}�~Qwrչ���q��y �eҋ��}�/~���vWԾW]B�ŵ�bǵ~�&�mFV_>%�ڬ�@�eo`:ԂO��r�����ha���w���6����t��c�@�����u:�W�b��4�]y����5%��R���Yy�p-�t��D���N�L%m�5�s�u���.s�N�	]��==Z�ė�-7��Ȕ|l��y�WT��A���1�.:�Y�a�-�A�2�`�>���it`�O7e,� u=��G���}vEKgbQ|n��P����%%��F0��R�\�i�#U;����%���AG�B���`A��� ��M��:�֦��MՐ31�bw$��<�w
t!L�.ml9i�g�{5N���>J������ \QIz{Q\���X��;�˳�k��}���o���3֚�|WP�Y����!��'���ӛ*'�U(̃��g���q3}֕��b��xf�R(�t�n��i����g�ӈ��9t�%_Z�	��\L�JO�ص5Ơ��S�/�	\�]��lqg����j�;�E)�4�R�K£i{n�Ъ@Ӈqӎ///�N�*8�oUN�*�>��uk�Y�Nm<�ȟ���M�l�Di�B��}�j��OJ��\g?�rK�\�ű��ѕ'���.>|ˣ��^ZXN����k1������p&�~���d��:Fv�w�:�E'�$�=����~�uP���4�RW_���|O����X�mD���ט��Y-�p����D�U���ʎ�:�+v(�.��?8[�����n^լ�m�?F�?xv��K������D�(��l�ѕ�w�A��l��wc���(K�ј̜72v-�x_���}"G����5`�bWڳ�ٻW5��.�,Zy�d1	y�y�l<��H&E��&F|�.P^���r��T��W�@�+��^)�{�B8W�F��)?��˥����������Ӕi�%Ϯŷ?�^t-FL���N�)5d�] �H�>�|s��ߵh�ҁ;�겑�Iu߽�;N�ɕ��c��aCƈXM�f��'[Nǩ
���O+J��HK{C&'4�k�G��'+�=�p,��7`;ۨ�8�XΎ�lb/F�UK3nf����f� vd��aT��+[�11�� O��H�sݥ����f
�:?��/*�9A0�o��L���"eq�+�є�/oT��Kx0�zv�>��L��-p�6�x.>�f����޳Hܭƻ%�Q�>KI#�6�GW��&���tnp�C���3ֲi���.˂#��D����������Ǡ�O��n�����?���/�{�0[�ŉ�2}�� �w6d�/M�E�j�F<^҈���Q�*���d�{��'L|�~���A�K�Xd����g���W��--?�L�K��Ŝ��A��`S���Z�Γ{�]j챩�)���[B�ʴ������}�p!5�od�N$�!_v�������-]0�e~3`�X"_�T"���r�B���T���	��5;g��;R�����ԗ�C1f��HH�'ܢ "B��$S�uy���
�R��z!��f�_�M^��B�h��~�zb]��G��Qsq�Vo�	iV\��ȅ��7{^{�O���h�<�:�z��1�o��~r�G�&���f��Sn1�|+�T%�9��V�� J9;�D:g�����3���⍴���,�`�4��o�V���P�kOr|
��MBF9��ي�L2��8�4C!�)dwZ��Fk�.�<	22}����Y��d.≏�{?@Sᢠөݤf� �+�Y�H�
0��
.\g�h�!��^��~-0�U4���ش^N�L�y��d��;;2�x��~�8g�tȹ��f�R!�	�� �19��E��*�h���*h_�$�f#V�٤ֹ<�����yGShӴ�S%��\Pw�w��LC׌?gPY���(Rʮ��9,���ֲ�$�Oa�=��nr�Y1�P�}�!�x�q/g���w^�Wh��i=X�z|��ǘ�<Z�])�Kf.�=�T�g��al��`i���Y��m"�}�*d}�f�5gg~��mш�ڮv[H&���	P�WS��ۂV:%���Q�E1{�C��%
��`9[x�S?H�F���jŀyj��{�jv(.�u.��*��rG�'�c���2k+q2���/�B_kݼT�5��<�/�F�>�v�2������x����1b%PT;D+,�d�|�
���.��%\R��&+/~SSҕ��R�̚($�:�G��G��Ԟ,� �{˂q�n�nߔ2��3\���l�
b}S0�i`�|Q̗+]��vV�}��ɖ!k\�����{Я��fΚ)����nþ�T�iw�E�oo4��ű|��^.�0�)����TrUF�����L����S���K����<��(1�������ݜ�t���$:5\~�J���$��}m��f�#>�#ˠ*_��Р'L����ax�}+���2�j/-V���ľ�&���y�m�Bf�	�'�mnk	�e��q;�����2��!����7P>�O�a�����5m��B-�GS.
k�,.r���sO��.�z�?���^�x@%W�( ��S�<�Y���^�i
b[f������I���i��٨xM��s7w��e=]`�XP�&,�������ƻ��4�fp�������mM���z��9�d �`���hUX��ڹKǔ��3O���n&+If^��}���H$�������!Nc�f�؆�T�o�q��r>�:�M�t�(��2:�.�$s��(!���{4��w#QOBM�ά'o%5>�tt�Q}�� ��l�a�	�	F̈́��˥}����d����_d���~%DV�����[�7C��><+Ǘ&���5��s��O8|��[7����r���p�t�::���?���>�mB�!kJ�)��s��伷�kX��3Z\h6<�ݾ�m}����	�8;��靣S7XMRj6���8��4@��⽇p��J���R����0n�t2�(�&Z&d��jOuF���0��ή��C�(��A.���y��"�Rh���pA���b�qj�ʀ�xw���~�������Q/���S���8�gHY[���#�x����JW!��6::��x��N����ჱ�52[,񮙴 ��;����V��3
�]�FȦqz�y����2n!\fa��a�o�.�Ğh����g'����⻔�5��6V4G����%�� 2��Y��iy���K{F[�\V�#yY��r>ga�/��Lc|���C�X���A����+cD9�Wb1�W�;�o�?����[�S��Ο4��О����-ńd�p��㳩	��.{��K;=8���8[v�0f.2r9g;D�X�o#�=�4y1�/-x�{8=��D�_]��$����q�����-FV!zPG�u��H�ӵ�����N �(�!����b����� K�EYq�zh2W<ǫU6ܑ�u�����k��o�@��#���EC��������˳�����@�C"ʘYHTJ�:�]{+K!=��w���o��T�|XSx=^����ɦO��(3
�4-����M=�Q�# �so����{��j>��H	�w�L��c9ʚ�����t.�yІ]��i9e��sO�������"����e��ڋ��]џ��"�r$9��)h�f?�XO�O�1{�t�J���!�I�d��cq\9&gՍ�oMJ��H�?5�e�]���B̏�|7�1U�̋��Q��V��Fh�2=��	�>H�9S�*ax>�~<�ȝ�8;����L��ϥ��η�3��q���;R��;���P�La���JB
��&ǒ������99��x3&4*�F6Cc�g���~ݿ�y^��z=><��k���s}>��z�?�����t1f�~�¬�4�z�PV&3����S�S���?!��e��אO��������_��_�� �S�_��'4m���0��c��yp��@��(��	�3眤P���SHH>I�J��h��+�9�png'v�ޫ�@Sꍚ��I���׭�d;����e�	q4V�9y�CXw���P���ͽ�Jg/�\�b��k�g�Cey��Q����l�<k�'g���ѧ	4{7' �*���.Ň�O��q�Ҥ~H�SiVz�Õ���`��w���H����]�$F�B�lDힲ]��ފ|S�e�f�����[r��wRK�ue���A�7�G|��`�-{�[ה=���K˩[2ݜD3��J&�l��c�=�:xed�U�����(�aSԣ!���y�w�d�V�
�K �2��s�G/��w]�J���w�J���ӟ��R���5�*`���n`���P�C��~�՞)��4a�Uro�?��3�	�R}��D��ћ#Ľ�ߨ�����N�Ă�J��|���Y��4t*�V,�e��k߃mJ��p�=Rw�w��	ocM�d�I\@�`T�Lb��x�2����G�r��M�R`��UJ���B�P���j��ԡ�����!��Y��Њ4�����x?ڃ��,[�Al_s�jԇuFo3���G0w�K\�m�a<�tTQՌxdס�0^y��o?���L��!�zݭ%⽍�l�M��k�?2x�g�K6�(�Q��`�K�4x~��w�u=�'�E�+��q+Lx4��[Ѽ��q5w�o�N9�n'\TB���m�u'���Y�Z6�|b6˴ѻfG��M:l,[���F�s{F*���mg�h��Ć�oժ�UZ��zi=�s���}W�ԣ��Ѕ�fql�/J}6��M��@�ϵ%^�a&��EC|d<�.Y�����N�\�1���䬸5��\���I*�������u��ZNl���=T�̈́��w��H���n�c��r޾%�k��bj�܍�.��*Yd��T��	@��Ӿ6B΢m��Jܵ	�|ь΄�E(�HjPl�PO�	\��7~\VV�<���]���6��)��u��4)�v�>��(H�V9�|��G���m�X�Prq�� �$�{�ן���-[1n�0t�G(�k�!D�,�)�Ŋ&���5���)�H�y��H(�*�� s�O�ʏ�� V`����.It�4�H<v0�Q�*���.o3�9��M��k_A�ǳ����nu� ��?z��P��
��N��:���D��#}�iT�`��p�m1�����a3�TUSA�R~@�2mo�r�ڴ�c���B�o˕�DCc���.F�jH�����s�W���҉��,��&�vT��4���	;D���������=�+	�?L�)[OH/�%�uw�;˜�Q�4�2������(������v�͘7����h���K�@v~W�����z��)�W�=/��u��
?����$ �a!u�:��NOva�-���u����ܽN-��8���rwax΢�����~?fߚva4<��>��&��e��9K�5���M���.�e&��̭��.�1�J��a�����Ŝ�@�<k�y9>����%b`��T��Լ\Ne���P؈�ba��.�`���� o��K�&,�+)�8K���^�\�5�JĀ��lC7�1\�T��EN{Tw5^�	�jօ�Gg�j����"٘�>��Z�W*Nu��{v�~f&��?����%���R�i�N\��qz����vS)IPE���R��2Z���W��lĳd�`��\NKt�_߄b;��l�T�d|I�a��.��
s�#����٠dz�sV�g`�V��{�C�I%z�S�a��a�ƣ�1�.Cm0�{��:�Jv�R�h7����\�Hgu�cS%��pS��p��o�$OˑC�Z�e@����	���AF ��Y�mdlϤ?�)_VmP�[Ɲ�8�#�����{W�&�_q5����7b{������z�K��y�Ұ>9��A�ܑ�v*R��<Y:��H�j��t�?�F*����m���݃��/���t��e)��^�����,;��!���|d���u  ��iG��ۚ��lC�3�K�vǏ�@��3�	?�Kwr�����8�x.3c[+n������Q��y&)PIP����I�(0�Ll�^�a������@��TTJ���FF�N�`�d�,�2\;����'��R#Fa9�-���P�ySJr���Q�(�AP6��Q`a�',�f�h5�)�.
ap�[���?I�#���9W}$d��H����+XFf�F�y�S>�9�\���������/vq�)ל�~�G��� Kbj�5o���9���i���|8k7 >�jfxʣq;g����I��<��\�U;o�M�ο��I�͂��(cF�_D�O�Lg�&�|s���8����TV�00���T	CU�2��g���-�k�/>�]�*p���L�Kj��i�vb���' ���+(n/q�)� %�4�hb=���U���-�s�~I��/�p>�qD�ߪ��#�D��{܀���h/��5[��;F�H�8���i����F��;X�Z֏w�����B�T�o��V��MM5r~iW5�w7y�����Jv��Xmv�r���^[��g��#��vj�ޒ���7�{��M�X��`�N�ģ�Z�R��7Kk 91��T,�+̒Q�e�A�ʸ͕Q�9Ft6B� �E'���v��4�'��?m�(���@��9	���xX�޶K�h��#�B��L����C�N���;,�Cs��C:;���\�v��������oJ[�ɡ��O�^^)��װ�{��,���j��?�ݽk�P�@�s�o�A��]A�0����x\
D�	ot���Y���"OG�ZC_폟�N�k�J�D�����]�B�M��E-u	���0�WS��G(9`�����HԀ��s8R��&_{�i�\h��8Q�1��g�Ŷ�/눆��z"XE�V��k6U��u�Wgl��̆�O8 ��⫄ɗ�*<��V��:��'����Dҙ�ڿ�;� �ޫ7����V�$<{�!���YS���X7��lY����Cmc�1T��*��=-�>�g*�ۤ@���IT����)O0JW��g���I7ٶf!4I��ҽ�w��؉X6�c���L7�%住;�b�k&���	e���5��_��"V�E��t�nKBؼnnZ�b} ��rS�y�{���6qE{�te�1ǹr='�7g'����Vx��@���ѥ��gp����!�Uw�����ᬯ:�Sg�8aa�T
�qs��(j���nو��X�I���&�k�׾c��F����GKt����H�h���z�|���'�T�l>�s�j:��	�џr{�0��:@KZ��~+>I,�uH����R^!$\����?;�U5ſ^7��#[V&39������]�"�������˫Ƃ��$ф�>ß�zH�>2k��S���[+�a�R�6�N-�X�dsS��z���7�Q��o��⨕�i۸F��|O͢�$^n*E�`m�1�����>�n�1'ȶ�M��ކ����u����Y���(҆#����7sUS>oD�;"fy�1U�.�]?yI��p�M�ΘY-����wVM���sk���H�~�NI��@|WW�����#0jHA2����1��Yo���w��+�{b�#~wb^>|;������Ҿ[hy�]�z�ο��fd��8�]���! �Qk{���'�L6W�7`�c������C���<����쟣�~���.��Ɲ��˚B�I&�2C�;�N�\"�`�u<7 (��{Ig��	}"$�$'F.Ō<�>����~�&v�%ڰ����|\Yo�^�ݜ��նl�c4���;��]W4���ߍ����/�sfSq�Bk`"�4p[��K5�`���US?�`L�k(7��-r�p|JV�s�����{��d���[��	�'��J��G�-׎*��q�l�bC�_������*;ݽ�}�n(��M�v/�� <�-2o*������S��G��b��Ī1YкN�k3���c�A\�yZ����y�'V�,r���҆{�K���_A�[���j3�!d#�Q2vp!����3��IK�'o�����d_�J���������mk;������qU/�#%�3ίQJ���DU���� �bԙd[~���=,�w�z*��[#h��A�0-ElZ��2w������=���
]�-���JWҳ��0�p^#���+��/��,�^'�'_K�sFv@���J�C�z7��h
k�픕������М���n�����}�|a��̗oq��x�ci�̤���7�
:h�oGaAWڨ����N'�S�F�/�eBoE���}�z�S��1{�l,��JD�ʆ�|���KU�G�-�R��]'4�|�8W=��c�@�ح��g+�_L^?/�!�+��H���a����d����ll�'I=�Z�+-R�>m%%gϱoA ��K�'F�J��7���pz����f~J�C�\֟����1dDwb�o?]�ɿ�}��#��ٛ�������@ �Pr*�2>}�ī��[�l�aڛ��ڴ��L#Ԇ�[s��aV,x��bjU:�`��ƌ�:,d�l��f<i��h��D�����M��=�� ������W�z�G�? Ư�d-0��f�Y=Dsm��3R*�.�*z��y|��{ʿ�
K�t���I5@ ���S���?k��sO��qg�ae�sd\D��M���S�_$p��8**i< (A{%U4��HJ�adۢ�svY��޷�$!�4\>]�}A�>�p(�]����L���u����B�D([F��h|m���l"�����~�a�1�K�����!��"$8 }�Ȣ~`�&Q]���o�X����L|+�o~�|m�fV���g��/��O�C�<1f�e��J�6��&��U�Ba�,�=��솖�j9��mƗ��k�8j�Q�O�!S]F([�|�$S�����$�݄gAW=})��!���������Qs�u��:LM�B������<U�����p��鶔x�ȯά��X�y���B�;V�_�p��&~L�/��b�~�{�ԁ����cO׊P� �y����d�86�_�u�U�f���S�Bk
g<�ʂ�_M���l��u6=��ZjX��e����o���:!�wƆ0@�Y�Y.�W^P�V^��v��EmOÇ>(	E����Pŏ{z[���ے-bJ��Er� N����ȭf�LV�#%�P�˅$e���З�P8�xt�iu�c*Y{�QnK��E��%�t��c�.[�[Ak���_�"L�0�y�Th8�8��}�[Ķ���/]rr�dSڋ��\ăQr}`��:m|ҝ h�m��ο�#:��_(�h�����@I��_�R�f>|�z#��*]�
9��D��?tXM�;���w[kh�L_|Ǣz~:x�~�����L�۸�B����"��S���L/7��e� �ۭ� ��2Q2S������ ܘұ��4�(�y�(V��ǈ&Т�H�t7��� 0����Ԛ�����x��[n]T��(y�p�ƨ�1���4~�ILn�n\���|�p*����ڐ��&'m*��l��7N5�:���<�J�䐎�DjAA����9{���,��|D���7n:������L�SoUE�ݫ?�a�ۨԵC��C��-�I����u��`���z�MwI�ڭ��zf�M9� �ZqA_�E"8�3�]-�  �i�� q���(>���H�j�W��C>�u	�� ����a��?����=>��Ǐ�~��838%�e��6ś̫�����v�I�UO���.N��@�H!��=��R��՜��1�]�y�۠���n�Rp��G�����y�[�#�'�
w��k˃+�w�����o��TO@�S<�e�~��̾������S֫y���g�E�R�������!��he�1y+ǰ����4R�OW��g��:z�
�>�~��!���zQf�R��>�u�c�.�F���z����ʅI���W�Z�=N �R�/�#rx6_�i�e��`NY�����~K���^�5��/uk����^}�š�u"��#:�}��y�;�����`[��#��~'�Y,|$�_P��%�LXO����Cr��i�1R���������޶������X���ӵ��AQ�<��(B����&�S�*�����(;��gX]��Wy%��>������
 d��kܵc��`�^2�� 8:�Hq���-��pD�ښD,�D��!���q�p�+k�r��?Vk�J�V�2�� NvK.�Y�v+��xs�A��ҠO$vT�ֳ �"��I=��
7in;�6���ű�IuWk���ϷK��'���^�Ϥ�Υ�Sor�J��OP�}`�Z�8���e!S�srKƹ�0]��L,Ys���.�lX����1�z3��f���/o?���O,������F����-x��3���T�k@��3�K�#��J� ���7G�n�(�\���"�*�(��[k01��J@�Fe��or񔉣.�+7��G��lW���KQ���5�!J͒���p���2s�����o,�ߨ�.�*��D8y���MNk瘬>��K�8��7 ��\�I��Q���޾5��,�>F���e�Xz}�|忷,F�i,� 颫X=�MI�Gdu~�����btC뾺؏����W1�^n
������?�_��h�f���^���G���(�̬J����
��A��ٻ����rT)k�{m����B�EMuY�����OX�U����jV�
u9W�s7(z��:gط�(��_��ڭ԰y��js$�t&_� y,���`e��Z�l��,�]k��i���\��1�^X�;��)}C�ld)=�|J�v-e$��ȼE�H�'cz^!8�
]⎼��9.����7�Syk����pn~�!�efG��:Z}[F}���O�-B�	�Λ��F-uc�soP(�]Cu@�c�m�ed�ޖ���bOP���E�M1��_�Ͻ�Ү��7+�3��/���f<�o6V���Qi&�7n��|��I`���h'���Ly�K��Wdp	�9*n'�2�o���슣�9��㝤8|���~��$n������-Dg�~umea�f�:7]�����.l�,����s%���w�P�|�a=�����K�p�W�mh^zv��j�� �OK7��[ь�Q{Q'eJ��'K��-�[��P�a�#�b��=��
��"��ml�	S�Cv�Jn�9kZ�rQ׎lZ8�D��[q��x��Z�L=p
8i�K��A���A���U��@g�����u����(�V��?��I��{:ϥ�+d��+_�:���GqK����uV��k�N���&�v�s�&~iM��Ê&~a����i)t[!|�C�7G�b��?�ٱ���oӴ��T��X4�a>��:3װ�'���*0�u;q|���4d�UQ��FE�2󋐏޻����k�D�� V�V3�����VWj�\��rCH�hT�������zs����z���ܼ��?*�!����Kù_&�zY;�{/����`A�W�x\{�Xx|Tݕ�ƾ[�Ҋr� /Z
�~4&N:ж�Q;x���8��9n�TI��o=�5R ˖�<O���8�7�*���w���i\��׭r\Wc@є7��굪K�5e�
=K�	��Ƚ�{��4o��q������_�p���az�H�?���z3���}m�W�{-,LN��9�.-+%�N�0�J���Z��XM�I*�K��x�ןXul��W���1+�\���.�s�EZN:���@��z�F�4�8H�����	� k8�Q� �Q�M���1��/���Eu��6Rk�mr�{��)�璮��"��]��Y���=3ȩ���ě�6����2g��;��u(z����H�q��?޸��k��g�5a�m���Պ2T\������{��^8��n�\�~
�yu�*UXamgË~T�J����s<�� õO)ii;��H�;�|�}���E�&o�����Q|������_[�>��F����g?
ȝ5�!�������N�n0t�4���<2T9й��}� 3��/�����a�&c\`�v��
r�5Eܙ����¢vt֮(/��_�/���)B �Ȕ#M��W��PY��D�}�~O�Uv_�HQA#TX��]�d&����Q{��J|h[V��j�����M돩���-nkr[�Xv����Q�8\�Tư�?����;��+(I��Q��('M�6�2L�Iˎ�C}A���	�B'C�C���S"�ϑ�!��`Si�^h(S2�B�����cc�n&�,SUomN��}=o�V�VĻte���%�Z2gn�gL��뗐Ǌ���|q�!މ����f�$q`�a�O�<=���߸�z�~�
�/"�;5x[J��@*@��EV�7���g����V �A3�t�{�i�vΌ��@_�FE�D#�ij��^s"Lj�CH�MJZ�ҕ��:2kg�R�,��Ղ�|�l>�X�%ʬ�þ_�?��Ď]�	��9�dd�U!���z��x�S�y�WB���f*�:j�MY���+,O��Ż)��������U�:�̃s�<� �V��W����*����X�ˬMN�T�e���'�z�X�4_���t�=�;��i=�0����?[Q+�O��`ˣ%ue��N���%&:�#��.�����c�^��@��Ʊ�2�5����ƣ�<0�~�aM�s�*��k�8����**�v�O�m���-a�*ۤk�\" '#P��2ꖐ>#���L�ĔY
z�:��\s��+>u��Y�}C��)��u��F�Ds�$ 7Jw"7�~�3����OFs�a`5���岕o��kM�N���c�Uj��CV�	�N�ڮE\�u�m긹� �wlC���jSС�.�T��1S[f	z3|���{hY���p�lez慽2&~Z�F�4��u	���N"R]��@����0����AOY�ӵL�ڗ�E1;ĵ�jp��9h��E	<c<:����n�U���t�3�&�uh�4�Ǒ��I �XLW��-`��]�]��q�.F���I(#���nZM*
L2(��\H��e���\��T�W���R�@��ґ�C�o>3��a��2?a��^��@\���qI��ޑk�Bb_-�ϓf��C!45�ę���?$�w�!.�����ZV�����S�~���h�:�����V+��pnr��w��D���%T�ĕ���^��oXf�]Pm­�ً/:zQ"XbAeD��+M��?�]</�FP���F�UI���dn�!���a��H��P��)C�\I��'� hʦ=�o�:�1���f�'�P��Z��P�+���0I
�^P�}�فgǆ�׸����Q���k�J�/�plJdei�
boF��k����%0�l����O�Ջ���Z�W��͝����8�t���)�U
I�L<�F) �]D.�
�i=���[5�3Z�rS��e�}�Y���EFoW��߽��]��
��]Y&Y?u��6�6�����ejڷ�]�)�::��C~�F�bb��|�֐"�G�8}30B�9�qyA'aBc�n��}V��R�8/¼e�f1���y���٪S��r (�G�D1x�YL㖕	�[�q��D�l?�q���)Ԗ�LyO75L�􂷋f']�@ą{��8\	�T�?_�QhX�W<~��y�ɒ�Sa�P a`�"�^���g�q�:�4BD�W�n+ �iO��_3��˥�Fqe����l�-4}y��	���7m��har�U*���-�t��׸��^7x�v�z��kḝ���G��9�0�-	]X��_��k��7���I����&�-{�n�@\< ]��u�L�槷!eo��! ��9�,��sgǕ���$Kt_xɖ�LY}a���_�S��4f�V�a��|��S���L��:gR�����o��9��Z���7���4g�H�Q�<�@����i���ۡ��y����%��ʟJ������^�'�&Wu����bi�ZO�#�?cՆ�%|����q�Fش���m���|��b1J����z>�&��F�p��Iz+"�����*Ƒ��M��w�s]e�#��篜
g�&�(V̲
ց<v���I:"J<�u�p���=a9,�~&aK<v �;ovy�>��x�>���_�QB��}籋���u�<���,(~d����mo{5��h�Y�F��\[͝�bz��o�ޖ��W������e7�h��Ƀ�Hq�K:�xX�B�������V�Q.�6n�>�X�Ro��O�����~�"p�w��ӎ�e��7мxoPfȱ!+��`�i�:��R�Ffє�Pw^�z�&������!Ċ7��e��~]߸rd1��2T羆����$g��ߘ7��N�ǋ���Ig֍��U�q���-�Pz�m�V��!�� ���b����	�P8�P���BgAȷh�7�Xc7䢝r8[�������/Xi�5�?�cksK�h��^�RXM����`�����|x��7�4�,�n�0N�c6iv��n�<H�ֵ�����Y�΀�.b*7���q���bJ��i��b�Xu�h��ޭK}�B�&����0�~a���`��NE/���O�_c����tf��x�(/���`������X(�h����@�Ճܰ�9*h���?ʚǍ/IaW�{�㡆.�k�"Y,��ڦ��v:7�$	]md�Ue(���̲��i�Շ���=qq��V�I����z�gX��KXnpF"��iC5�q��ߖc��Q�^��z^6'��.u����9/1L�Uw$H����I@�BÈZzz�b�c'S#�d�r�Zd�0L%��m�b���o��K��i��[�� #m2���u��f�D�޷��j������?��`F@��h�]�_P�f
��ܔ&Nj���������;"����,t,�DI'�~��LRѬ�AG��+.��3���'m��� ��aǔ����7`��p6~N��(u��8"Էa��U�/���t�j�e�n���k0�r0�j�ю+�O�h���ᑞi)��������xہ :�{�ޫy\�W�#E;J��72h;��Զ��갳�lz:�w�ڦ��U�P\��Z�m0V�b��D9�0��d�+�T�H�Zi9��~za9�4g�F]ٴb����F�1,�uFVc�a_�Z�[��>`��gE��&�I�z�}g�D����k��O��&��j��=�W���1�aps��lwW�@�k�m5�W��9��:�r��ׁ^�v�c��GQA% ���u�nZ��(c�ܷ�����=o�a�u�į��KHC�b�D��C�Z��u8M��	֘��V���a��T�{�=7ѳ�Ҏ�֑�r���6H�{����������oD�Hq������T�2U�2;8	J������]��eLq��� E�Gm��h ��=f����ʪ�Q[��*��Զy	�><������u}��7�(��~��x_�0c�
7݃�-4L%�Zs����UH��=�ʫQ�{`�4�΍�V'ں8P��(���[��/�BF<��E�׬
0:"&4L� yp��ݶ���������v��fj�C�,)
U�/^��zu~��~��l�l#��ֆU�t��ӉE�ާmgY�"FNrL��vE�����LS��O�uE���\�ﮗ��f%LW(�(<e��OV1�܋���
��?�W���]TC�e��
�T�"=9���@��j��x��<<7XǬ"'�f�LVk7��5�W{���&�������t��cGU��if�8k,j6�DwY2��Un����o@��U	TLF�
��S���Y���=��+�x3��a���7F�Q#��qcC���鍨{�i�un֩&8�b1I�*	#��fG/Ե;�����A�i����G�W�7���K���X�ޮ=�*���Q����ͽ���q�ѱ�`�u��٨-�e�#�w��,[=Պt7p)��u���-</߷că�4��B?�Lr�/��ˁ|}qQ�,/���im4�f�k�9���Y�'�K�՞1v���$"��eK(C;����.Cy�4��ѦP��C�)�_m����]�t/8a�]C�i�h�d�����w�����,�к�Ul\���cKYY��MR����fɊ��Q����]�z�"k�ז[��V��ye��ZW)�W�?�ܥ:����;��˒��L�9���Q��A\����KѥnϾ�+��C�B�(���4p>NݲƆa'��M�4h;��M<��#� @�)DI�$ɠ��8�"�2��$Ϙ�Äux�,Ω�n+�̿�]�Ą�T[�$�������#_�)�򂾼6
!~.��A�|\�j�K�����B�{�[�BOi�Y��_�<h}�ϫub��]bPG�������t�xJ��a�����M�^Q����E�����(�I4&bB�#F�#"�gS3F�U�ތU?����(�[��a��l�H��T�T6�8j|������Վ3ޱcwlR��vDk���bC1'�w��5�8"0#�:e/7݇}�qu�+��Z���^~6���Ҁ��.kS�C�%��wʕ"��l��b~}�#��st3��ם�E���5�&â{��2v�ѠHj���@x�]��]m~��#�b�PlּXnJ��9�2x�\�>�89f�u�p���Ywi7�3z�2��i#���"�Sni���n��UO�e����:!��6vΕ�ՊP~����j��Vm1NKq՗9��v4���jb��~�� ����G�"�ܼ抴�:}������6:��e'�a��U]~�>�c�m������Q�qI}|�+�|��ӥ�����;4P��Ɲҧ��x����]��C3��b7�.���d_ms���ׇѱH�\�?ŗ�V1{�ו��S\S�J'^�A�O^���?N<�'4]��^����t����y	)��*�JJ�ŰC�U~�w,�����bn�qu�L�k�#��o
x��pd�y�b,����#N�z���b�Ő
ҙ�bV��p�}�A�j��¥\�2`�#-��1�k��]������PnzAV�"}|>x�hО��1+�;@���I��Qгbx|`��V���"i�M7����Dl��af�!�����o/�F���<�b��B]&�`�%���S�]ͧ<4��P��=���굧�SP����������T}�d�mu�U�!����2���JM��M{2��d��7VM0%���"��߈�����Yƃ��Y���C=Ly{�
6��e��\��OǪ/oVb�+r+2U&̤j�ny��M`E�"0�#a���E>����8�!]�(��Skk�S�����y{v[�nL�b>���G��p���PԇVN�\��R�Iڥ�)n�ywQ�(�E��/3���r��ԣ���IK�Bp��P1��̉5G�&�W��>� ���v�<�#M��qe���֡5��]�u.�n���{���̥pM�|�_��8_������d��ޭ�<���`+��b
O����2� ��ELci�sK��Ǣ�>*(�L����bUoJ%n����rk�M��Q�*���Z��v׉�ZEq4���[;�L��3�ȇ��D�&~�O��}g�[)z�q]#J�?o��;���E&e�h�]R�AΥ���5C�ʮq�5iW�-�J.�ۓ��w��>J�e���]�5����:~�!����ch����\�1�a�	��Wsy�Qb)������#D߸�O�\�z��Af�U��#�|���D���[�
�2���w���yj��t��&t$��t���K^À1x��-Wg('^�hB��{�e#p5!'������ˠ0t��J)��G��.�קh��tL�{]��[�G�Q/�m��N~�Yj�1;��W\�}����w��*��(��d������V�����qJAĢ�KHRhp���")�P�Ɣdߩ2����	������CX�8��F�+��Чg�l�L�#x?�)����$m����ۃ�0���7����d��F�W�w�GK�BB�c��3"],B���?��^�-�*��q֓��I-E�/�i�Wf}���.���fU�K�Ci1����Nk�c�s�Q����7�4|���j4=❎}��\&Ma)�g����q'�o��'�t��f�Y������k8��8:P�o��>�����7�O3xl�>V�,�m���<:{5�瞱�Y���Z���ր��uҾ�������#�O:��wb�n�vr@$K[!nCjⰚZ���~��ҍ��d%�>��!��E�1�����Z����z����6z�qb�G���E�/���Ӑ��!=(���p_iwG
k�����B�V(ic�B�����䪡�Ӎt��J�=�8��-�C��Οu������{Z��Q�mr�&(���*�h�k�ϒ}W�>����+��F&IY{}�2���-ȧ3b��ό��vߛ�ˋx�R֭�A���xv����ydb�hପ�Zm6w��x�Ni��pXV�ds��Q�������f����=�6�2�O��I͛x'm�ɵ��ФQ!?gY����C2I�Lc\Q��n��������H�D�N��I`�����)��ɖQı��^��:����������=C�}�3}Z�4�U�=:���E*�)�h@�d����B��M.��:7R��#���5)LcS��r���'�v�7�AaJFm�+\�}ZH�G�%ڼ�Ą"���k�X�˜{&�y�3��q����m��@����Oʻ��r�+_�?����q�o�K��m�F�1���
l��U��5�hoX�l	}�SvJHꪉ_P	������:({�xy��8/����gؼ2P|rEg>.�[����g@��|�M�W�/?�����<ѐ������RT����"<^4��K���7?���I��cwdJ8C�������(������+ �e�h��8�/!v����XΟ�O���ЉK��\J��u}���4���4V�s�q[ �DT'�x����S{���L��8�J e�*�rzP�Gts1V5&}��̹������`ľ�vLgt�: L>��mr���[Fng��@S���be�_
�:y��*��~>�aǕ�������ʒ����"�aC)9����e�e��1oE�dݱ����A��Z%��״R�}�zk?�><Q]�.����XX"&;D����|��ϟ�=1v�߭�+P�&��9b��v�k���א��n\�����5?�Sz�\ƍ/e@A��S��z���p�=}��YtRۃR<�� weu�xx�bqg6�D�7Yx7�3�73��w>C�|�q��zG��Qq�����Ka�-��Ex�s��OQNH�X���eGm2����x5L ���]6/R�}m)l55K�'�9��{�T��$-3���W�jQϓ_ݗ�p�vD����h����z�J� �7�i���㼤�6��
i�f�I����V����Z�$OFW�s͙}��=�旝Ϭps}�[��ɴ&U����߱�Q���'w���T�J�o<���d�M�C�rv>�Ə��OȾ�A�C�A�n( <J-�?,]��1SF&z @�*�����&�%5�;I��.��I��8�?;Iպv �:���M�n��]�w�s�|�d�`6�a���o�G��}oR7o8��
+�������|��/xK���M?�7�*=�;���5�ۥ������s���<��S��Q�S�w�Q��ַ�1(�\3����BbLǛ7�`@��@*w��k�X��(���W�����^2��`ү�~8!ߛ{�2ZBԊ{�m��{I7�u�%���.T&��Ҷ��|I`g�� yA5�(�#��A �F@��F0�U*L9z^W�AAo����\�`�6Q����#��(؞g��ǌhe�jk� .3��m�
C�]\���KGg8�'��j���^���o+^�da�8�?<~�=v`����g��PRHP�����wj�>+��-��EXh�ߝ�ED���q]Iյ�@�,�5��7U'�Ɏ+^��挄ܫŊ�۸!��Xx|> �U��F�"`�\��.j���Z�L�e��(�R�{���g������F�C6������A×���??H��2�[Ot.S����dv̅p\b�t�����ؒ!��=n[��%���'/�@��֯dDZ-[��cp�~iD���1B��L������~S}ꚟ� E���q�m:rl�MÁ'�ˌ������]��rr\�|8�48���ƻ;��[�|V���=��H�����Ƞ��!��ԣCv�%1��g�=.	�����I�V/Y�ʗP2v}��X#@�Ӕ4Jh�ڿ�!���}���dt˴3]P�3�U�)qU�(�Sl�:�`	Fh�����17��|�.��D�l���ʄ��`H��F�D�>q��+K�Eu�+�u�?�4�X���1˻u�����߱p���b�iǵw�}YwO���wb��&�8xtΏ>���'�b���.>:Ĵ_��̺{;$[}߻ZS�����_O]���g��;��~x��v��/�[����+�����hͣ��F����Z/���yyq��W������H��r������_7������Kx��<H����e�SB PK   ���X���l��  � /   images/30131ebf-3f05-42a3-9ad5-e2b3b9511573.jpg��TM�.��dA@�0*(H�q@$���"�%�8
J/ A���sCFr�0�&������s�:�{oM�Z�]�U{�޵�gw�7n��JQE    �� n�o��{�� �ELLDDLFBr�999%�mJ**r���i�����SP߽�@w�����o'��g��I��I�(�)��?\;@s� M����p����� �� ������W!����&�-R2r|����B�D������"bڇr7�hZ�<r�{�)��-���Z�G��܂I���c���	�S.!aQ1q	��
�J�*��ut���,�[Y���ٻ{xzy����|��5"!��o�i�9�y��Eſ��kj��;��{z��'&��gf�ͯ���llnm��"�ON��/P�W�" 	���/����u������^7��6�!"~(p�VN����Σ�nѽ��Q�A�&�uD��m���]h�1�j�j��N���_��ߊ�?z����GH�̛�½�%hة������_5QC<߶��㰿�H��н�nc'/�:���S�J[�q��<I�2�Y��P&》�k�jM3��Z�Η��$�#{QLU+M>x��3���5w�Ba�mPmx� �1����2ɯ��[�WB��w����@8�2�(V������T�Јj�+����@�u�kۀGf�\�XL�3Z�I3��{mm[E��h[A�x�%Ǌ4jkBP�M��q��k����14��"��Y�/���*�]@��H���;�y:�/"�;�=G���_�p�#���5vT
�@�#��!�PR�8�^T����hz�������g���)�s��(N��@^�q���JRi��8�Ms�
#�dk�3EEq�T�������{�%�Lՙ������h�,��`n�ę0jZȁ{wS��s�~�A�ǛK8��&3�u���+S��먪7-�?�R_��L�
(OF�",�Z-6�V`���p����%#�Iٽ`�N.];�O+:ʨ��*XN��}'߾ra�j��V�z@�����!?��k�j����Q�,Z:��G��T�n�NA�Q�!e:���(��j?�Bƞ��]��3@�.�up@pn���F�<��RM�T�o��+�/K_9��V��?�0w>��ǄU�&Pc�l�Z;�z�N�3��.��`��O��s�{��h��ʤ��ړ?��v�E��h�d����,��{<ό�4;+�Q��2ɱ��0�R[�2��0#@���|F�n��y��q��H}B�uS��d9��L,�_�%F��`��|E�L9����Y'AT:�0	���Ձ�8�����!<)�E�w��l����S&�	
)�2�8`�����T[{ܳ�3����W\�=Bө��5H���N�؏���q��'m�2�K��f��۱L_^@�CLjˎ��k�"�϶�1����e����6�ex}D���va�'�Tn��Y�eB�n�x�HήƆB�4�*$k�s�]ݹ{I��:V9H��.C: �E9;a�tg���ܔ!�����M�3�@�κ;��������_�M����WXe��~s�v��F� �!/s��n��șz�{[�T�oR��VK~*
*�z�� �wJ�Z_z���\É!-�����a�Z8p��I���츉�k�zT�8o�w�h� >��F�*%��%5���<��26#�?*�q@{?�M�2��m�	��s02{�/�<�O��V�~E�M��5��$u���aZ��B���3�&P4o1dl6���� Ű$���� �+|3e1����']B*�A�`d���i�G�?�dFl��0�{$�p@�o�4�(#3*i)�\�u ~`�̅������R���X��R�ʭx��>�����4Dk�����c�[����:J�@�$����aG���~��ۙ�\p]�z����F�i\1
U�)�3Vvv�
�`�o��W`տ�P>�a���y�f��G5�O8���ՏdHV��cs5	Y{�c����)8�S<�ƿ<!=� ٣N8�����;���/����� (F
m����O�LE��a�J�m�� y>��O}���ZU�Õ�J��ZI-�N�E��w�-����������|/��RR���U��f��G?Yf�YA)ʐ24+˿����E�Ku�u��
q��
V�鸆��y,u���q���?���$J��N�Nv��=�uĭ��3��.^�MC���_w'v<�֞��}�?�>=�
��ivu��{L��4s��S!�i���|m��d,-k�&4Դ�q�B'$tog~z�m�o���8�(nG)���h�� n�pK��py��Q�3_^ț�4^�Ww�v{��#�������I����w6�E���bW�k=�߮�����1�<�1�n�\�e\��_�ք��̬*����j�>�.��21�<^�'T}X-��Ֆ��*G4"(*K���yg�P����ӆ.�b����yr_�Y�Z�[�-dX�(�Q��Χ����,��AH3->����#�T�{�:$c��h;�]�����
�}H��݄�{�J�bD>ذg��4��M3�%D�[�ZCB��4m&����zǕ$���4�{-z�G�C��
"��=�O9(�ɋG���{����(��t.��$�^������_�6�^W5o69�_SJ,�^�tTvD�2��j�#�[f�_��3-{�bzZ&J�`���(+�gث�X��)8N+��e����T}�襠�;�FQM�^��R��+�Ӟ�H�&���7�-9[W3�h�1��hK�<���dQ��Iи�R��1Dj���緫�S�Xl����@b�^^./���|�fI����������j��$B�7�Sԉ�C�EBs&�]��S&/렌�wm���4�0�úϫ�iqx3�zV��>_w���5�M"���ٛ]8��NxFG�z��͡����P�O��!A������+֛#Z���!w��8��Rt��+c�����M�+�p�׷Pc�=���նG��B���P�іo*�m�C��*SCy���g���MrC�O��=9v�S��L>Ygfyt��uY��Y�2�&�VyF\-a�).�g�e>�ًϔ�{��a�6;}�'o�̓��hݵ-�j��xŦo��y�������/A�H"[�֗�0Y�]�/�3x�X���d�[y#f�o�jR^�
%�#���������$�p�:atG���W}kT���Bg��h��Z.���9_y'-��9��5Y��3�O瓇鯛m�l��U;+'��ג�Dv������W��U�Rޟ����8����Vw�hQ�Pq�rJTSD�\�B&;����K	�Ǔ�/s���:	�����)^�T�Pҗ���M}��uQ�ހW�T�#�����雿�zQAd�B��U�P0��Kc-�+0h��9���U'Uh{��e�������y篠�eǌwp@�!5�2���/G"�(O�ըQ�
.����C)����oų�H��!!�HN��ؠ�D�5�?��7t�˔Cz�*
A���J`��p��:�1�E����*�q�Y�ˣ7�'�9Sf�, ��I{�֕�<����X_6�kr�6�����;�c��[����҅���\�Z�x�|��k�[���M&�=k(��P��T
�_�.{�&��z����Tț�3�<�ݯ�5�QZ%�0�,��BBD;d�:;�������j��?���.Ա.D$�u����f�",z�b_D��9ѵz;�;�qx>r�H��S//��3���Ƚ_����z��Z} 3�sS���<��}�VyEP9�,��ں��S��wwe!U�dx�6u�1t?X�v�G^��B�&�QO̵6���3UGB���"����Τ�c��mMm�b1fEA���C��G��s��\��ܴ��Kx�F�C���=l�ⴧ��!o��-^��ܒ�Sg�Ұ��tֆ��n`g. �m"Pd�H��t�S�"�A�8kAq�Zq���V���Ve�9���������S�̛���j�kg����]2D�EZ*\�4��jI���հ�aP��AT��7�V�B7x�~p�
�RK~���	\[��[�qx�c�,B��܋�/{���8��Y�4��t%��4�/��I���ɳ���\��V�k!����3L�3�wp�3�+)�2�G�a��?8 6.��D\�����!��ʽ����L�Yz�ù����L�ԜL��	��blh��W��X�6'��|��&�ýy��NS�Fg�����;���[�f�/��z���Y#c�f8��n���6{�w��67���ʄ�3�)�:�&��]���\լ�c��:?�X�q�u� &H�+D��m�W5�O3m��)GN]�`�Y���b?�-[U����4�O1��V_�y�BQ]0ⴂڇoR#�!�{`VruJ����{#��vw�0�m�z��d@;��O�OXՔ�n��̽f>�Y�O��p
��Q/���k׳,j�)����p��KW�嶉�n���A�/q!q�`��ɦ�
��M�4��aH�lyq@����8(H�]������>���:uSs�Q�?&����R1�M�S��,���$aՐ��f5���e�:�"8�c���C.ʌ=�6xr��t��kZ��HC��/��91�m�%��>Z�_�k��-���YŰ#7,:���{�LVZ!(�!��dO3����1w�_�,v�{�hy6�>������U+��z�m&��m�5��[�rx1��1W];_�g�!��J:�A�Y��{l�v��2B���Ӯ��{��O�֪uB|K�GC�?�81�mL���� �?sP�E�l�R(s&��"��Z,�F\'���M��Q3j2��R��K^$��("'���m˯����?a�<����,n幓8"���5��oL�*�̓Q�U��@� 7Ֆ|�!Q~6�}u@<�@�IQ��jw�4���;�U��(���6�\a[:7�EY�'���M��D�q�fQ������{[]���]#�P8�.��<��#k�m*R�q1�o]M%��6έr)����r�8-�{�5�u�fݲ�tݻ ]���zl�qO���Qˁo픨p�̧����������	>}�v��̞<9G�{ʕ����������W$�	�ؤp�^�mZ�l����_�K
�v-�-)o:�����_��M���d�� ��WH*h��w��"����#>"9��j"$q����p��ӎo^<J���E3{?����s���J�e�ڛ�8�P���%T_F�O�(f�[3�[��N�j�i䝮�pcUZ3u�y�C6�S8Op"�j�Y��'+����"�-C)E���í���@@�����~�~i�SorOڍ�x���6�9����w	%�a�ho�^�Y�Ҷ(�����������xژ�O����Kr�W��k�
LK�I�@]�h��
��q��+�_cD�y���_Y�Fh6_## ]��C�����P�)��q*�+OwAy���M[ �E"7f�<����݈��	���!Fg�J�YUBX��ʳ�DYä��5�@��i�@��y��q��"��^�w�����mGCGj�J'�I�'�����O��/��v������f�-��-jD�X�������q���/�N}���]�h��teL|bY���7-�^�S�Q���n\e�]s?˵��;Q1��x��o,���&,�'��h��GZ ���Ι��ڏ��4q�%*-�r�TP����ؤA!�e�P�w�$���@�Ԝ����Km�3�̦.�=LߍK�<q���Ӣ���s�,Ov����o!=��_z'���Ro�3��I�Ͳ�K���|&�'�kX[8Q�U�Q�Pc]�����6��ZǷW�P�\����Sd����.�����_�S��c�:�����c��	�nV��I#,{���1����P�f�cX���t߱d��+��فVΙ�3B�t��Iw!�<C� ��QV��<�GA���d,$$����G� �w��Xі�_�,Yd�?\�;6�gL뷄�!���j���#K����CbRa������
�%)#[��<���+���&'i�#��ô��-����t</o^	�jfy)������7[�#��2�f=����K���08(4�F��e��J���%r�'�#ܡc՚
�d����8.�?����J��(��f��B�>�Ͳ�����%0��i���"ӟv0P�{���L�'}c�㣂��-j�c��˳�|����Sj�ԭ�b���(:Vg�� 1 {�E����}^�Ձ��ɩ���
1T'�6> (S�ԗ�3���{띄c��F��g�ʣ��<?�ƅ�ʪ�lr0�@��$�tO+޸|�ws���{Y�nL3�K�e�RtۏrH��ԉԐ?u"�ͷ����=�@�^��*q<k�@��,��&�6��$y֥�:�C����I�WΩ�������5)��-!.(q�
5��6��|&�h�M�$,��T�e��?o��	��'>p�6�P��7�߶*�mD����I�_1낏[F����g����"���}w:�^J�Ԍq��{�M�c���R�����6<���^a��Kp�DD�Xf�I/�~w�*�5����	p@����L+�Q~k4k�`�'������[8��֕~7�Hk�IqM)=S ��z��Ë�*lm��É'��<ZA�G,
��"o���N���ġ^u��k%��b�#��/��'���,)>	��S�;c���f?|᤹a�_� ��-���W��QؤI�Kّ����wP���������[-&�w�i�f��a4O��u%;a�c�:ڶ,6"h��e��S;L��(�Gm���'��X�����Y�;e���ou\!멻/�	,IB-���JQϷ��~D���A"Ly�3�V���Px �Q���A�d�������s�DMٝ���J��>�&1�2Xے���bڰO��#A�鯿��
����mdõ��[sVM��ܜ�N}�e�ٙH_�p�DK����!|4�o��)� ��H�<>��!�b�>��l����V2�J�N�c�R8�/t3����x��Bt-I<8���U7����x����>��b�'ߟ5��R���^���:�e���;��2��� �&�5��T��W`[�Żނe��Ѕ4yWּ���½8A�J ��F-�����]|��z}!��?݆Rv���h�i�k��@�*�������)�%-� �gl;�4��Uq+;}e��c�r;WY�ʵ���7�6V��TR����>�c��2O[#�n``:|@��LW'(9�Gڱ5N�a�Ē�� 2��(�>r� ��6?��F�!�B�p�L�9���!�y�7��M� )}~�"�� O�;�gޖW��/ǖm�]m�����fb6���u�� ���G��9��q��+��4��~�*�
&���W1M�R�����ub��־f�b�"�|s�3pZF.�hkI߬h����~��s]�0M5��W��ޣo�Qq��1l���oƝ�/)����oх���x/��b{?ya��>XΗ�s%�̡�����s��r�S�G�qJ�˯�U^�;����`���Xͫ��X��1��_u4p���V�Y��Y�%*�}�YS&G��E���HC?�Y�n�ծ;jr�m�xc{1f������)F�Q�df�p���{�>%�T2��'xA�Nk�����YQ-��&�r_{���_=�Ө����E`�͏h��xz�F�=Q��e��}Z���B�೦tņ�q���[R��4j���O*��E~�=N�]pq�=�]�?�gм�RF�gK�	���<ݓ#�G�#y��c�,��72"��<��XXj(E6���	]Y�T`�X��V&$�2o��LY���Ã 	[�t�Fl,��3��A_�!K���� ~{`�t?��񚇡��$SO��乴F���?����~��a�3��
P�;����!���s�ݓ	�-3�_]K��81���7~�M^�y���:IG�<���tJ.��P�P�I<-*of+������9�2�1�u�����J���v*�M��I_Q̤�`%M��"�Hߥt�9Q[.d�\�!�b�9 s���y�oX��A�ο!dX��p'�J��W��17U�z�U���jᨷ���shU�R�
2���Z����I�e�����#>}f�2���#�9f֤)y>K���1��so�r�l�wzן�֬�E���GH�H�n�=�->��CK��| ���i��7�o)��$�����3���"8i���-�+�kn*�n�3�����E��?S�b^_09$�8��O���|��uXgjJ!�~���7��ø��-��{s���;Ы� �W��܊A)2R�bf�lI��#���tH/��ҟ[�����v�.߯j��5_�s�-`֯��a@�n�m�����~������%��� K���� �X�w�����m>�h{`�A���������a�M:rt���Fd����c�/-��LG@4�_�N�S�SeioSl��봑q�%)&~Q���vX��$���
Ǥ����	�����c�~�O��oݮ3��*~���-jh`�}�����v1Gp��e�̢���v�]��f/���'t^���_l���N�,Z�:��&��gF�w�`���s�I�|-���@��v+���.��25�"#m��Kڇ>g�a/�{<�~5��-ճ]i_��Z"�A�C�}�`��)�7^i�8���coj���߻����<'J���,�����|N��Tk�騼�����@��ɕu�W���W�[)��z�����gOIϚ����{�x��R|=�M��r�b,Հ<Z9���Sٗ�y~���j�	�Ҏ�T`��v����dvGw:�r��(�3+<V�<p.���L[f�����H�6d�Xʾ���A/�#v0�<���;���w5��\D��f��N���X8E�@�!��ИL���4�������U��,��E���V߰��c94>d��e�Ljh�Ʈ��y�[BT?�9���[}[�j���4W�/����_��Y��w���w\��Z���ٳ#^g[/���.R��46����m�e5�����fU�`�wT���*��AH��y%���5�J¤s�g�1�] �VI�M�����{_㻟�[o>�1�MьS�����2Q�
�~n/�|��j�x�eX[yP�uZPO��u����ە���|���o8�<gN�GM:���ԡHa����XDb�#�n�����a`nL_��\���6{|�@l:�6�]0�녺��Z���:I%}�^�{-bD�!:+��O�� ~�t50\�� أ-�&�u?���mf��@ϟ�ߟ]Gs��搞���ݚ��ČUj~��֧���|�!m�P1�_���su���J�<�d�q��ɉ�!�K��PVd��)��B�',/ ���<���IgR;�}��j�o��C7����W*�/dX'��[;��?���<ed�k��������'�j�4|s{����r����j���>��0�X��e&��ۺ�茄�1��������C*�b���ߎ9�g����/H��_��� 價��W��G�e&�XZ���c���'�A�5ɵ�*��~�9e����;��wߟ�[FR����3���Џ
!�}�S�;2�k����Q𫩯��{�k_��J����5�X^C��~�){uQ��Y��{�?F�7����Oַ��G��3p�~�e��^���6�4	��t�7ٶmt!є��!�^e&G���8��tc+HMP�����q9�����}1Bf���W����4��+wLI�{�;�:��2M��[]�ԋ��/Y�9Sp�����)����
��1'�̫��l �V�=���<Æ��)W������u1[ce'������凭R�.��8;��^�q/I��-�I�r^�_Ɛ���ȍ��#c���<��ʛZ0���P������?�i�غ��5'��[��4-sO;4�$cn�6 G����m$�_�n$b��Jf-��.�󒷹�ҍg\�B�2��d�,e�����(��a�M���:m4a{��x-��/�j�H����4�-�^��y���%ڵ��Z�7���C�E��������!���>{S�DV�F���d���"�I#����`��j��Q%$>�s��LQ����~KUM0�3�Y�Ѳ��>�x�H��^?YU����Wg��"c����{|���zc��#c�`[�R����C���/:x��dB ���q���"��C�(FxY�'G�'P/��O��〽�qP����J�7�(ocY�`�!B���^~��</~E�*�����_�����b۴ �����6�{l����L�8t��}���J�4�*�p��+%����@�5��mJ��,hR��I��������\ ,I�F���A���~ڮ�zُK�"��AY�f�݈O�
�u�%��3S�f$t��˛9��7H�m�m�L͗��˹��m2σ��Y�zw����=��;�kݛjXmj����r�~;�q"]�?n8b��<�����Eߺgr.���mD}^,b�>�l �,�ɩ��OK5X=�.Ӽ��e�@�X�����5XC%�cn�{eL/%��:nY��u��VY���D��p��?�}N>d�/�e�|��Q���괙h�Zس���*����!B���M*��]�e�>��֒YCV[n�:8۲�,\��u��<+ܒ�����R���q����aK�72���Wm`q�V`t�;��������_}��u<��,���x��Z�ճq�������`VG��x�=~q��kr���:���f/��Oh�+?������8*ѫGyeҏ������1����N�R�����a��oE��j�!yc�x���k^��\j+�����|���Xɣa,���Eh��!�]�J=�܎�Is�������Paa�ݪm��K����?�#c� �I�ޢ���u��L��\p�{M����q	�9��5�^�imw%}1-�H�$�Qk��ur�8͢fq^RO��}��#����׈[�h�G�$�LcHˏ/�[Q��ɫ��-�,�J:�������ek��@����&��.%����S7���H)qR}�����Hh��!x���O</V�*qA�K��ͽ���sf�?k?Yq+\���^���3��*n��q����h.d��PGU�����<Vޕ<��Ij!s����i&�dB��5�Ŋ:qҁ{��ߍ�S�|Z�>\��Q�E�V4�˨Nع�2�3Y��:�L�A��&�]�����j�FTyG��������!�3��Ju����~�p�Lg�i�6�,'^b78ؽ��+
���$t�8�^��u�)]��#�A���ؑ7]Ϋ��X�w�!~�U��-@!2�Q���/3�hB���|��d=;7W:w1��ةS/7p\�^3���+�3��F=
��yh�VeM_�-%�*����M��T�t)�D?�C�� �P@r��1�>��dA��]��ӵ�5?�|��zd� c/����hY/����6>��a�+�$V9���H~x�����+��<\l�:�^���2}��kaU֐��N���?5����"j,فE�&�V*�j{N�LAG9������s-@_=N2,p@�ag��IS���qV?X/q��;\�@O�`Z�G�8 L��Z�[��!^�^�B�M�#�>K�bI~���`Gv����:Pň�DP�̍��S:ԪUo��]W�çz�F�V|�}_E����РҺAWv@)#&J��#9(~��n?�ʪDZer03 h�ñ�*�4|���ǵ���|Po+IUsĪ��2^$}����)����L�'8�+�qh���,�miJ��#6��x�L��(b��V�?9ؕ���Pd�e�	��a�īL_������-�fF2]�N�����]��ڍ8�?Jm�	u��@e?aV���I�F
��T�)rNq���̴}��_��!�O��FL5�oUt���(y�I���'��L�-jX~K�Q�R�϶^0b�T�M>ϯr�"H�|L�CE˵}O���F�Q�Ib^�����D�-[�q�n!��e��ءe�����7�{G�������RK�ߪ����֌&���{�h�u�:J��a.A�K"��{b�G�&�Ju��W�"���u�Q��S���c���}FY��u������Mf����[q1���\�����V607��>��R=�e*�7ߢ�
��_3��#�R2gi:��]�R�p�옉L,Xl�Y�e�,Af���O+�h�EӚ!'�hS�����y,ߔP�>Q&�d�f�
��X�L	Y'����ݙ�B�t��O�Rpv"�'��q�� j6��2���Q��e����F�t�Ok'q@%ܷ��tG�i��!xU޶O���x>�W֬2����GF?��z��.�d�>��~�t�ƻ�j�{����>�~}�ܮA��$||�}�w�|~��'���ɹ	V�S��2|XBY�{�"���ڏ�R5��*�`��?��Y���>>���1� �%�|_0rX�2�m4㮒k���3E93q/Ƶ&�J4kF��:S#��Ҳq���}6������t^����%�k�=�z�,Ϻ��9	���)��Ӗ7��$M�he�yK��"1= �~f���;�'��'��O�bi����7T�4��GI�d���O��K�k���	�[`9����� X���*��:�H�Pܿ��1�UŲ��:b��h4[
\h�e-�ì�/'=�J$rڦ�j4ΨT�(u�vi�Q]���H�J�7�����Q�/H��>��Ad��.M�5��Һ:�aY�b[G>�en�`�TDr�,0�7�]\�P�Ɠ�ݸk���-�=�%�]�ۓ�9���꟣�m�]B
��O!���-������%ä�̦�ӯ�n�8�n۹��"B9*�.H�t�>�t��L��-i5�H`ڈR-�a������
������&���{�~].6�(V�����G,v3�*SzW|,WꌲOD����wTؾ�Ċ#��3��a�R��$���	�
"r���p ����æX`�wo�na�N�����#jì���A����SIڮ�qp�8�p�p�����HR�����5��0��$}�\�ڿ-�vh�O���%y%ܜ�3�˫�.9*����׻�x��z��\�%����+�v]���S��rO�B�f>�vfk��Q�c_�+�2	ݸ��2z�������YE�V�Nes���ާ�	�F�ÓG�),����𚬵ٶ�Ikt���e)Rn�_Ҟ	����]+��4J��*~��(v/ԉ�+�7v,���2��u��3R(,S7��nJ�	�1�N�v��J��	�x�j˵���ݬ�.z�����|��x�����(�b�+sQM�c����gl��@�,����FW�$%+�2E��#�6�0Ԍ�2�;�sF���"r��n��=�H0�ߣ���g������?���H�g�_�0M._�<n�`�󇩊�OQ�q�3�*�,�hI[w����J�����{�W���C�i��KhE$�¡��)�+;����r�@S���"7l�{�����,%�7Y.p�n�/H���3[���?���<��8���{pQ���$��qpZ�jڲ������G�HP*��-�&��C�GxbaY�35�MV��>u΍�E\�ġP=��X������nm�}}\���V��|�$*-Y?��3J~Q�w(�PPe�螥贺%L���
}]wSn`TZ��vm2г��o�����,ST�^��__��y��%�>9���߁�����/�ŷ#�����=
��N�0�_�s�Z�c]z��r-��D�?��f�563⦹�iK�VN���9Z�7t՟]��p����+�3�Mi�S:�@:�ޟ�7�b��GJN�KNJ���D_�/��!8����Iߺ�!���y\1��bs���1��=$=���Úk�M�O���ta����q \�
��}4�;�va�kW�}���]�0�N;񺌢��
�����>:=4���<��b̖�;zRl�����ص7z��8 ���Qr0~���ɻ�/�Ǩc1�9j&[�.�v�� �����gb�h_����"��B��"זXA=��?ա��Ri_ӽ�z(�%��ħ;��W�O0"���v�������ߏt�vz���C���"��5��1��k<�J����4;_��W+֖+�^č	u���raY����ئ���Bb���،����R�,��y2��tzc�Pl����RГ^��8z�WX��x����wD@u}��hX�G�<�X��V�
�f��w������s+o���A߯���.��m�NM���39z?pp��r��p-��"��q�=�TMMk����Ǜ}�����h�W����U�X��}m�vFo� �3�Q���ĵM�m���]�.A_F�e�Ow]P��U��}��E����j���k<]G֥z����Y�l��n��$ʬ�<m�F�'�է��L��jZ=O�ݣ3��Iᾠ�?SL��*-G|M����R��� �Z)]����f�R>�'V6�����ౣ)���Ɨ2��5�	���^���M�VD]��O0/���V�蚰v8.����s����U��,����R����-9��i���R�Bu+�����(�}�V�(�G�������z��b1�N<]-��hP���wO����_�ag��[��b$W���)`��0�v�ƈwY����D���6?��z�������.Jg]������>��ş��"�����v��k��-�o�=X=ݺԑH�� 7XqL~��}�E�/��ٚ�Ei������ar���<kS��匵D�uͽ�׍��E�8���a�b��e��+dT$\5U8�9�h�󺣐`ي�J0B,�����>i���7.:1�Y�rG˅u3�R/L��d`چ��1F+�BZE*%�6l�I�������٧���'�=����B�����D��G�~�$����D���F�}~�u<'m���d5��{~_Z�"��6�����\��G�Ǩ�x{�s��Q �2@g��oW�x����F���O�}w��I���X+��K(U�ziz���9"��=��н�Ѡ�;1��f&��3_|v6Qz@堼�� �(���:�<�'��Y��Χ9����%=�|HB�r(K�ݸ߸#���nn�p=ۄn�����W&�Կ�+R�!d��ݜ�sf��(�R� 
�j;�;iN�-� ��oh�\�{;�6�<r�p�4���yA��5{[ךY���Q#���h$��GkK�ۿgyp�؍��n�!��FM�d�P��T;� z3�fO��2��1���󥢄1��{6��KZf>���Y��lR��S>��K?�p.���|o;�����,����~�Z�.�ع�ݹ�2�2(��'��5���x�D�Z?7�fX�	����[��g5���+v�l�'"~p���5�ѡ���;�h���z��e�Z�p&��wI����S-��׫��L�d�A\��B2��ގ@��E��ԧQE��v鿯�����(�[˟����f OX�=4Hk{�wÒ��F�]f〱�6y�9;R:-��#�9�נ��.zm�]�`;�G95%�m\��#,q��8��<��V����Ԝ8~�8N��%�XFё�(��g�~o9>�S�>/W���i�M���/���v�JV�X�U>|]Hvlq=bM���5Y7@�g\º��V؇(Llԛ���F��'+f�zͦK�)73���2ߟ>�7�콝�&XF����� ��b�}��"Ԭ�T :M��v�;�:�#h�_s�_h��S��S���9��Y�Ƽ�B�C��`W�h@��N��X�J0�]o��Tt�pɨW<4L�`�&lm�M*�����ꢰ�sB+�o^̣��9�>����Rq?gTf�$j%?v|W�T���������A�����3�]�ݩWtoP�y���<�Բh����+s2sҘӘ1�{}�2�Jb���)޹��� �E��(�ֱ�⽂�$�HSډ�i�!r}�
t��ЩQю<��;R�yp�>]��4�'�L�������ƻ]��@�1��L0vO�}�R�m�� �2���RR��_=��Oc����H"	���|߈��͌���@W����g�\������
���r��v$h�o�!򍭉��N�7�싁��@�Z�϶f�1獣��{4��6�{�D��Ɋ�㊯���_jx���s�Hj���k&�@��9:�Agxө�2w%g�G'���G�ù��ݭ׿[�4��fM�=ί��e�-�p[���f�ǜ��5>?�Ď�� SK�x����k�,��q�ve;�$ݎ�[�.�Ҥ�Ɣ7��~����`K��E`�������ǇSսLxE��#�4�xh���/��;���}���AzP���J���t�^��AP���*�!�&%�5@��PC�����]�u�]Y�?f��{�^3��u��5���Đ6X���S@�w
�c��r�����i):�)��@6���"�T�i��)���'�蟣�h̆ ���|IE�B���}X�A_i��l`�q��*�-!�D�����M�z����W����Ʀ?mPo]g��kƧ�+u̯}�#GP�9I�g��B���a�#��+i9��Z�(�WY�{e_g�_�����K,���:�k*k! i:F|Go��<��.y}@H�RВ��{�8rLw>?SW$�~������ny�,�I�i~�On�O[��� ���Vu\�TJsR�6dk3�2쿦7]x��+�[6oj�R�'�Z$���yp5��8X�o�P�N������r\I�1�z�tV}��׿����F����:e�.%h��_+4Y���������ce1g��8�8:�9�l�4�ATʌ�w����3R�s���#Ð��=�U�=�n�ǤQf�Zg�n=��:�O��'�x��'�`��W�-6�k�����#���9+2�X�:_m��O�}��	9V���̜.m�Xb}�EɓH�����-�����MQ]ruuէC_�ɢ]rZ?���#�P�4olhlB���xS�7�+cq��dc9q�1\~�����D`\z�x>��r}���e�dT��%v��qv(�I\wi��o��k��;r���F!�;B4a�`�~(f���q?��t=PXɉʀD��h�E���y�]�
���q�n(3�gU���n�������@P��٨�����zz}��b�\�aC�\p!�Y��z�wE�
ԑ������/1ΰ�y��I(,ؼNw�s:�_\
����-tw������Y�<���C&�͡���j-�����bޫ6�%F��=BƤY��n��)��i1�_��MZ&l���\�sN�?WtiM�<���\��ӫ��QL�xt	z����|����_��ɘM��]�f���!��y�jf6쏚����b�����q�{/5x9�/3���ٮ�(-{|�s�a��x�u�ٿ"~�mK�7��p��� ~?z���F\B��ħ_�����p��ig�ܦt?_}mk/�������ec�Q���Q�c����/��i��M褒W2&�͛�����{+
�<�>�ɢ�Mǁ=	J���&����d���.��Kb�K��=ǎ�hDT��&��y`,�g��`��K���W�Pڶ{������y��Ct�����u���}VL{,.r%u���t8�X�k�ܤyTR��/��N]$�x�S��d<v�� ���E�kzo��Q��)��4X�b���:>�pH����y[-��l�M}o �Jz7����l�	�E�}���w���|Bd�u��8�@l��L��X���J���Wӕ��um��8��WL����+�z�:@��a.�U�IH�ˋ|r�?7ր	@V�j���R�B�d;���[���/{��D�v� ;��*�$4wK]�Q�L-k-e�������m.V��5d���֮�s۪�=�Y2�c��to��^�zSD��NFb�ƫ
�����~)��o
��;�]UP ��C6Rw~Q�r>�����^���y�]�\�2���w��@���_��! }5Q&򟌓��;v��n���$џ�	h���˪�����M46%����~wgO2H�V������	w�C��z]�u�Ċ_���%A��j�̽~��>����L�'%{g������4��D����T�A��������;�cE�6;�ʙ�Ѕ�M�������#��
� >��"��м�c������N��S�$	��ÜQ�.)e"�U9��{ }+vݟf��A�>}�dtՔMr��렋U�1;�֮p�>��V��,]&�oOJ��\���u�4��h(��VC�=�@����D��̟b�������l�Awض^��� �Q#�l�gD�1��/Y�����57�Hl��dGgK2aM�����r���:ʝ'���֝��3n/���j(��m06�����!�	 Ѵ}]�zt9������؟x��%�AM̷Si�wδշ�o]�+D�f��.4��1�5YyZ�o/eO���4��(�N�������n���i��ILl!�1��ڏ�?Ňd�B�!!��5�5}Ǆ�M&��6y6��_:X�4���݅і�6ZFk�K������y��m���>m)2��t��A�T�ҥ>̻�ݿ�/���r���0AsqR>q�S�	{��-S|���'�i�P���ۗ���O���Zإ�I��+A�[j�^nu7�|���
D�.�R�lj��)D��v�~8 �)��\��͡��=:�FɆ�n��O���N�J��s�J����G�T��u.2ƨ�>���io���#��Q:��y��G7�l�|0�$�(	�%6XP��(�0��-�D-�j�C��7�7c��R���hO��ges}���+�N�ge�V��LJ�p�wC�RV��h/h���nBq,�'����)���h������1s�f:S�Ua}��h��wt�,�E[__���83�YQ�yR�Al���ȝ��T1$i�4��$|I�v���Nc�����s2	o��_�O
��z�,J�ԏۂmu\%���y����ugG�߃���܍�Z|hX�^�r�;PZ���D2��<��8F�� C�G�P��u�����Lе�r�#;8�L10k�cqg!�Mq V)��
�CߧiY5ׂ۱��~�@Cr2�nr���(�.��˥�U��j�.�)�+x&:�ʱ�«����nt���N�}���w�t�F	K!x���R�2D�y ��qwI�^����ۡv�N8x�3��fm��{�x�,?\В,��ۃƈ9
��ABj��O&d��4ϵQ��%>&w�]ν��4ܧ�p��f����%8���R���dڅ0�q{��r49�[^xϘ,'���SD�>Q��b�G�ܕh�Xr�|���m\�y��~�u0���pv�c6��!���s#��@�,Bʇ�C>kcgY7x����U���x�����9������Y�>��Le��9:EwS)�(�����cq�vʔ�7~n�x�����¡����l�v6�${�o:=�g�h����n���%UK}s�j??=���)����R�=��h��+C��5z x<��F� �o�L�@7Q�菂�.��ʐ�~|R��Đ;}��聀]��	�[��<	J
oIu���<��duV��q�y�켍�/�U�Rڞ$Gu7%���,��� ��w���7nE��B��$sR�WU\mq	������i�*�lӴ�_���:�GO�-:ݢ9'3�n�,�o��k�܈_�������p�r+�r�����3��5!�:iX�煚Plb�n���]q趾���c
�̴�P�8G����d}�i"¼�?E��J0�[~�f��˖w��+_�T���=��Ncf赆�'�|Zf������b%��3�f��Q����H�Ω�?��IoИ�ι�^WkB���*�r��#��Sj�F��G�oy���<��d|it�P^YO��#��EqmS�h�`&�~R;��L�`��*,�s�3��]S�˻sA�ۻ���*�<����bH׌��4n�x�B"��	_���Y[�ڃZ�	����	薗�+�&R����s�R�7��<QE�,�@�͖߫jp�W���*>M�"�0S�mT�H��E�	�7�[$������7��C�;::B7�ر���ۉm`e�!(��!r���韓AO�[hV&��^5��D�{����+��~
\��	>7��aƾ��z���Q��0�b�u�\�3��}�䊂�f���s�F��H(�O �_�S���E�����`ل��nه�h�#`��tw�*0t��Nނ�?�["�ʏ�E*���-�1|�%�%�WkM<�t�_�
��#��"�z�&n�mˑKt:�Q�ak*\�f$(I;ob2ME��Y�H�!���8{K+Hcu��IE� ��"p�ĶE"�}m�綺I��Pف�����`�H&����S5��C����A�#C�~��z�:w7'D� �U�{�LK�Jճ�G�0 �s�b����hE�Jm�.���&N}��V����]�]�.�J��7 ��� ���I�q�Fb�+{���"�_��H�wyw���H����3��mΟ2�����������`X�x+�wu�Z�2����JČ4
X�G��l�;fW�:�쬪ؖ"����%���]��;�\�!��N(G�#*�̞l�N������`H ��\��\��V�ނ��  /���ߟ�33�H���ˎ��3���n�*��)�y[N����6����H�8]��
���]��Xe�d^H0MA���ײYTD��Z@s
O�j�ԗ���Oba��-(��4.�a�ǝ��"�/���d7�4���p;��v<���Յ�Ђ�����i�ѯ]v�RK��4�0�,{;�V��p���j+�}K	1S��@^T-�K��+&��ϟ����1n���
ug�财�Q%,�Z"R��ʢ��#�s��s��1`E�}ّ��$n� B"ܐ��ܗ�������Z/X�����-��L��i�+�ß�-�Ou��]pJ㒆��l'dqh�;��\�u"��>�pf���h�x@G��=a�ۋ����?��#X�]�,vw�5�Ϝ�Yg�F��b��w1zo'��$����刁*�bOoנ�?K�7�m�ǿ����u�㿠!����Z�����Hk���rr� #"łwx�ꔡ��嶳!����i�/�.�%�h���mϰ��A2,L�͉���֛s�u�i�l��U��t���j(�{�=n2ǘHD����?�ٯk������:(�������m[C����D�bЩ2[|xbw��RL�+
YV���0��5��\*�����֗�h�#8�^�c�� 7���@��ד��9\̋]ݐ%�fz+t��uX��d�$ǒ=K�=W�,�L�qm�Rgv�\4�J�h5Ol2��K���ỌI��tG%d�}���Y0W��;׿z�m��D8����TܠF��mBb�ù_�̩�t��g�B���i5-I�y�����#�в���J�D	�'�/��^@��N4?�P������qc�������@%������Gq�s+�E����CD&���C�W��( ��۴����!��hw�!D���'0
K_���r6
���獉�-��s�A�������E�7>}��K���?"=Fk���}��A��_���8m ��'�=�A�T����Z#�};�F0gj�v_�/'�T_�(;I`�q���� yp> ʯI!X{��l�5���gT��i����'H�I~�E� 0p���z�f'ߜ^^k�c�'�e������K��$����G��}����N��C�y������l���H���'6�)?�.@y�3�������o��_�$���M������$f�[� �=��lP���b��y(�mKĘ�d���5,i�yV�d՟YXI,��c�vw[G�M�����wwW�هy�r�&��	�a�z�����z�[�t���7��$��B,̱x���d?:+m;���R�y6\��,çPL�}�Q��Oƶ�b^Y8b�E[yA�{�0�?Aܘy2�Q�s��wh��xG�fp!���J��v?�H5� ��t��O8����Y/�EZ�@��v%�S~4w��@�E��{������Ϊ�[��>�hf!���za�q�������k�-$�I!0RZ~ǿ?���R���8�1b��F���R�k����:?�l�wOi�%(�(�>Lq�n��}���'U�aF�8�B�D�WAcY��Ϧ�]/���7�����n�Q.9�N�RҼ�L�p��d���\'���Z��q2T�n�����p��% ��K�{�"�|*f{D��l��'W��[����(@@�����d��o����r@]Ti��t{��/�����A���Y��d���ޕ�<��?�0�/_��7M<"W�oC��x���X�ٞ��j|B�4[�����H�G�)�0�4��j�Ϻ�;��S�&��T	0�\O�:�A���0n�B�'�`7�[��Ǽ������J(�&�E��2x�,X��������}� ���XˎoGLG[���-D�yk�$DL&��B�=�K�r�λ�+_Z|�tF��o������\�{��C$n�*�b!��>�������O��.QwˮWּ���ce�AsӸ�#C"M�P����(���dUGAx�D�ֵM�?t�h&p5ovpð�.�Տ�/�����~�ߪóV��b�m�I��x������ն�xd�n^�VD���R�K�*��*P���N��
O�2�`���˫h�ι�������gtsfBs!�
�;�%���uQ�TD'������� �u^YQ�F�t@g�ՏD�۝�r"OA����5������{NV���ciI�g�4�y^h�ԏljGZ����D��i�5��c��ҙ�;pM��h>�>~��L���ɥ�|�2A,�����oR�qPC���[����md�pk��m�LBl�fO4�4��W\�S%{%*� Ɍz�Lbtm�̾n���փS�y��R�^/��lI�Gα[�iٕ���)��Y�7 ����[��6<{��\[�~�ǌ�*X��Y���g�q� ���ީ����XYj�f�����Yl���,p=(�*�'����-ӕ�g��ǝ<�3��8 �� X���A��m[�g�p������De�6>w��r��	�:ۤD�
��� �|xc�.*���VZ���bwH�r9��h`�~�V�O�5�Z��E�}Գh(���Ø�v�/,KX��h{/�d~���(?���H���K�Q��{{>�,e�B'�P2�֓}�4�`�����J��;ы䃣�+��D{�лq6݌ר�T�����Ky�G��]�q�^�d�3�H"�Kw�㡧!���gj��7�k����BWɉv�]]�����_��B�m����g�n��}$���Y��tmʪF���Wʪ	�|�TM�������q�OŬ�݃S���v2/'HP��wX������r�N�ӌ��x�0z��r^��������̹&����.�ǌq�<�[�m�3�C1(k��-�7h4>6�=w��J�5g�:�˰7�^X����ۿj�%�8���I�<D��v���6^�f���Y#��R�:��T��,:,�L3�!�Z�N<��O��v��k��[C�C*�ҧ�'O�D���a3"�����w��;������:�+�w^�Ӣ����� ���
��J�D��_�S����Fh�����׷�e0J�7;��*Jl��~4��T���ՈX1�^,����A��&�۵;t[�3m�)�XG�+������-��z)�so ��J��z/�E�yN)�������V��k�L��!���ss������ȿp޶����;d2��!�P+���Үi����O���s�_⯵Ǎ��7�h,�h���b�c��YT�Γ�z=�z�����-E`�UU�H�xʟ��.@��&Agk����8��}�4�;>�.����Y�q���&��r�c����~�h�$�:�u�v;����d�f8��9>�v;�+�� '��u�6B(���˨1�uf�,�=0�`��_�1�V�fk/��;�}Ba:w�R�X��|�1k��P�[ͺ��[~1U��*�CMeT|��ok�����E9��I}��ܽ��ԡ�쁖ԁ��4N|a\�$��^�%*�;�e�����d�]��21s#��.��---Վ������T#~��Z����ܳ��gf�m�ɻ�?�Vb����܈��cUhu�}��8��[�+�tk����p�u�=V��[��Ϸ�_&I��HKeQ� �f�ڈ���`8���Wh��N�hr̖,���?w0����ZK���n�@�T�Z>n� a� =]�>�l{�hI�KXM��s��c��*}��;%C��*:Ni����)�]��1���y���~��ᡉmW�WJ��3Cc�X��
!��#8�9�}=�!���l���f�����[x�0x��B��-7��-O��a̓Z"��a?q�H�aou���;՟d�h]1�J���]��;�hs��X�?J�C���`ۥ'o	��Ȁ��=�@�ۛ�u�1�CAKA3����L�A�ky#[�`p�-����a2��r��q$|%TCPk{�cjͨ�1d��0O0�>"[*�ϡt��0��!O�=�%is���I[e.K�#GK�d���)"�*�F�S:j韟�4��DoAM��������$Ԥ���x�s~;�IF ���\E�ٓ렩bA<��f=�$7�m��F��C�&p�CKv�c�ТR��L?p\iզ򴰚��πw�37 XC�c��Q���n�S��e��H�QF�/�����[=���V��H�*��B�h�laW�'��ut�P���l)�4ƾb&Du�E���v��p���1��+�K���HtQ�\j4�\0����Y̼����e2s43��EH��6"����_������F�p��f�Y��e�{=�$R�hme"A�>�tXN�AuA���ow�n��LK�ɇ�o��ѠNwu�-�=���$d(�ֵ�u����}�~��j�A�Ƨo�9�Zmz��c�	��o&��.��� �}�UE���_9^��=�����c����M�h~��9���4}_��_�Y��8�;!M�^�0�2�e+���(e��q�8=�f�E;{��{j�s�[ieyB��E�N�:�o+M(hq�C�o���_O�[����h�_F�c�7�u��G7����d����&?�ƛ�ӅfxF�m7]iX�!�|�>s�=�]c�Y6�h��gg�|ێ���?����q�1-�!�+V,������Tk���[�l7�}���U�#v�̫���fM�������w�G�F�͈$�p/\ҰX��x P�uVJ8�m偔�Sn�^��p=��k��z�iu_�THe��W[~h0� I/�/SJ�I�%[~�Vn ��޶�k
yY�u�����Pv؟�|�<Wr(?�HElDg�A�5��RR�W"&C�b]��7Q9�e�>Q8��)��dz_���K[��S�q���pF����n��΄'}g�r o񜁑y6�CEx�����0A�ɡ��j�<��Pc��ڳ��r4��o�Sf�!EGT��B�bf6\���~���O�$��RѻE��o�~
œ��mq�M,�9 vO�1�/�O@�Ot����Ѻ���.��H�� ���Sw�(�u �J2*��c�/�WNL�����R� ^��;�fb�m���n_�R�#>l����1g�8Ś f�������*�j��IkV?Á�~R�s���	>W�A+��Y@����Y�~�7��x�g�T�Qa6t(qH�ܕ{�1_bw_G�����F(U~��7]�OҬ
u��)m9*:`��4Y�;Ul��Q9Z,������Z�j���r�wX�9k�]b�p�+&�6��+$�-�F���	��Ε�ܬ�s��A�R�W�xp���B��Y[Ֆ��#}b�ˣ��v��!ҲWlh�P���E��ͺl��l#A��Du���8�Y},���V��g�h�J>��c�qah��k� '������0pʊ�e*D�3*�~� ��g�m�Ko�z�s���eh��+J5Y�)��Œ�.�?0��wٞ�P^"�D�8��;�[���JP��}�Y�SH��E���DVv�H���#G�e'�x)��8/�).���u�J�����J?k�V��f���f�P�=���rW�;Ͼ'Y@�c��(�QXe�&�5O�Ь�I�İ�����x�У����μ�$D���'�ꣶ�+m�"�^?����ǈ�Y��7�dKxB�w5iijv'�^ԭJ�Cx���6~�TLE7:lS�HB��N��z��}��¸�����!l�����=�+VTP��7Qc������
%C��̸0%�*������&{'�����SV恙�C��%�&#M��?��{�DF���Nc���
?�3��НE�{�nT�]om�Y1�J�yu�ɟ��TW� V||3�����?�^[�Fm�Y�ϱ���jj���3�S���0����٦�����#��躟y��?A���4�"��@���C�@�%��{}�%�z���e2��6�ZK��#�
0��-��]��M�Юx�l�(�j�Nn �JX;�C�[�l���y��Hq]��z��Q�}��yVXI�]�ߣ��"7d��ώW���z���F{���4�����[G��V̽j-lN��߱_xl����6CV�`-���w�f.�*�2�7��UYX��|�E��c�}��	@#hpË|��]��X���Fx�YSg�,6�:�s7�v�;�W�IlH_�͜�� ��>�$È.�uĠ{֌٦�%������=�G�4Y���u\�#��%���ۑ83�w�dLV�]?�a4%k�zy�\y�5�R<�.�ǅ@%��7�����������%Q���M�T�¸���XMEW�� �p
��k\y���������>j��t�B��Ί6����m���rS�/��ˆ��_�3g�9DYLM�_ǽ}�sh$&F1P��񒽎�������zP��U����@e����0R��|ѩ:=D�۲X�bA)0���2�~a��O�	��'� ߮Q?_s"h�m�&9�)�!�)��z���ڌS�vZŻ�p!���"yM�j�ވ��O�_��uٜt��<~h���F��\QF�V��Q_�^T@���R?O>\���x��jJ�|A!��n�ex'�>=0,�Z�s�Y.�V:�OZT��|ܳw���jF�7��a�[Me[��͛�0��;�ggl�S�J�B.��_a�}G8B$�s��
c2>�}�O9�
~g@^��B��6��A�i��3�h]��P�v�J��k����6�Qn��(g��Apx"��vJ�� �h�C�2/e$��!C����G���-�x�P�K�^�=�iH�2s�`�c�vHY�<]�O�q��<Q�&t}���Hd�ԡ[1�ӟ:��ڽ��h��(T�nn���m��ϳ��kS.�rw�P���IE��/G~@��%��j��~<-�,c�l��+Q-`��;�ɰ��y�]�&(ި�2[��㝻��E�2��%�8r��~�)�ˉ��7$��|��_j/�¿��<H��2rv�@�b)5��'�[�M	L��������h���ҷ
���U�5Ҽ�,��B�J��A~XCxD����`�I�o֕�04��=������3Y�U�{�����P�i��B����N�����gQ%�W8��)������C{n�A��k�l��z�k�f�g[��� �c�������R����;wՈE�^�SuU�m����>�p�^5�s0|���>����n�bw��5p?pmU�*�E�7� Ww&̡j{�{�*���(�W�R�`.�^ɟ�"
Յ,���
:<M���y3 �:�S��y���7q��Ϛ>��2��W;>��r_�x�2{����V�A��.5��\��B@5��Z������q�C �:��8���`)
C�`����>	�*�5&M�0�؞(N������L�;&�� 9Z�&��Ҫ�'�<�mc�J�S3�oZ��<d$ϙ��?�%L���p��v��U	��{Q|�R��t1g�W��H�$ƨ���>0Zk�c�񮅙����3��t�]�� ��6|E��re�s��Z����Zw� h��`I����~���T<?�luRc��
���1���S��v�_�0y������V�,��??���26; �C�]d����H7T�%MZ��+#Ō��/|��6r��c�P0��0�u-u���<#J+�}-rG7�`P��|�U���t�A>��~���b�m��F���nl����=�+�0���������$֡-�N:`�#�P���)g:s�V_؉�H�������A��d����"shO�y�����D,���P�CY�Ti�.����-�Es>.C�"��'}%uއ�D���cP`�T\8�٥����l_�'`�_j?������P���J�~	�q�*���.��N��b���e�+�Og���@�2w�� :V�l��iq���7��m�W��cm߅t��?��ޕ�{�(WJ��_�cP�!P��yyn�8�H��W���!�o �������&xg�\TI��.���Z��=M;+��'���V��y��H�KR5��ȉY�b'Y�0ϹN��Y\u�cK9G���*Z�'_�#ql��@��]SV�����<ä�c>L�V$K��7�W��}+t�
�B�0�#�[����*x�{z_��΁�\����63�4�W12����`�G�A�����9h���x���8@5������/�	�'��taԓܘU���뱙���~͏�$���>zh~
��x� (��=]�9���x�=��S���\�o�N�{�S�͚���9Q�_�	���C�bM�L�nYLy)��]���ƫ�8�:�Hf��p��D��r�q�M}���f��D*������7�-���/R��o����@jwGT$�\���2�,��^��~�J���ڑ�p_Aj�"�"o�pL���b���j��'ʡ$%��[i@����;����?��x�z�,� ���o �f�c���Б���*��P��\�h��uN�Z�X�Ѷ6*i[���$�<�
^��򷇙���Sacyгyײ6j<զ�	$B/[� �W!Z��w@�`�G!����3��Wu��tO�*�VٛRe�h�!�@��۵�s,\�2��|u9=���.�	�a�X��,�fx̞='���n���������PU��Ύ��I=m�7�A�1���}��<5���}���I����}�|Y�H'Z�âE�2�=;k��N�2I�mL~.>�\��߂�撂����6��	�t��4��/`�Az��/�_8M�@j����ɑ�'A��^�����ܰa�?=��-��z9
m�ʖ�|p.��>��v R���q�o��Gq�^L��*�Y����<�%5���8��(��a���D�["z���u�3ݵ$��0�0�jS�;�4�4mn��b�����a��Dw�tͤ��b-~�t����>��`��%�cߠ�Vy-<�֋Q���$0�Խ�s��s�a�Y+�tV�,Af?��o �ձ:4ӯ��z7�'k���-�`m������Y��)����x��a3,(�ܖn9<�Py�fK ���\�}a#Q�>_FT0fCdyt��6�L����1 ⴗI�����@�J�q������rpk\w[����p���K��O^q�Ꜯ�,R'��::u��w$�֖?�BV�:э-o�)Č=� k�,ִ�}~)Q�
G�֛n v�0N����Bo��������TF�����L?\op�+:	[���ӟg��8\7<#�\H��b�(���6*e�SaV��NTbr�n=*�β�]���"μ�j6
o937�Dc�vPW%�J�UFrM��[�4�l5����QW���""���(3E�ZM��&�Bm��X�b~�����-�����(K�K�K�7<O�/����\�K��/1�H[N��w�FKQ�l���gMz;��P<����K��!�R-�/�}���GY��	�W;vFd��C�r��!��b��`Tuۮ_�#l<! �ͬ�j2�C��A��u�Z�/��?No9▘���~���$����\����{o NPĕ�Ok�@�+_��~�q]o䲷�:q+a�/�H�1�ѷ=�A��VG2�q��5����!m����t~��M]��«Vyc�a�p�Y/9Z�tz��gA)�s��R�HN���.�����SkY�ҿ��[�Y)�$/󯒆݇��4 �dr���XS���S�{�?�E�C"�����Gg6�7X�ǳ��	�8��L��p�4/R#mU�M2K����������i��U�|�4�؎N6T�e�gq�����Z~��x$49�9>����A3��rs���ZX#`שl��ǿ1��g&	�QTܮ�'��)=5��g��Mf�;c�KщW��a_>�ǹ�g��\��j֝V��q����m�?q&����1{���W��/r51J�@��hec�ej)"
?�-�^�rK��	��7��r�)�-�ڈ�REۭA��s﭅��H�)����O�L�����7�����ߑQmv�,T�u>�,���D�u\�44ё]�x���� m��0G�ܖ����+�����!Aɱ�/ax���z��]2�lT��Z,�&���L�yڽbF��Q�b{��l��qs�G>��<3}�OM5�/�FBA�E�Q�t}Qoz�G= �9?_��K�46 ��C���ߤ�W�e/m��or�9[��\�-5�F�@f��=���P�.d�i�*/ӢH�����5|�o3�ka�Ty�)3$|�gJ<Y�ٝ��X�!p����ˮ��b3? �Mb��&0,���묕��e�G�- �F����He�������Aq�Cߠ��V=��i�����4���i��l��_�De�%����;Us~�V9� Δ֬���]MW)r����l24��`hŮ���D����_���(����(���'���J�����)."u�����Sk&���s4��ϝ�d���0YC�O���F�f��3$��tf�o`]��P���?�I��b�j��C��_����8�����0شx5��X��y� ���Z���	��_���'o*�~�������� �F���ZN�|^ �]/ہϕ��r��O쪊R?�+�}�NU�a����y����%�ؤ ���u���U�\��� 	�Ļ�����C�KV��
�m{Sͩ-�f��P �{S�nv�,Ksɤ���W�ɛv%C�r]� �s���S*����*Y͌����KHøh)��K�Q؄T-�?	�zkQ�	4_+1b�{������!GfOF2Бh ���nq�����[���&_��C?n7��(�ٹ��ŷ��u�� r��W���H��B�m�3w�n;!���B�����[Eh��;�����O_`囯z���r��Q���7�-]t��EĿbx��W�C��S�Z�S�����|˱`6k޳*�B������u�)�oY)��Ȟ�3Cn��[;d���X��� �{�2�4�v����q?����J~PS.�`ɜ*a��Z��e��(( G���δ������[�C^���@�F�wx&��ǜ����p��*s_��<O��҇�6]�g�N��Nk�l��	�v��L�xs+	��&��Э�_�	Ȓ�E�-)�Z�f{|�����]��4����⸹[9�?�s+e��~�!��Fл�Ҕa*a�c8���rGu_���c��� �_�Igi8dy��%���R��r�ßeR_,��sT�gZY�}�WhNe7����*_Z�,6��%
���؈�Nm�}+���+��k�x(L� x#'�[����q���2�`K����ȣ��A���5�������x݄�}��<c1�u/W��r
��)�F��."W4�:K��`�+��XZL+�@�ΐ�|Z��ۈv|��(�ڦ�&}e��JL9������Y%��ͳ$�Q%犻�%�Y��ncLH� s�0�Y�����h���(a��8�������M�X���-*�na��,�ي����2�S�6��cW��;�� xۊ�9?š���TE'��������kWr[����A�7F;�/B�F��͈G/��<ƛI�w�Rb�dx�G8���W��&����Z	�c�lK'����x��᪨�o�Z�yR[�Y�Ȅ%�M�2��i�W8�)O�����XpRMUWZf�C��cQ9��j��ʶ���h6)D�v��Q=2���e6D9P��KD��	�߼�a�<�c��s2�9��'�7UYI׳l�J���+��r	1�K�ϷFĺ��[�Ƃ�7�!����ͻ�[��L��1
jL���M�ɼe����ܰ��@CB�����Q��F�Jq� �D��D����j;=��
C�P�->���R�H(,w�M��^���΄��[Fw�f���Ѕ��cB'd&�*��~�"�=1�Ҟ��:� {FmS��Y��@����}����f��2�E]\��y��֪9D��R����Mf7)����g�",B��@C����x�~.�>H2�?
�i�-f}���~PK��s�B��oN5e��˼��Ryt��E��O��%��M# �Mwh�*�p�p�1�*�{��z}a�^�W���
�e�:���"��u���~�=�� a���`�M>�x�h�oz�ɮ�_�ˮ�ug$��������=����w� (*MA��
*��^�    ��H��B�i�����"5���$�H�����]�}�����u��'+�dϙgf?3�K���;�T� �z�0�p}���� Q��-]��v�l���,B7�i[<JYL���AnW6
��U(-dx��.-Jz�:&4
P�t��ζ��@�r��G8���kwʠ�E�p�_uݲ�l�Ϗ�h�k�=�|"�P��G�u�[�cg���p���4+�ɗk�4��j�J�C���[s绊x����d�Ll�t���`]P{i�[���;�R��������M�
_�
��D�LI��c�ב���
�ĝ����`>;��yU�	��.+Ǟ�%]5��E���?5!�QU.��R9��Iz�n��E6�iɲ����]J ��2ᠳ��N8Zl���ªEL����j�M�ϓW�&���a��K�3n�n��u��-�ى��bw�#������큗��{F2���J�W�]�_�U�)�N�	.SJL��f����M�Y��H� ,���V�L��p��M�
��DUi>�O'0�^s���f��b�вޕ翀���?7g�i������D�6�ݙU' ��	�����+�Q����'��dɩ��1J&�f�];o>��,Jv��Ҁ��"����ꇫ�|�eʬjK�������oXx.-%�&@�U��d�J�������a�wMS��W�ôP,^������<�L;�X��;	�א{�2!�Y����K]�i������=xMQLO-��t�$l�� �=��؎�^C܏Ckv��m�Y���Ĝ��T�pN9�D`��SSZ�-��#��� E�t�#�
�w'`&�j-H����Һ����P(�����F�-p��]�'��u�3�`��2��u��ޱ�>�:�V5�������D���G��	Ƚ����c������J{�JnH4�v��aG�3S��E 3X��� �]ҡz)F3���C��]x�T�qQ�F�t+q�$�V=�Pm��٬���*�m�_#�7G\����ܩ0|� G��MW�^�ۂSu
�tH�M�f�v�2fVbX�/�}�{�s��7���u�W^R���u�v������b�߷�Z����}߲3tY�P�9��9;�����~c��E����zH�d�V#�Lxڷ�ߵK������W��s��Q�`3;�]W7�=|�s�	q#?�n1|���f�L�$M���5>씖��%k��׌�M�.���;��H۲D��x�H�
�Q�nr?:��z��q���{�Hɻڤ�h�
��w�E���5�QkG���V�R���l���2[���?�4j�)tk4��p�.�@�\�8%�}��S�C�:C?�������رE�x�K�e�\�T�)�%K��������3��_X�YT��v�NHW�Z��[=W���J�L�C?IO�j{�4�[�(24_FW�Z�[�uӜ�Cj�X���� ��.��?�w<X�Sv�������&QFP��SBI�	�5���RM"�-�jb�'(�i���'l[�\*��c1���g�K��ݶ�e�cR^僫�Sӥ��%���
g����o��-	{XKH��՚����K��uXvkNR5�I���-�f5ܵjI~Ow��	%Տ����!K^�l�M�|i�0�,�9�ـ��*��[U��)�Ix��,fff�:N��}�t�%�V޶y�D�@�$�N�#*,M�x��m�a5�S��nr2��zO���!����ؒ�����K$3E`s�<��Q�������~~o̥/>��ޱ_RO%6tg%������096
��WNfV�o��D��O
�|�s�"�[�9���rb�
��ro���BC�%�ˈ���̆':�r�Q:a��hS|�c�n���4~/l����Y��e�;_�f*���g�c��i����p�=K��@~p�θ���-2����iu�Y0ea�+��#�
�ꉇ��/�cn�<��g@6�Okλ ̇��'Ez:ϙ�D�b�4[5�8�/���R��ʮd����Y��=�_�����#��f���O�=6-��\���JU�e��YS�����W��h��yc�0oE�:1��R}A_���]3]&a���1�Ί"��:IP!%$p$�FT��j�S"������t�]�ݧzH��䪾�F�'}N#r{��ʢ��i�>_|��'���!�ڹ�I~}�=��B����r.C3g+�^��腳ը#+*5��Z�k���ȉ|�h���V_��e<��J�{,�"d���r�gRDU��	_ \�e�1�C��l0����C����7�L��v��\�^m�2?szd\	o���/�(�	��W��3d_�S�{�7ܷ!�N�ыq���v�M�Y{yF_���3���ER�W�M��f}v����S3h�Eu����i&�V)�P�3t�����鑂�����|���>�01b'R��o��z��R
<��$�h~���P1�-���Ɂ��-�î)�aqE���a��s�����/�*ox�{/b�\}�!8�y0�<V����
-�1��m�XK�Ęr�P&�M���ɩ�G�*;Ro�Y-	N��){��Ǿ�^+H�{\9��k%n��?�ϞO+��LN��O*qj�,�Š�9��x������A*�B�eX����*��_ �=P�i�$6�띰�[A��g�{��z����+%. Q|n"�{��s�{��	��G�2rGt�]�u�/�U�$�Ⱥ4�D�"�&Ӓ���r.�kS�i
,��9�B��PL����\��:��	�Q��/��v"s�ߑ�^ʜ4��8�@�+,S��yW$b� �w���w\��~0_�bܝX7�ӛ�rnW?�s���@�"�0?Z�c#��=�Cr����Ŋ� ��Ot���˃��Bx�2�4�J.ƴ��[�x-b��it]]�\������t��8ϔ�٨��ޏQ��S�7*������נ��w��n�Q�R����5�Ϫ�+��6j��y�G�K�E���Vm�_�Y}*"��I��e�bk������/ ��8���j�V�	e�9��Kˀ!�]pof��8x�S�H����w�A�K:6�|���B0����lTP�	�/��Vڏ`_ɉ�c䞄���iX ��m�,g~�>�K7�ӌ�K�s�Ki�j?+�:��qؕ!O����Rv��kz~�� �p���K`�������|<nB~�C��FmkѪ���/Ŗ��e��LT,�5��XsQ�0!+�x������+���5p�P`l�4�����X�h��D�͝�83�+ec�G"r~�X�Gb�|�.X�� C��}wUR��H����-乻\�I���e9��يoi�����m	>󦸚�<��o t"7\.��*VLv�e���>�~E���O��Wç�������q�s-;�?�x���b�M�]�@��-����"`��1"�%v��T���˵Q.0X�nx,Ry��?�I�fx-���SܦfՖ��/�M�s���k;��L�[$����	�Q.�ϫΞB�`��\�|�ȪXW��$�!�N��In�����Aߟ@*S+�G��a��	�ݬ�5֙�T�Y�+��D�Am�'P\�!�b���qb'����{��\�(�S==����L9�o*�L�����I�oB�b��rl昙e�=����XR��ET��u*(�����Z"��A�:��oǩ��M{lC��I��S��y7A�&n"�*�r���WVYH�[4Jx_ n���	�ڒ���e[��Ժ���k�-�
�Ч�4���`�kƣ�{Ae�����l���n�K����5f��䇥Q1D���`��@�Dl��1�q���y�T �|1\�����)��o�qjZQ�´G6�;�[��sŮ�6�IIdEp�2��]���O�����~b��nv_	M�r�ò��`N�Oo�.������[7O����k�3��������"U��P�l��C�༷��Y���w��yWn�ѓ&귫����7|�ɬg��e�6����=��"8�N�NS>�����`x�	[Q�8�q���L��[Z3H����y���t!��w�k���K��_[hP�3��Ƴm[�&��y}^�h-GQqC����\ZM���+�Y�ۢ�-�s�5 v��/�krs��Kԯ��a��;��_} ���>���5��
�uyh��%�а�e �� ��$�8�~��AKZV��W��%�a�Z?\O��+��+CviJE�+��3�5\��ZTk�������uW/_�Pѝ�o�'͂�+6u���L�b�i/�����
��#.�\�o�n(:y���8R;���G�kҖ�n}k�����xiD� 7gŔ���̯x��p�Z�t��N:L )�a����D�D�jg�1K� ��(���S��$:�8��鼺zfѫp���Qvj=C�nL.�J4��Qܲ.xgi!b�H���?���״��Z��:݆�Xt@@�~��}����4f�~ݱ��zυ�<S�����G~J�g���o�D���IWˍ5�#/I����|�P2��=�D�6�otN��J�~�*
P('q8��ᅖf?nv1�[t�}�5bz宺�����j�����[S839��M	H���c�Ӑqv��a+e[v�|AH�
Õh�;:X�U�5�79ߑ1c%�[8H���o3�}	��1�A��yc�f�1�@����:q�q��`�8��N�Mτ���F��-��Mc��z�7|_�AFk�0.4��:�Y����8R�L�Cr�N�S����0[;F�V��c:/��g��_�x'���Ӈ''�������E[�N�R�5���>ĝE�n�^�o��"��e�d�B9Qz$�Wr⡿���3{������m�o�
�Q�����ݙ��O���re��XƞA���2mCN�	�[K����*l:�t㌎J�bEH�N��P����&�od( 9�m�J
��{����>6]�����6*;L=��ܷ���_~ϡ�ZoY��m����9@SMƜ��9�D�Ӓ�k��S��X�C!zK�
�f���������CqE����5�}���U�cT� ��B��c�S�a|C��]��pFf����Dc�\"
?�eN�G<�z���O9jA�*�m`�@�fX����0-���p��I�&�n�m���Ւ�O�7��/Z^B=��Z�fz|�g>���<UZw[-\h�s�ꐕ�[Y���� \�,/���7uG�����������@�Z��y���[5ԇ`���������S��<�7����k� v��$]�����_�Y.���Wn�� ��(��	2M� P�.0�����;��3ttVS'�T�� 9:�H1�f�����\��@����>jrL�<~���L���j�ZF�h��ʖ��Y�����֜���-�$aX�֋�K\���o��Qi_S~#M0�:Y0�\�Ay ��\�,pM�?���Mn[m�yM�Ɉj�eK�,H�k\J�Y8L�w�[�!-��僸*V��z�	���^9��%�f��c�ye;��:��	���9y���m�L��k� ����GnxTMY���5�|X�e3mVݴ����p̈́̽�t�p��j�TX��j�{us�u���je���y�������)oe�L��U�ʯ��6��ssG����������
g���JQ�o��B��~���%�����X�(��9΀�'��lr2+E�g�f�*�<]�8��� ���F���ߦk�-��|yt���i�۩����a��樏;�s��y�Qf8e�vt�����+��8���4���ɇ����Z����I�Ȇ���g]ԫ�I$��l�c�af!픴-Y�&l�֏8�O_�M��V��'��Z�G�ٺU��o�����I�zR���]��}��Q���'uog��(#�*��;聈�ۣ���o�?] �|`���֍`N�m��ǳ��5/�|�N��!��f��l�N�=i�N~C'9Ԃ��QR�儇���{�ȧv��-e������7`6yƞ}z����<`�D8������U״��VG���&[���qv�
���o��ocJk�T�>���~�$�.lk8y}�|&p�˖�ۋmq��Ӭ�����hXp�IJ�V�(-���Q*�w��㘧Fl��ޯ:I������[iCP�S��6�CC��qB.�.3g߂�6���<ﮬ�)�B����Sk��o���. ���#�a!q'�{��g/��ҽ��ucYy�[�1-e���"����mA5�͹��i_�ɫ�
�C�����ѯ6�W׫܁ǎ�{]��vĹbS*xO�(��yŎ��f^fBl �nç�U$G���,Ҩ��}ӟ{�NPʧ�ΐ��ۛ��aX�`��� 8�<h¬�Qy1���Yb�s�� UL��Ba�ƣ�@���UP�}/b5T�F�����߂��<(� �U'���!U[M�J�#R�2o��w}4N!��~\~7�����j7��[j�5���1��Y���!��s9�K�ǻ{�j�˻L�%es��5�|j_��ݩ����a�=Z����:{��b?�p'��>u,�j��?�|��^���g���轔����=@�T#:C��'�d�e�ͱ����ש�0�?:���sf!��,ue�ө���W"s��0�[��+G�$�E�٘{����' �'�{[gf����r�?��h�d��V��aA�z�hv79W{��|P5�h�)�<
��3R9<m*�R�s^fj�����o�y*�{EX.u��l�,P���A7QT���oU����%�q���h�d��c�����H��1���*�|Ç�ӆI�^�騼6V�d�%���aYk��Z���m��J�����?�nO�`$=�Q*�½�Uv{��ڇ���5M�Y4����t��>�֧|���7dj�5,^����pDg�s~G ������ �oi���cюn�����Nb��u�՛Nr�Z�r.ױ̰A�I�ɣ�Ď�}�w�����W7��{��2��N�nh��:)��"��j�n���m�e�"������� c��%���;�y~�.�k`:g�����c��^j���XL݉�Ds�yu�`?�&�@��\-{5&m��VA�ܵ��7��̚�6��T�Q�űY��7���v_�Ĳc�Q�G�������e��NX}�?������5��3.
����Rw��$�gH����(o}��{�ˬt���u�ɟ��{'� -v�/��0���4	-�]N�/�sW�("jA�r��dc��	ɳ9d�|���Mw�A�ۧ��ֳ1Xa�d,>F5���#�S���԰�(@⶞0E����W�Y�AW�R����'	�1�3��(@Y���Tòst�m}�M|���*gz��c.X��y�qZygСx����z����yxB�B�	X�j^r���`?Z���t����U��ﯺ���]�sv�?��6������g��:��y1�?e^y�ڊ ȅ�s��Y�� -������ךg#�H]�+/9 ��[	>�/ �ߨ-�qt2C��xxM��ү������yG��fM�yF�Ƀ����/�ө??m�2#�j�iF���(�0��j�U��Fy�Wڌλ���'o2�|<�Q�|�~UЋ��t}��庑x5߆�_�̇)�4���%��:����I�h\����Le�˹}*��1d%��|d�ZG?.+�a�����v#��L�5%�x�n{��:
{�f�ϼ��{��S��Z���p��_�Fޝ��ne`r�'5�_�����מ>��)UDԀ?���V@�-�i��(��ޫ���ql��xIj]�m�'��,rCh4�ێ�P��ڎ+o�>�x��aG~�����V�iW�=�����hf/���G��0/���9Aތ�r�V����K&��gO?w��$֢*z��
�	������Ϩ:;��T�w���q�_M�^��[�s��_���0K�6:�Ţ�Z�r��G>�jQ��)�b	u�


�&�܊,�{�3��=�c����s�?�|�6.�&k�V�q���CT����\~c�����f�`{�u#WQ� ��鸅�;��תZ�M��e��yCrY�-���X�I}�pM������LXg�I�)�oc�d��c��h&鲻ݶ�g=�L�}f��v_ �f�l���Xw�ɰ�U���h�iZ��Y0�#?�؍	o�,b�J�E�둇���mN�V��5)h��мG}���Kv�k�ɂ���:VdL��YFZ��/�^|HC��]$�5̀$Ͻy����=I=�f?Ap)'ô�OD�s���c!�{A�*���9=H����w�Ӕri$��Z��^� ��0�,.||�4�#��������2[܇	ngS_H�:���Q��`uT����|p�d�:F��D�n�Hs��I-3��!�~�Z�/k�E+�b��:�lK5�@�P�	\Kv_�
�O����ƅ$�V�e-$	��#tK5?��!��f��S \�=3����0��S��`����F�xɇ�`V�g�U\w��B�n���_a�8��G�A� �q阹}k}Jd�O�|�?&���.z3����Q���$���Ld�q �1�R�j�v�>qЉ�&M�?Wޅޑ���F��tL�1b�86�sfr���+vF�e
Nv�P�B�5sV�\[/� 6y�)V����. 5��jr���_��U�u�#�߾�ӥfXv�|�PmTǨ�)�;)b����8)0�,%��O4��W%�WFI��R���Y Z�b��5y`��� :!>�����tgn�Sw�RglҥoR>�Z\O3O�V�ba'G*oZ=3�ߴ�߼ �{F1)�w~��;��uN��u�R��߅v�g�#S}�9��8?<�W��{��IN�^T��o�����8���~�kw��s�o�����@�CS����q� F�R��s>�����{�Ԇ�ԩT�Cw�Dώ
K�G��/o�9�����
uX�0I��m��!Zsњ�)M�;;~Z+G����c�I�w�-TWf�z�~��uK�JTt���qP��ԃ�<���ُhZ�͜����'E�D�r]. 玛��l��th*��@$�ך�f��~N�]�f��d�c���@a'B�0;���'�ݫ��6��d�֌����� �����غ�w>�BQF�y���oȫ����/�)\�&Wm,�v��J�
,�=R��ez[���!5kզy�������_����v��ҟ����$Yn�� L�����CF���T�-��s��19z���
�Fفd�LW`���eٺ���?���] ���z�����au'��"*�g� �9�l�˝�t�zF���R�.G i��ؓ �@>��F��!ݽu0 ���Wr)��Gz�#��M��|u�LJ$,�Ɇ�%tq�c�P�����-˳a������r�J�v/�lS�L��� $qѭ�_ �
�n;��z�q�o.5N���O�jr�&_ɦ]q�ii�~��q9p�Wh�����z�\B�7��2����1�y����'�|��M��̍�)'ht�nZ��F�ι;,	�0�鑽SA1��+.����:�V�o(�8<ێ�������;�l2P�:���I��^��;��[J$�m��jT�¹���ok�[��|�1�9P���8�nB��r�ʴ'��D�y$s�X�Ѭ��B���4����:�e. _�T������n�գ��L�Z������_h�&�C�C��]ͪ?U�/G�c��x��$��='[ #Ĝ�=�����GژN��%t�uA���] �]?����ڊr�P�4����S�
l*f�3�6A���g���ؗr���!�$��ھ�1Oof['�#(ؗ`��=��X��\1�^L�}�s�sǙ��M5ϕ{�Փ'M�\��yM<�u�W3�>�7���i���+1`����AU� �}�Y��mԤlS�sU��lˍ�`�K�q�/�k%�>2��4!׀�YT_m��l"�kޝ4]� �i/QD���Sr%�yې������:M^^�O}a �I�H�#���Ӟuu;�o矫�s��[�<�>a����WH�ܔ��ֺ p1������T_�Ԧ���qHujJZ���q�����)+&f�<P���S�P��g��OG�T��lB���N��еf�n�kss�g.�g���v�Q��=���,Df]��ZM2���x�0����JD�e��.:�L�_KA����u��Dx�W�^���΅���ڌ�ؠ,e.�ٴ���#m��>Iל,=�!d�7�t��J��[��6W^���(B?����M�`��������j ��5� d&��3�SVK���x������<��Cq�SѬS�+��1j��@���F
Үa�*e�4�Ϯ���/��RE�����_��7�}�f1ɭl�X�1u���O�#AR�f.���ڛ��V����I��@z��6�\�z��I�wc���	�,����e.:ah�x���od��-����$q2�L��-տ�J�!:2uu�ޱI!^}� T�:JeɑP/���fHV�Ѫ��8�~b/)�He4�]�b�4�R��-8�'$��C�(�|1���3I��j���C� ��影s]7��(��\'�i�EN�U������1�vـ���E�-4��1�q]x��6���4W_M �o��#m�i���墢UJt�R��Y�a��$��V��ͱ���lZ��гY��N��Ow϶&ͬgV��i��J�B��!'>Q�fr�������[�u���.�z��ۛ�e ����jU�,օ����T����-6�
�8��,D���Ut���Ȫ���5��Q�z䌐)�;?*�̙���"r�]˦�Z��*-�S�-r�K��;	��<����e?���*�2��Aq,�^x,"'�x��/ӌ��ׄz�j��
%�+� t��Ԍ�#�x�	�����\u�Ê��!���*3(�����5T�\���c���H�S:.;X� D�C�j��X���M�\}��=(EQ൵ޯ�����"P��u�[�K��I�4󎕳0�����[F�J�_�3Ϊg	��x6��i�����?�3��`��4�ǌZ�H��tkiɧ峸֒K2V�ބ��9C,�\m�8w�)���+��d_�����1�}ϙ�(]�2-��W�$�p9��k�T2iB,m`B.�Of*���N�,ua��X�I��>�vR\ݗ?��k�*�;�)��+P:��*ו�f@G�56z��R7q��MO?v�򐪡��hXnN1�Mލ�[����k�%�7��]�W��o����A�5�=��E�>���"���lH�x�?��W�����Bw���{�
W�bH����*S�9��A>�l�n�.ӵ�[k��D�
}�.>���f[|9g�h<���W�O����2������p �80
=X-��qw��h�̪]�ʃ��o�s5s�f^��~��D��q.<����s~���S�ݳ��y_�ԏß�u]�4.���+�r�н��r���ڌ�Z���a�Qң����y:s{T��Yz����֐�r0�6����L���t�y����Pp�?��I��HSA'��QǩCc��_��XS�
Jo��[��k₺�g�1k�)�"�Yv���8p�Ȩ�p&��,f�%3�2?�i���	���� �n�i�搝쟯�5��N�Z�Tn���?3}d��5��]"�`A�e:�Yb��l��U>�{}Ed8#O28@uχ}����ݠժ��[�kL�9
 �Zz�,1RB��e]�q`=� D�ޛ$rb���pKw�kFՅ�$<�3{�����n������#b�Y���M����
��d;w�iy��D����f���7/ m\�y�P^��%:4�-�q˥���y�����xs����r[ilW�rk���b3
�+q��ٴ���C����b��R��ڧf�ӐM��f�ĳ���_K�o
�MO,�d�\�F��̫�C�����k�?�N2���?[X�{o�E���)�� l��aG]��;�L��}��1��7W�YE&�Wg���qYM��N+���np���\ �tt�gT!�j��g1�7�0��?юC��	�sG��1��]6�;G��҇�Q�9�7��/ ��ү�Hll-�@��9pOۊ��T����i�J��߷��Q>�*�k ;wR�G9��(�/h�U�w�~����� �N`�|f�i�@e<me���7����r´,�:N#����,�c�S»R�'.�;� ���$q�B'��ެt�_W���Ơ��W. aɥ����
w��. S�fK��9����$�.w'�J
�z��l�ڹ���	,w�i�.!-Ӂ09T�y��"�u������`��>�R���l�S�H�"�c@���U6�D)l%�1�j��=C��t�{N8o~褉D�+���H���i��vR����4�4&���ŠKo���
7}i1ռ.�/���*f��4\����6��-_LJO�Etj�#,�6����-@8+	c�Z��o"��:8?;Bo��#�jH�uM��jZ�����n�h��e|hG3�+� ���m��<$v��� ���Td��TI��`krz0���J9lND����d����7��u�C=^,ϐ�"J����� @ް�;�u^�q;҄2�~U��	#c��ڑ��1%�VIR������sDd3Z��;E��*ho๋7h�O4�\� ��Lv�k<����{.&�OK+��k�G���g��m��G�)b��o���Rq��Ə7�0Q�f�f�>�?�7���/_��ؚm��c�`�,\o���n�������.?�#���[3?�8O"y�3=d����(�q��bU�),#{f��� �r��	>�ק}�Y|n)9\�PI"ط��`a�L��ɧ��e=���)8�����:8�%�卵09�x�|�6�}y̳��
��k܇�,�N���ٹNl�����=���rM�C�D��l��̑�^����I8��$��w2�*T68�V�n�W�qEbr�rT�n���0*�׼�G�i�ru.  ������䋧��8}�hi�X`��F�	Qi�1M���� Aܝ�3�m���4�G��wڂ���n�0,\B�	��ثziR�p�:�픥9�Z~dCT��?��	7��㖦��㠤&�ڸٿ5������.�nE��r�+��L2���DQz��"f������9� 0tto�bb�wc]�󘲣��J�D�nd�����r��zV�М����L��c�.�>�Uni��P����@���#��ߝ\���2��q���:��TN�_ǔ�p6M��Q|"o�ه�OoHր����6���n���: M{��Լ@:o;�ۏ�+�6�X�}���e�}pڟ�`.~����<�� ��P��������7��%�C��\깟J��s��E\�v��kP칀���W0Z~�f�ި�e6�,���4p��[�>�nbj�?�:�<�_�~H�����u�v_-�U-d�(]��5(g1�B�S�`��\X��嶠׷Lk��m�Q���[��[�G��^�Ϋ#QӠ���[⥁���^Q�%{� ���?(�nFWuCA�n�x˛ؒ���{�MۡY�3��܀�8�b�lwh:TɜP<�@�-����%rD��F�VШ���� n!	��;f�M@"����G��̔|y/k?
���}]������(	�{\ւ���Z�/I�Ǫ���=S��iv��, _�s ��94��.>��7*hz�E�a)�6��VC�}Gr�]�xqo&�6߷g`�y�ib�O�+N S�s/h�۾rJ�M
��w;�#��i��C��,��i��Q6�#�7Nu����=�
>�k�Q�IN�Y�c��2�hN8�3w�Z��_�&K��>�(g(_~�2)kȃ�w��~�e~T��r��9�3��KU�k�(L�Ƴ�Q�0ZH6�_�E��_Y! � !󟞽�]ߪ{kAmX�l�#ծn-�f�=񹇵;}#���Y�ȿ�{�м񤍻�m��1U_V���
6-��:��w���y����D���r�<��V�ςm��F��q���I��{����vRxd�i<���Ep�K�T��S+/f^�U���/���"�9���^M{C}m�ɿ� �Y����H��A��)�+m�K+�s��yDr[N����I�'����"�n��6�U�>$�{��.q���:J������@\6;a���R�kl�v�h䔮_PTd�}u�z]�ȾO5�&�H0�)zu�֙bJ�[�1����� �UY�4�~�&j�g��\��eo�d��ri�j�hn0"ޔ�,�}*�w�0�'�b7�>D��<��pz��j\���� [����3\��U�G<�R�~W�"��v�����m�^2D��h��Y���� K_O��Q�=�
�bVb6e^��5_�t�c-7���~ھ7ɝ��)gc�8�Dq�ܩ��$��D�)7SVX���*������z�6%rk*�f�ގ�=]�;QA���v����xe*�kc������i�C:����Q0���''����:�J�?���_�l�)���
<o�������6Z�6��F>�Jt�t����Y8[���꼛�5ۭ:5�[�	��8�<� ۹ p�����L�P'��N��d�ۛ3�F\��E�YV&�_��*��F�ub�x�L/�n{sarbT�m&:�U��?R��eԦ��V��o�'��X�q>9�ߜ�W�W Z�؉'��P�G\������^��ɩ��Z
���&j+Լ��>1��q%aZ<��	?>���`��sC$�����G��`�o���۳�+]K��z���[LD'L�mū�Bf�7Ʒ �G�'�jl/�n����z����8,�T�)�B�K��K�y�+�=�{��(�c�b��������e��H�$��2+��\�29�
������m�R��s��/ �ٕc?տ��b�'*W��z�?��Ɂ�'t�t�يJ�Ygv��Y�s뫜+ny�C�R�k��H'� �|��9۩�5�4�����ح6�����IE�}+[A7rI#�s_F"K7�QW��&
L�j�ˎ~�-�g�� Kƒ����B��ɘ6��mN���'W���7�](��)�S��9�]$��t�v��&X8�?��^r95d�M�
�����M����gq��v5~�z_�%����6�H�뾦��@���JDz�o��j������@&��#�ɰE���廉�m�[���S��#����:�g�(�� �q��%�~������C�^CbS�{�\L#yS�T�*�Ԝ�v�v��-q`�=]l���β�i����:�  K��x�w�D��/��Or`C���>p�4^�W^ ��
G��Lyv�;W/ ������2�8�F�x�Q4���6�
� 0��X�;~� �{�L���ys�)Ex�*��+�E�������E<7�
��6;��H���!�tN�TNk�r���ޝ����$W�;_qum"�m�]3��|Fˍ�{�pn�l��+����Kf����<�ar�6��u���O�1xm�ny�Hwu���Ϩ��j�Q��sa~��_��
�@7UAT�WhJ�iPj�������u*)�������ɐ��1%��6��'H�Q3ʂx}E�g[�_V���f��-�;J+��?�:F�%��0KQ>�3x_z]&��c�g�㣪���ЛC�Vmk<���+�����lY7��(���4�K&^�d���J��9rڮl1�dZ�椛�ɫ��NI�߉�=
"��U%Y�RY ��x5bjO%�4�9�u�J�e�fPF>6ײ�I���\��	�T��r)�דI��!;n[�����]=�A���ؕ�EoЁ�bu��0�d��5�Uf�6	�{�u�WU.�`�W�T�ҝ]�7��s{�d�r[��	���O�I��,�j�>�qb2�q�0�qc{��ڂ>~���Ͼ����n]�	��l��;K��#jf��m?���pwӂ6+�Y�Q��M�`�a��L���m�� �Z6ifK9���g[b����E?���n�!���Y�F�jd)�[m��EN�)�
e�ۡU�Zy�'Xx	/���9�ك���؃eP.yY�8���'�����U��S#���G.
1�R�/������C��r�SKqʓ�^W�:`vx���2b>�e�%!�2��mE�hE�|����H�Sɱx���F�A^��8ˀqp\��!��c�Ľa/`L��}�=h��6!��S�(Q9�d��(!�v�)y�a6�r��Rƙ\j��PL	���}�a��[��lC�J�c7���Wه&݌�)�;�,��>��t73�"�eb���@��T*+�E�D��qX��~��=�0�ߢ�&�7 �^�GwT>����_��wXS_�-��NTP��H��I@�Ko*(D��Q@��Q�(]Z���B��	%H9���~��{����c?yv����k�5���i�9�e�V���؅���50Bfu
����5��_c�6���^��F˼Y��R��P�6��44u��;�,:i6+JS�{� :qOeɗ�>��>Q�����6��������1}�T�J�
w��=q�B��o�3�W��a��F9��/rz��d��3K�^���HgZ��l���ܻ�'��>�~������+�ݣg�#Z������I�>�敄P"[�L�i��)%���B����~eW^{}��j?����~�]�b�Nr\W<�m��f쑬7�V�w��XyF�����j�P�.��(�p%6�9�h��N���½m���qy��l��H��	ߕ�L��Z��i�Ы�W��gZ�SC:_*ىN7ي�~�g�n��]�0�|N�2x��%��b#��s9o��ǖ�e{���'�l�M+Td��j)�m1���j�9��i�����։�آf�Y��ˉu�3{n{D�>��c���`���j-s���M%�Obǔj\���)*u���`'��8�q��[��Z���j7{QN�Q������>��?B^���9i,1� ���X�h�����*�{n{�C,���;�}x���s�j;b�����f��K�#�?�rO�Q�բ[��ini��JY��v���\�qQݳ�,c]�cǪ��RC��ӟ�\%��
}�����ѯ��CG9t"ۅ�ny�Ƴj��6�D�S��eS@b�Gn�!g�z��-Cf+��"zw�3dy�.����%�����Sk(է	<��RDs+*�s��n������4��Ň�R�D{�n�> ���r��:,/�79U�a�E�L>����`&,��C���>o�*���Z*A��jo������e�e��� xlRH������by��;]%�5�8�%�g���K��9�ܼPk	ϰ�O'>5�@}�a<�Y[^g��T?��|Ǟ֑��J�W\k�9�h��֊�4U��7�ʘ�C'��V�ؒf^tV�o��'�p��	�b�'�������7���X��r����k�[@��n�h��\��wԺ�FCUH@�u<Ө8�{��وB��MڮEN�F�m��S��3Uv�v�0g⃯�J�������}����Əڅڡw���`�X��VۀO����&]�;�b9{@��u��O0E�'�cq��qĶ�k�d�Azd>Ul?�W'OL���E?r�w�����{�O���-X?��=�)��b[�-q#|
2>�;F.�v�#3�����u����8��Sl�jO��1Q6+0�=#�� �|n��~�-7���HAV �������P�E��ә�h�Z���U���ZB�C��Kq�Ԗ��WB֒���*%&�����V=��b�?�k�Q:T�u�3�u�}~��|NEw�C��6�:��{e�V�Et���<�V�D^�x����3�2 �7X[�� 󼹌��H6��W�_��tJ�H�<Ί:�s��O����b�u#��4�s��4n���u�w�b�b_�r<*Cng)����*6y>I#W:�Cx�p���ЄJ�ߡ�����v�7��D��q�'S�|/�j.����s�����Oml�������5����0��I/O?2�<�kۗf�V���y#f]Z�r𵊮��?�ڽF@ך��/w�p�⍈�聘�Ơ��xuE�y�yDQ�9�>2�c���F�Z���Y��N��n+0����㉫�t�U��O�,l�ٗ.s�hL���~�s�&7W��v[Ɲ[7lS,��A��OF���~Z�����%@�v�"A����S�N��J�q�FCyDn7cn�����R_"�δ(j�,FLC̺��ff�&2�Q��b�z�2l����mp�]_�����a|Ik��.QyN9h�I%����^�Sz|N�=v\)�b��e[��ߩN���e�*&�<�}��i�K��A����Ԥ�#�ě�\�ۮ��	X�mn	��=�����@M�'A$9�c��Ҷz��G��L�:X7㚱���2n#�x��C�1A�ebbd�V���l1���U�p<�2^8&�l��t�3�oxQ7��_p)k��r��7�D�zp!��7�nx@�K���<'���g����+��ƻ��K�Nbs:������T��e����0nO���M��a5�|�7�s���t�Cp��~�0Q��l���-wob?c��bߧ�l[�������G��iI�SO_���.��̾�5�ľm��Ix���]	�7nrX��r���#�ۻE��˘W�����پWy� tS���Ocn[��L��zKl���ҳ�س�Hp�����l��ӟ��W��B���*�� �⚒�Z���Z�b����΋A�˯|�oX>r�����/厴�ܫl�[����.v|�l�
[�Q�B�係�S�)��ڰ�0�����9өO�S��\������d�g��=q�Kw��k^��n	��ز'�[��v��n<U�z�ʑ�}����ŉG\��2~~�
k%1�,���|��B+�����K]�l������p�X�H�3V:��;��f�����)�`��E��o2��-zSs��l%��c��+ĥ����W ��V�1���)�̅��J2�T,}ĮS��pϴW�S�>MOKe����c�鯶�!\_��Jj��-3���!�MGC����|0�m�m��K-�6!]"����<�h(�~�#?��>坌婼�Ny^}u�u��sό�`��w�H��'j�iw�5â����;��@0%�a_ދ��/E`@�<�K����c]�կ:0*F?�9� ���T�5��%�H�禑��Vv�R�����~���
}��u��541��9�\���!b��#����]�䞍��*�)�}g�/�5��6Qb8D���6�)(J�zHpƦc�:|�D�L��w.QdG5U� �x�]�yx�dV.�w⨬-��;���4C��W�~����ˊ�E���N|`F�I3�C�a-"�`ڠ�*2F����,$�E�ђD��O�~N;�j`H����ǃn \� U��ȁ���;EB�cj��Sޠ'ix���v�ŭ^���j�����有���ŉh�@'�[X0G��l��*������N�b�����@���)3��,��I{�Z���(+��D�q =tE�׍�ߒ<Rh�M� uL����confy5\�5�����4*퍼�z�mZ�бҬ�̧~�h-�_D6�r9Y��*PtU^��������y�x�0�M%������H"(>���<���,��dJ�f�����0�1L�0y�#}jYRb�`Y�=��Y���Rjڇ��U�׸2�~���;�j��M>�q�t�������#�Q�X�&.H���3��ζ7ѧ�����[5��f�qR�s?��:�9�
N³��>|���ڴ���~�������j�p>NL��@�+	߻��wY6�����̇q�V��&�*B��nu�������g��T$~L`R%$H�z1��4,V	�w*o������3���� �����T��n���\v��Q�W�&*��[����7��:=� {!�_	Nѡ$ʸKe������P�4�N�̷�$~�\�`kx�E����������-�69�d�jz	:rl�u6B9�v�+岁?�%Bp�Kp朸����<pG��������x5l�63�ugXq���7�`�����o�7]���h�ft�V\�,�_k�_뗜"F��f�+C�2�ݥ�eWJ]��#C�7�ř��6b�B`��Ғi>�d�'��ٔ��������Ы�0)�p	��^�����l�E�X�T�YN��TgnJi,�\��r�����0G<��Gi��{JC�NE�wuM��ٛ�02' I�����`TZ>��YN��{ǈ1\��;,���c(�
xVt��
\z�ͬ�����7v��R����t�rhEo>������{��08z�y��F�o�k�gy�>�U���W�QW��՞�U�/K3���2���詥{�W���I�-��U23ե�Z.j1ߓ��\�8=�I���yf�gU�Y��Y������LL��cF��&���:���>lZާ�޸G���G8��(�z��n_P��hBHըDp���왌�n5A�㯟ۮ%�5)n�M��[ޫ��U��֝�Hޞ.�aH��Q�z�i@ƘBYj}\O��mA���"�;���<D���zqM �m�����j�x��W,�sքA�d� C�Y5���+�����5S��' ,u�~i}n!b.����|�KO=�KW쪎΄�R�0�|�	���2w��J���9+Т:e�]��^�ܽX����˲�V@��tʁ6S�r���l{�L��r/�C�y���X�ǻCǥ��5�;,��oD ���ʝ��[G`��)=l���@�՞�ʄ�oA`?�����֕WD�1�Oօ���Kf����Pѕg���I�P���r���hK�nu�Rl�Ke�׳�_كWH�|�P��	��+��bؘz�p:��1�Nː��էy��Ό3��M=�6��Z�����R��j�X���ؤ���i�aS�f�;��fbZ��7C��B����.�Y�\f�hA,��N��S ['��ec5OC�`�����<t����%-75��`�;F�"��'��"��j@�/΃{^�75�bl��T�k�39'���E:��Phx�DTvel�ҹU��[_�l�g�Ar���7���a:�q{�B������a�p\*���,�_o����'�}#�x2c4�ZQ�[xg;���غj�IQ�=�ޖJ5P�gd��+���2�(�~N2ɂ��$H���<�*����m���(��Ǌ˶E���-R�1K$�6mP�E.}D��;�q�V�Ӱg�;P)TX��0	x��C���qRɰ�������@{*[�w}�f���<o���#?�m���:���-��ex }����gq4K�FgE	��?�H���9N���-�5,fn�zL�,,��`4:;�K�R��_�қ��.La{I��Ouc�Ѓ�n�	v�V�T�����A� !��e��BQ]3"��N�J����nX��ubۃ���{����V	���.���yV��!�BWyP�S�=�@r%6Կ�Q�K��.�������O�@��J�h�_���f3�Ui8ӢZ=*����2���8� �CPx�����x~"OE4lk,s�w�Vz�U�Pb��GJ�?Vm��<2t���=�@�0�c�����n[��%�m��G����''.�^�����z�_#>��	�c�̦�c�<��{ꄽ��Dݝ�>�i~��:�?~ں냼#G���~O|=rІYEx�,�kڿP���D��s	d����X��	vc�VV��`k�R����gLk#u�Fz[}����Vd�
&÷��^�P�1�l�_d<�~�}OX��6��+��~t}��5>�(�!yW�-V�m`u�VοV=Q}ܽ�\�,{�}�ȥ8����>��g�p��Gg�2�>�ՄH@�r���;�,��3�-o�IV���6��N�7ݍ�	v���]�60	u�d6IY�8 �iI��Ä+��PI�`�s�{m+X(��!O���ei�����6��'�����)F�)Ԧ	����b�%���v�)�$Ɖ�J�Л%����'�z��{��	��4�/�x��T�,E�zo�f��9;e��UK�9>�c�0Rpv�� �{d���c���]ξIA���n��
�����N�������'G
�O��:��qU�A�UZ�i z���=��č�Q�N�Y��1�5Dp
 /PE������j<3N	%�;�#$Y�i�*� �"�u���q#������/��E���;�ɵ�����D��y���`2�a�^��^ ���Cj��+�y�� �����K���K�9�7SK�=��MW��gK"{vU��j��&V[V+B�q��O�`{��2�ʑ��/�8y1���2��TfA�r�"�Ֆo4�\5x0�zu�ະ|@�iܢ�2ֲ��S�רN��n�����n�$��Z�~s�c�ŗ�xg�8y�&�]��Z�c�W�{�B�k^\V��)=�&]n:+�:9��{K���;�$�駋����5��}�)��W_ȴel�Gu���'�K�|4�z37D��u�mbmԛi��c�=���O�R����9i�NU.�G���_"b�ˤ��^W@��U&��%�[�f�M�*�����չ�B�|!�~pW����ϡ�����8��c��3pFec�/=��0�u�W�bσ�0v�1 ��@3�6���z���-�f�|��ǒ���t���A��2�s�󨶓�6����Q7^##j�i���=�R��]f6I<���������yqgە�Sq��oq�ӾІ�nE��i�(y.���Q�7OIM~��V6�;=$�߯�gzGdm��!蓀Ps��Г#�.����i�<������#B��1שf������t�z�o��]�������P�TF�(xB��qUv�2����{�xJ2.�g��M�աg4ś>rWM�ċ=�а��Y����t��?�8�w���r�B�h��~�	5/�q�Y�]��4X �=C��$G����;�mL_=5ˀ�m�_�l<��aB��pl91-̞�c�����#�8��s"Mu�ڢ>%����4�������3�n>��jV=����$��mi�<7�F�c-R���ݭ#���bDk)�v�C��UO�Vm���r�u�I'*i�{���|���P�zv������?�b_~���|�x�Q��xj�Ќc�H��E(�V��ĳ;')��E�s�]V`8����;]!Rl{�����3�#)���i�M�\�1�ѡ�x�v����l!��,�����m���f��݂ݵ��㒢�=�f��]Y}�_�Uw�UV_P��tT5�#�j�ECjM�v���x7�5�k���u�g$k4;�(L"�dZ�b-��GL��&s-P����8k�U�(�m��_Pz��:�)	����(�9p�#�~Fc��g(�j�7\��V� u�]T�H]n$N������s�F�#���'2����������1Q��C�F��b�2�V���TC�����ۥ��Ɲv��Ŷ�P6�l�9ӏ�>0�u�@�N^�7����
_lG0�� ��������;�y���oE��2��}��ڎŃKEs�@�p����A#��1]=o�:�E���@�JPZu�=7(mP��H�a��x=і��H4�XZ:�Ao�G����#J{~�Sp��핌Z�H����?���˙7�� �!u[Uȟk�}ʕ�����&�b8Va�lq2���2B�*m|I&��cn��K�B,�Yٽݶ����{��h���Uy���5ӛs�}Nߴ�����S�cЍAb��o�j��U{�?�X�i�$�=-a̑��G� g�?{N�h�Z�q�����(A��E�ߊ�_�b2K�TW���ը�ws<5�f�gf����ڽ��cϺ?,b�V�/���7se��E6���K�.����@���JL�,qXLD}X�7�p�T��K���$j57�{.h�<
���gC2�}��BNɤ�Q����.�
���"��tB���N��l��p�-|�d�N1$�o�����5�|����X�E	;���2��9e�6�L�p˹B�u�'F��,��Dz�����3%�Am�{R>(�zvKn�Et��q��.����Xa��
�r��<�zhK3�-'t���r�cȾ�h�np r es�jʴ�S<�%����%��a����)�eb�����M�0S	�/����F��Wf)]O�~V�_Є��G��4�H ��U=�
�yO��i\L^&3�k.�ֹ�{ђcw�z�m6�� I?��l��fvk̱��%pN]�Z;�9 eq����+Յ��]2+��X4[wF��z��;�3��u��I���d�T��g�
z �m�Ȋ�ib]��K��_�������Aj��c�埐�L�����^�����$��:e�c��`�������f��W���f����M��a�>���X���#��A�{Ŏ���>��|~g�"瑛��
hU֯ Ķ�Wm�����ÙC��=���oE�ʁ��*R�'�ئ��`��e�����돻K,�CF�G��cܡ�D�wD�-�W8/4/�\�q��̶��
^����o��|e�_"�'9	��/a-��D=x�"|��t^4[��^8�Np�5p���@S�iKnЖGz8M���T�k���-�ˋA�����M�MMp��?��q_5�i�0�&�Ӗ��w�Lݽ:�ls�9ŏ��c��X���*D����
j�jZ���j� ���¿�o��>/�K6�h;s�tw�����W�_�"rQn�p�e�:����*��]܍r||p ���k�1��ܼW�?��$gϣ�O1��I@)�v7	���s���G�g��]��A�坜�{0�eD�GY�w��}��$K X�W8����δ��&�l�L�\��o�@1�:k +����J���)���4�A�}K�s��ȮRt����VY����޾�i��Z�������q �Q�kO�n~��ϻ�Go��cY^��Km�HԖi�&��G��#�2!��_�u�2��`���\&_󖦞=�vPm*�d��B��m��
�R�y}v��)C���V���,5�V�S^�Q��?}��u ��8��P���~�T�,��7}�4c�D��7�ܶ$XH�?5��U	�Y��(���Ŕκ�TXk�o��{�NG�0�����=8,W��S��^M����	s�*����e�M�t�v~�w�Պ����=�L�Z�s`7��=7����M���58sg'o��>�7�2<��������˼���Qh���7T���"ʜ�:�˲��H�� �5�����;3"BI�@�H�U�R�|�1�ڙ"g���%5Y%d�B���&�F�l�Vb.���8*4a��mH�ǽ�Ŷ~��7������0�u������_��&��|��V�yS�a�,��T���Y���^D���fK�H�vj�,���mk8��O��i��P��A��c�۳k,���JG�p�E�d��4x"��?|��[�3��nw5]����+@��U�%M��Bj��������"�ڳ�$ �n�6?+4��l�9�Y�Jлoя���e1��ѣF��fi��<��,`y�B1��8}�f��M��'Y��f�}��x&v��"��{�lW��۶����(d2vh�[�8*�C�Gn�G�������F'Ȣ���'F�R*�˫�"��N.��{�z�ە5��;E(��}ۺ�f���wA}Pv:7�����8��1��u�3EF
����dTR0u{@햪2S�����'N�x���pbe�����\���h��	���ْ������J�(o�����/�9J$�,����n:�R�Y�>��,��k�/ȸ�ӕ����������q��M�x������1_��Pk߸����O�X��ߴQ2�x��k3U�P�:~3���� S������moV�]�2���I�7h<�$��N�|s��7��Q�Kk�q�u��p @�)�X��J���>ܵ�p��s�Ϩ������C[}}C7H�eǳ�cs���C2}��r�Z�+^H6(�Ŗ�����%��?�j��q�b r?=�Yj�m5�5~�w���]>��⾏V5���V�yq�-6%蕽�%s��3�/%N'I�LcI�~�#�+ɲ=�Kdn���~-�A;շ��hP�7	N������K���<��	��%oH���%��f8�{�c>�ok+k������.�l�8��:��ٿ�rY���f��ш`�O�6��.
�L1��F��T~�)x��ۯ�G�e�in��nǻ}���� �.�D���M7TR���8��`l�H8��W�ݞ�B4��?H��C8W0֬�/ �Fgߝ�ֈ�u�]W�C;d�
�m@VVc�_ѩГ��ߵg�BK!��b��5�3�a�U��q����t��J�sF���uժ�(���o��Č�Ub��+���JYJ�AN���'��!��8��&�6��/xz�<nq�S�8�	��Kȷzo�<a����m{�{�y8����L��/�p��r|r^oN�p�+�^���m�_]��_#����*��uÙ�N���vlZ��ҳy��m�O�O�.7'a�j����#��wk[}݂�	��y�b���,�np�uM������a���P�~�P��:�+C!:�dɉ��s�%�m.�ٱ5��N�K7����4��K��#6mv���j�h��]_�'>u;А��$G'�ɘ�ѣ�!׹��5%K�NmKGV*��v��q����F���dm����𩠋n�uq:�A��O����Pʜ/o4��(HğxS;"�MP�ʹjԻj�r�.���{}׺���G�?�J.Y������P�E�,�TC��CZ\n�~�fh�ʎOC���1�+�Yl��^��i�1��&��a�"*U��\y�lr��y+'������q%6��?����|�W���Z����sY��B�eCS�ϼd�����1c�<2Q��~�P�L����6ʦ�|G�����ڸ��â1���5Ð��`��+���m���7��ͽ��$`!��v!�Yeɂ>�`�=w���_�6B�k�$ ���S�;ԑ�dh�Yh/�E�<	h��|%O8��s�G7�к+1R	�P2�Tl#J���U5I@��¥�c�RƮ�T�H� ֩��W���m�h�wHk�~0UX����e~�Y���j���G�
�$%��T��+����N��>iI�u3W��>;Pp�B�>�U�-�GĊK{[�ʿsW�VWR�Jc0z稵�M���������y��]�����:�������P�`�b�C�\㴘����`FY	�4_����ɋe}�Ӑ5Τ�LϦ���x�ܑBWGmNZ��aZv�VQDN�2����#o���f�QO�!��2�� wp����4���[&{��H��ߎS
��۝/%�S�����ZH����%�JYխ��ś���V^�)H��\���D�8�2qؼs���tK��9���{���:��p�ࢰ�NNoތG�\P�ݠZ��d�zЙ�%>�q�ٔ�:y��O�NM0����;���(�}�wtL���v�MM9/����2����	���M~6��Kß]�*�$v*�MJ��Ժ�|�.JU]$_�U�E�[����G����H��^P��\C$6�(����V����0��KRs�}R`&c_������)˺�(��ɢ2�����s�pl�/������:Q�+�(R��1,"`-�v��H�;/�#"��.Q�����Jhg��[3Wi�lOQ�!Z�Y��ץ����+o�_h){u��R�#�,?��U�?�Fx�������s��l���u�旲�k<�oʻq�ox��kd����'1���A!��Ȑ�M��	jԇ\z2��
Sy2���We��/&W����I�f�����u����F�)�s�Y�m��M��_�5���S�]��e���&ī`�t�3v�� hCn�]ꀥ�*C��hncLdC2)q��\�b�ư5��G���]ٙ�pC�5��'���vI���U�'֟�}J�W|�g�i�
k���׃.�I@{Wߐٖ�H|C��)��B ��Ұ���];�v�B����;���y8K2��� __�D�$WqP=�F�zM�V/e���`gfn_�-q�LH�%��ͦ8�T�B��+�s���ws�EZ�!K���*�{��g�s�����:��6��ŀ��h_��XCz
�pa�x��߂G�5�����w���ܪ��5��u��F��x�|��|��]�C��M[a��[�ՠGN��c���EtE@�Y����^�.m�k	�}�w3>��&��V{�M
d�%S���)3֎l��{%>�h�._�������[3RQ`�ɝ	��k���:Z��ҽ�Vw}T��Eh0��ס
�9�(݊:[��RǝB���[/��%��GU���)�d�+�+����U�f��\�r ����zJ���~�!,�젫{���~�l��F��m���
h^j�d���������M��:o�õ����
���Yc����Q��\ü�w�<��k���i��݌I �R(�/��yK�b�ey�������lG��$`��W���H�T�A�5�_�d�>C.T�Yi��	�F_���@�l��zMc��c��0a������)��̗^(J̵��W�԰��j�����Gn�#�'�[�Zv��Z���_QU���c�(����廐��=	n-[1ß��|1eMtwP��VٴS4�8���,��v��d���jC��g2tI�/3���kA�^��\�/a��� �S�FN�	�4�W���XEؗB�l�,�\��/��_��g���J ��<ps-���i:ed���i�-�����_��O�Ni��A�r�d4�U%�ظL΋_S�r[���Z�6:���+��t�P-�qc��i��Y;w�-Z��x(;'�Q��?��|X���D��W^��ވ��v���a���vX8�x#M"�#�|�	���v�Z��	��"���qB~������
Ad�����8�^���
`�@��i��\�ħ�J���� �>� ̀�
[3��/��EӋ�7��a���z�Z����O"\�*f}[���؄N�YZ*~p@��3�ٴW��[j�l���/҅28/�����3�B���k�+��B�������|z���l6��#�VWPe�b> W���� O���8k���|�X���)&2���Ln�?L��K�8����!W�Nx�٪!�����'Ԅ�z�+C��"�Җy��n<3����<MЙ٠k�d�v&�"$�@�	���^�׊���{�s����
%;�2��Et`��;���c��@!�����Ta�c��v��e�.�CmY�r�Y�^�A�r��:ȖzmP��E�n��p�U�f�&�gI�L�Ȋ;p)�O2��"��n��M�8@�����d��r2![��g��aר���s���߽�)RQ /�63��ɺ73���BO^
��qr�\�t�8;�?��p�I%�Z�L	'�3Z�I�5k�j�X�T1H&��8��;F]�_5��B���$�M�`�,�-(Ϟ��Ta�,�Zs�>�
c!x�0��ķ�DB6� �Ս���>���"J�N/��2�k\;�R$�ֈ/D��Q>�l�a�D�&i�4�:X�D�	�,�C�xJ��{��w`�BC;�_���� �d�U��Ye��sĪNB�MΖ�
��^��۞����b�����J ��y�$d��7��D)`
:�C˸r CA���+t�w��@s:?�ga8{�[B���d��B��>�D'��!�N~I-+�p��˲vl�E0{�3q�JaR���E�A7�a:d�Z�ú��Y����YM�#)"��";����,��	?��]&��/S.�u�2XF"?8�/+?�{rco��f��=��kq#��(�%0X�N�R�Y��]g[��c��]�`E�l�@����	?	�&W��u w�	�jcȏX�ÊM�v�������fʠdg�\�E9
��ݎ9��њ�!�J��h6@�r&��eX�������P���QŎB����wp��뢆�-mt�C�6��gJ�t�[�[�+ݙ���탎������l&;�D.�����~eY��b#�$����>�0����w��5����7���I�lf�x1�xQ�s��XMƘ(���Nh�9�"��s�ԩv[Kj��������+��g@�����k!'@	x-Fyy��>����yX#�ì��	ٶz�\(�@-a��s�5�{y�d�c"�	/��xNZ�Ӥ�i�}r9�7���m�^���S�QQ���	�s9���ؾ�Ѭ�=r����x�]�G}�8� ���	�� v�~[�j*��0��,��~����M���ą�Kt�&5��W��zL��lЃɷl���!@����aPV��� _�
X��l��w	�h~��7�v�%���,�j�i���B�I��]��:��t
	�k5V3}�|7`���� �%�.��V�@yh����?yg�!��W��J�d"���
�6-k�n�Q�y��=\�sWc�huUt_�琀�7�lr���l�� {�@4k�ˬ�Ir�&@�q��9���J���\O�y�vmΖoX�#��G��L�ӎ��]��� �Ye�n㣸�%TV0��ٙ�J��y�O`�|2��Y���''�n��]��x�7+Z�A�&h���˗'k���&r���9<=��� ;	���jX!��{��`�=��/V@���Ó���d_��nÑ�+�I� ��J�O�)�T���J�J�`B��u92z����@����&�jA<Ky���]3���v�(�W���|���Qj7)w����z��o�G����`��D�\Fg�M?��$D��)��;��'�T�0B"��J�<��<�]�akĻS�g%�^��h�;>���e9�Z�� _�>#���	�*ᵜdBYm���E���0 ��Y����6N���+,z/[	���ڳ����J"@��R����M7>�&�PK   �yyX���Z��  f�  /   images/34701e0f-fe0f-4ef5-a5e5-12bda4ce8831.jpg��UT\Q�������$����]��%�[�4Xpwww'��H�������/�=�~[�a}c�=֜oko; yi9i ���x� � ������¿�������������������������������C���O@HH��MLBD@�G@H ��DTDDTLtL��g��pQ�X�"��h�p��q�ކ�
 8D���	�ݿ���QP��q �����!�����5 ."�{N	$|53dZ���/�����Pzns�T4"bR2F&�,<�|���%�JI����khji����[XZY���ٻ�{xzy�|�����INIMK����UXT\򳴬����������c`phxdtl|baqiyeu��������������?��a�p x�������;x�������O�='����>-W0
�����~T:nu(���<=�.�������(��������m�����qb ����dc��\�m��h;�E�2�Z��]�&���`lڙ�$�5�/졝b�I�͊�{������t��[��jT�H�+�6��〈�B ��k�1�n����
�r�قTH�T>�[ �qe���m�"�S��8ޤ �"?�/�zˏ�A�'�[J�����'}Av��8�_.D+�Ǘڔ��+�>>��G�U[Z]٬v���=|�4Qc����?��G�gZ�s�6շ����S7����+YB��z>�Հث�
,�&�ô�y��ʄ�ρC
���A�O�����C��Ѫ�g� �����,M|�����A��o9:�2;�Q�Z���Ҽ������e��1lD��Ξ��V�AOV��5�����hJi>d(qד�.�����;�n�*�T=��[�e��`���\��=�1��}��_���Y>� �\��X�x�R��'<�on[��S��G�E(�e ��9;V2m«���^�V�������Md�?�V����} ��A��n�KI)&p��W�����o&0)?䂵�co�N���É��&��3��I�ab��=��z.ϵG�1�d��=��7@��P�������a|6�)	�a�_�~$�>��(�w�k��&;%$��:QB�s���O���=	/�o �'�וu�B��׶�L͑S�s?SU���� #8.���HU	�Y�0� )�#_�ӂX�ǟ'�/��V��zeWE��H�����*�3�ъ�јQh��'̗8��#�B9w�,�ɾ���,l��TQT����pѯ0~L�����Ǫ!A����:��b����M�KMF���G@��=�,=���xw��Ev&�>��{FԺP�fєjC;�qʿ�#�@��=7�(m�|/j~�р���V�oT�u���z%����,�A��5L_��OnY'w�t��A��e#ު�-����iD�'�a��2z¬N����Ĭ`4W�c��a���d�)s~��g�]� �@��k	rŠ1�]W���!pu� �����k�=�����_��2M��ϒ��{����^E�����q3�Ryl*h�dj���֊�d̷p�����q}� ���I�v?-�����%�NY\M�`8@�D����*G:&(2^����� ���ă��;�^���w~q�
%��VH�ZI&r�\�a�C���U�Fɰ�h闾"� �T�#�����P �׮�3�ĩ�:�7�C����oMd��)��;B�;Z�˝L9�Ў)n�QT\
a��Y�s���}I�`|�\���J!,v��V� ��7��X�5y/�抃ȰJ c5(���=�����薏�ּ\������Ǳ"z��&wc��lɋ|f)E ?��w��@�ͥ�H%^�y����(*9M�]�0@��b���.��>����$���������Ws0I�� `����cܫr��6KiI���t�0b�9I�o1�h�CL�8-�r�����$d����}���_x�:( ����)��spG�E[k -%:��f�p폃oG�~�0��H2`dX�����+����fbv���~�=��������=VՁ������_ti �GB��V�w� <��-ڈ'��^Q��&Q֟���9r�DQ
l�#>��|����Fo �B�!\2х��o�o���<7he������B#f[��3ɏ�D����X*@Ybs�b��~7.��l�z<<���=������5P"p�׮js���iY��Q�� /�&�3�W��DON�-k��`c�2��A��-��C>IM��_q�����S?S�Gh�+�h�v+r��ڐ��un��0z�-o�Iq	�_qs��F3������Y���v0�H���a��q'1���^5��%^�	$4���H,7aZB�3�����Z��v�ɽ��=χּR�	u��F<#������K����U^��`3��}D{R1�C�\�9S���Y���7 �Uj��הI�Cg�A�Y��6�v�j��� mqw�9f�g���:b��N�yq���!��T =n�D�,�ʠ��볤>Ӛ=z�y�?�&<�sH�{�n��Gh8'�ej��`]��]�8�鯑#��:27I�ѣ���H�3����i��\�Pa�tԭT;ѵ�p!΃���t���NF�	^���� �B}�{�c��ӆ�GK[����ӑ|��"	�2Q���߉�Ǳy~�q�S�pf���[��S]��w�b�F��ޜ3i�� � �Ѵ]*B_��Jb���}�LT�+=YF�;�o �gac��E��?�^�^�B/�����g��X2Ǽ�)g8H������ƣɹ�ҟ������uh�srj��Q� ���2�Cg��{�<�x��ˡ�rq�]�f8���2!B�&
r��A[r{ԑ��˵�Hmbx�[�KW�;�t�W��3Z�����*4��|��lh?�\�FE��F�3*o��'̯��m���A����1����Y	,���?�����C�ɚ��F�<�ٌ�����?[ʃ߭L}A��{怟��d��3}}�˅M�݅(���군���խ�Y9ݫ���c��mt��ح����}��gP���K�Hb�A���=@�$�6����K�3�q#m�dH��/^j,HN)���T��C���x� �äo�Ӌ�麷��N�;89J��6[��!�1��%SX���8U�um�DX�㸗YqM�ُs����F��"y�:;�[���_�DS|N{M*s!���M��U�*��V�����;�i2����^�\�2��e���jF��/�pb�{Q�@D���{~o��p��KD�Ъ�.=������tO���a!�J���( f���J=\vX�+����
�k��A�4
*���ʺ�aq�<�r	2ǎit����KN]u���7��ٻ��@��^��s���|��z��Ul���O�)����[;Z����1�w�Z�G!#S�QG��-p�>)\3�� =���rR�L7S�\&�r��KyN5\t>�R�,>�e��2��~�|r��0�+���`>��@�����Ư���S EY$	�|�Qa[��T+�p�8�p�s\wLu�V$�2��O��&��#Qzo��e���Afb\�|�mÐ�d��d�#҇#>���Q�I�-��_EfG��嘇%MS�5wb.~^!�zm�dw�<�%hƟ�c�l��l��̎����vʭ6��C�J�R�Ѝ�hzm#]�����/׆�P�D=#H�3ԉ���2��G��\;�\	��:#VH�-5jx�.�~�:Sc���vR�#�08c����H�-���t��T	�k{< W��M'S��_�Z�DO���4 U��Y��h?lZ��,����\��G�PG�>	=������ԥ����/�=z��O������G�J�,����د3g���Zf'ι�~Xu2�̳H�8�>�8���MZ��H<�HEvf�����m�g��>��p� ᪞���%V�YU��æ������vvB�@٠7�D5�?�S�
s`,� p3�t�s��N�#���PU��sqh����Vl�R|����A�����a�E�.Q�AB��=�i���܉o���y9�t];��,���鸂W�w�����/A*\�����2K�;鴮��ec Q�m�[cn1%�;��4��V�}����,j��}�1ף>2���7x>�� h�� ����;�I G��ڭt�:��aR*|Vy{�����bQ�jmn.��J�4�-?;�`�9�śJ$��_k��]vI����!��f�0�1�C������d���v�c�Y:(ֺ�Nϸ�f��K���uv�
K�L��{�i����j#��q�U9�sa�t��0�n>�;�힋�gˉW�v��[o�D�h߷^֢����@|/Gm�ϐ���VQ}I>N�7:���F���#��t�3�vf8iOD`��� �7Z�����[Ř���̤�E��0�G��]�Y�/��h>2������g��!}y? ?����u��#�q�w�k&t�dx�l?�sz�#�: ���i��G\�	���������}u70Ǵ89�`Sz�*���2B �P��>��V,Q��.�ӼT��촎A
�u��a>	<�$ta�+����Z�KU�����毃S�c���G����'�{�h����z��~�.�"��R>���̐����m�QEcx�r;8�^D�9A�%oKh�@Ѿ����n���y�SvK��G��6̸�T�a�=�:�Ri�^���j�s��a��������[s�`b�4Ø�q��Jb��\�;n��0�X>��PI�,�Uyo'�S���(�uڡ�^�`'e��O��$�;4�d�V-��P�B ���9����)��=;�3vw��?�f#.��j�{!���B��\+y
&F��X����xg�^1��M�KjC���W�1��X�!U�.UN�_oA���i��5���4�����g����H���V��j�g��w%4@�x��!�i�cA���*�3(ɬ�+�6�Od�"���pAS��u.�Q
���K��w��]���7/�w�?�<�Ww��gm�XZR�C�H�恰rs��:J��k��m�̄�4Jm"a�b��Oh)�F�Ӣ9��{mJ���r�3��5D�tt�/��ZP\�N�5��84�j��^C�L���K�߿�i���?m�ǡ�l��9x҂��8e��{FMf�'�u��;��������Ł�mQ��嫕�{����2)lk��
���izx��7z�t��i��c64� ��S�3YQto�'�=����[rBM�~ژS}�m|�M�?2�E����A��Ȅ+��jo� ]*��@?;3��n�E�|�Eݭ������)�_�'��$5g�#?��U%�Fư��3g�"��=��u��MM8RM�~!*\���O�s�
-�Q]������ݡ�@��o�dO�G�[���.�JÓW �1�O��w����2&����1ˊ����9�ݳs�����v�̈���Z�u�;����0IU�/�Ry�k��I�no��L�зG��}���ܦ
G:6t�����e���:���3_{���#	z1�$K|�X��PCta;��0�,�����ᙪ��>¦0��6ST��q�E��H�{ =���X/���ҙ�K����uP[��V�jfR�������=��
���;�*���̹R��PM��|���ׄ�{��Sd>��e/��H�N�6JN_�z~��7�-�_�U����*��!�JwߧX(yˑ�8���,6�o�Q�'��e��1\U)S4Ő������y�kh��IO�Y�eC'*�A4��,�p���ԙTգ������>�x�(� ��L�6BxU�z��Z�JԻ���j�=�S��֊���5�z�j�s��Q�	@�	 8� <Ȳ�s���S �ʹђ�?G��B�ڗ?x�tXi�p��8Z.rf9�3�O�VZ
�sypyЩk�mk~�Ԗ�Mo,X�݀aO�z�v^�m���8^�lZ7)��F&��ᐼl���,�H�$4�u2��b�SY6Y���n�F�aｻ��޲��u� ���'Ǳ��Kۍ8�qփ�+�ަ��	9� GX��U���/S��-�̜{�F��5�ڂ��l THM�PN�t�8Ol��
3]���"�?�%���1����4�)g�j��Xw�c��6pL�i�����:H�e�q�8�	���R^�4�%r�����"�,�����}/>��܁�@�'[Wĩ�Ž�]t������e�"����2\7���u1���n�K_v#��3�Lx����*"�	0�����e���
\0��`��~�t�Ԁ�6F^QA���B��-�0#�n�^n��u���GԿ*�As���4W�	�ĉ������
����:}��W驔81l�f����eI���!�wA�Y�P��������Ir1�kM�kU1�)R�;n�6�E����z%t*�lJTV�Qz& �>��Ԏ�@X�"#�Ţ��77�8y4��r��eL	�	�/0�}��_�{�K�����a��_6N��~$�� �u~��V��LH�2�����Ϳ��(��z��C�.J3�t�DҘ8Φ�O�τ�$�ǌ���^��[X�"�N[�8����<J��0��6?=߶��v'��&1�\(Y�a~���_���`�,�ۀA�~b,|EͅV�^EU���.u����(��$6a`i6q&� �����?��N����P���7Ya1�e�]��ٸ�ׄ0�5f�:�<���Ei,��ǏS癴Z/^+��?��N'��َ��cO}���-v F��c&�1?��C�د�
0ϡ|x!F�T����(l�U�% 95'���;a�ю}�� ���l����` G����%I�ٜ{�o`d����p�hCj�#�O&��n���^'#�����P�s�Ǘ%��>�AE�=��yɴ��[�J��D�	���~k2�G���溥��K_\B��*��eM P#<���s��èI��ϣ\����nX� ��<���8��@q���DPk�.��oM�|{HZ3M��U�)�X$R�{��t9�f��=�5A��'a:U}���w�<B��w�������c.`e�DR���>"Y�1��X!֮�͠���X��2q��C�<�U�����"s�B���<��7p9�������k��$���I僰��`�bT{%�ޟ:V��Q:�;�4�(v<,v5x}Z���8��idǿ��NݬY�J�����kޔ�|�+n��װY��m���$Mj�6�d�L��CCiz;���SE!܉:�H.j�3�׽M�q�0~/8��ZY�t�0Fc0����P�e>��ы�Ci�␉cǺR]��o,�厤Ii���Jt��X�����\��U��.�u.�uE2!.�?��s0j�mH*4�[���xr����B�#��जp�c���!�ôt9yA3Z`ߌ��m�ѧ)��V
M�9!9¡��ݺ!q��|~<�v���V�� �tD��V���±��� f�q�}�I0� ��wm��9�Tk�66�L�K��a�+��ì_ �B�"��N���@��K�F�J��.DV[L�{�Z3` ���%���S]&���G>���k<Ч����?*�~t�01�%��3�U�������cp�!|����,$T�n��=�L�M�?��S�O���Y��I�_�4�v�H)�G.DزN�n�B-h������������MI�g�v�{T��~`̺v�����8���"���%����j �;t7=���$+eR��)W1�㽢�'�����&B������/�
��$���1D�?��+�A�灚��؞�ޢ��>�Dw%Hs�F�F�����e��!I>If����)�����j�o/�y�w���/��A���k5d�zI�f]��##�6L�nUR���1O��_�(���G^�!Ӓr��*��x}�7pt�e��c�8��O� 5Yu�M���F����n��iw�
�Ͳ5N���[�uU�B]p��ʻM@�$����+y��P�״٭�3����1Q�$j$�.��d�H;��?G�-��s�,P	d�ŒC�*�'��V�-�}Q$��=ja�}� �]6b�]�W?��Zb�:X7�B6�f��x[��zR��,?Ho7�3M��Q5��b��^S��8L�^�si��s�?}�R' �pC9շ_�d��1:�K��'�[��� ~�}��o��ِ�8�Q=H�6J(5ѕ����h�Ѓ���^.�4�p�i-�65�}��i$����/g�=,����p�sj�	��#���w/����� 2�>q��7��hK�/����~t�|�Gk������!�^��J�V�/�Q����"j�Q\i�2v*�[�p�:�h�R�o����$�c�� ��VA���ĶGx��OR��S!�ZQ>��81 �Uy��2&0�oS�0���쯮����i4yhx�@�`w�Y������L��gدz�S#p��d�-ϡ�,�"�)�����
��ß���2��놁X�J�+n�Y�z�|iO�F%��s,��I�O4�N,����%:=�_ZۏWו��yS��k���Z����A�3s�'�"'Ox<��&W�
>@�1T�4N��Y���aT�ɫ�!Μ1�~ɤA�3�.�Al�9/�{�Ŝ�&Fܔm��{�*`�ã�(]��=7m>�g
ؖ�J'2�܃BW� �>��U^�:���\��#��7\��(V���9���3�������m|��<��Xd�³юo�l}ӑ����F<*�,��x��YR:�ͅ��4�Q���Ձm;�:c�����Ɩ�yI�a�ߕt夈H�Xa�ࣞ��Q!��}�:��Ґ�ס��~WM8QP;�f*H�A�Iޓ��aw�� s��\�e�T\>�Z�2�+�e0��O����J�2K��q�wJ�XQ��ם8�x��"��bc9�3��=j!�%`�����g%���k���H*��AD&�czh�sK�Qd����]&mRMɒ>3�dX��DT��� ���6�h�˿�7��I�}��֘/zQw�t������:�便���G�~,~�0�-o��Bu?�f��=på��fE'��.	��6�o{�l�9S�Ǫ<9�h��ޏ�*Ѳ�ﬧB��:Z��uY9�6Kc�Zp_��V<�(w���?�QI��Ow4�x�����/#
���Ah{��D�9���ua@�~S�5��(�����k�3i�g��	?��}����Y�'Qj��b���y�ZxMEDO�$�~ǔ�ESv'͎��������.?;{"t��]��U@�A������Bz�@�� �l�2�=�}��P�B����|���K�'L�I�Ž�����U�����t�B\��B�5��	6��^���|�v&��'�6�.w���=�h�\�p�Ι�{�WQ��ݑw���-_�z�K!"-i�_,���C�-�h�J$��︨yL���X}~<~��P��֫J/k��
�hC���Խ'Nz�O寁�Ǒ&N���2��}��9.�]B���=�=מq�����<i���k�hC%Cp7\$��@��?�!�7���݁w�&t{8�~�T��'����E��ff�n.��+�n��nPW��-�$'�b�'��s�;(Fʳ	?�/]���:�;���4K�eIIuԘ�WM�dE�������_����/i�Y��WV�pO'$~�U�����u�f�9��bJ7�Iv���䖅`r���}�ƒ}�VFoOQ�}qM"���}�O_�s�B��t�Ɉy#�I����*ۗ!��x����o�d�%5�6|�>�6�����C��$0�8h��B�%�Y�
�FW�{7'Ɗ�>_����@�m;ϻ���Xم��,9B~.T�w(���Z6N�<��?/�_�<�pӏ�?�]2�Q�vK��-�u@�4T�:��� ���:�0��/6oz����� ޮ%:��H�=.$O~L�P���}}�	ui~��{�lۇ�����;���w�0���� �[C�܃�;ql�w�]�G�«��u=�"l�6�y���2a��%�!��Aj��-<�ި.T �8�}��aAv�0ؗjD�U���_L��6���Kcۺ���Ѳ�CƯj`'h�� �6�,����ŋ��Z�J��g,=.2u�ߒ˳�}�lR¼{�w���e��UX�0ݾE���$i1.�f�2r�Z��Ѓ��t1�.X��՞%�x�d&�,�d2%&�"g�BB�o�cpե��J�_�ې��Y&���F��XJ3���5�����)�T�q�e
fOE�YRr��%:S�Ho�V�P�K�9�M\�f���m�����Ÿ���Fð�Ծ*C�گ��d�g63̊c�?3�90�.H��I�JƦE� �bq��_�q��M!�RE࿹���S�
���rAp�1}�����_ �� ��o���7��r��`M[9ַtf���'�Z|q
���\��Ҙ$�}�-�$k��*� ��}f��0QN,S�d����Y*��3]^���~�V��5͖���Oq�F෥�L�̥��k�b��tH���#����~��u+hFy1Q�;G�ˈM��L-h&��M�:��+��&���SltmQ�N�@�2S]���Q�*�����l��ل�i��Ș��ǒ�<j�̆%AG���q[�ʞ�n�����r���������gZ�CuAN��XW���B����|7*i���+�
�3aߞg����;���e�!>~$Z�a�[�c�n��,��-�<H���������:�b�g�GE&A�0P胳+��
x�.��hu���'-q��>�Q�&��F��-�y2و̭@����7@�v��^%Q�� ��V�PG�� ��9+ž�_���
 93f����T?�Sne8�L�D���Zfd��)6��2E��O�!�=4����ݝM�F۶��OOO��p���*qc�JS���B w~|����ml���*�ѐ߸�[�jk���7=�t�t:�y�v�	]��y"�:1�A$͋�ՙ	���{缍[mwbGFM�ǝk5�&<�귴�_��I*փ�� �x���n~tGBL��gL��Қ#�\<:�����r?�kw��vP���$���$���Ʃ8 q��Ͼ�l&-�Z4ٽ��������H�	�yjl�'�^ţ{kL�0/�H�0e�+�,(FH8�H>;��*�XV!����2���'����j su��o��.n��ވ
�;�d�D��->J郼��AM�=͘k=b-�=�c�}�֥<.=v~ҬQA~��Ctlfe"�U�^JwkA��]^�&붻�
>|٥S?Q�W?Ҿ�'d�L
Y� O�� X���2;���{�7|+7Ӕ9�M�:���ϙb�����~R���[���;�|ǃ���v{��!'��V�C�Ln�hܸ��/�f(}b����W2&���UK� {Q�r�`�L?���M�m ^�"�}?�e�������|��u�������6�_�J��O�V3�RCI�LA ɺ�w��N�}�U�U�-�7 ~͏�x�D8E�]�|�s�f�n��]���\oCf��Q��3�u��Ͱ8������j��pS��W��	sE3�y����L���K�/������x��<ai���[�5����A�]�Y���l�y�J^�Mj�mN��+d:ބ��\�=�8�­��3���;�t�D0[8�VL2�+������u��!���Xm�U~��ϼ��|t��q��Cp�Q�z|\���|�H�z�����	�����3����$+a����멲�9,��g}��15̂8ʃU	iV+[��m��}��WV]	b�7��F.);!�`�����%噅��)���/*�/�ٚ��J�!���Q�<���I����Ou�ƛ���8G[��Ғ2��N&g��m��ߋ����=�e���m</m3��,p���)�j��u׽��0L������v�?ܒ��s��ﲞ��%�����KJn`�W⊜�-���ſ�@�tf�B��r���ua͐�>�Ģ���]=���T���{m��N�s1�[1s/3)��������,{�R��G�}��of����艕�~Q	�����s��pB��
��
+�O�(x�>:�`��B�g�N�0��9^	WMWϝ>��(��|r���6��l�0eSD��7�&��C%��:ے��'�N?YO��+;�<k`��j!�.��K�l���U���{#�)�oqKPnn��.�_~�6P�`!	"���I��V��u�n`ձR�����zQ��W�6�} ��2�x��B���A �s񮾜�9���g]a��J7� 1����xp�Y)ָ}�#�Rm�q�D��$���h����ǣ���;��?o ��Fʗ�!��T����\eikQ�p�j:.B���S�:"^Q`f{*�~z�~�-^d�5�2��a��B�Vq� >�[,ӿ��q5�%�O��@uv�fnD.kӭm����ٌܬ8�ܩ��I���S[��	�E����9¦��X����&v�~(��ѽ����e�y�X:i�`�^֖�v�$�����#�!�ih_;���J�G�;��RNƅd&/��}ğ��� ��/D�w�-��������H�掤?0���(I��T��m�衷�#Wa[�ݰ����	P�P�W� )����T-��B���)�e��4�R�ׅj8�E��<8��D=���*�|��@ӕe9�!Q�ްA:HY��^a��r��|dXN�����,7��$�ګ8%bM@�终HR��}�q��Ld`�wr�~����WB�t�w�R�a����=Z�8��D���q��d������@e���mժ�/���,V&و	w������E)��x�3_D;�;�Ծ�|kf���Ä�����U���>�`˷	ټd��=�p_���[8����aR��Ŀ{1���A0s1�[�%��X�����K-Ίʝrx&Ԛ�:hko��"̣����?b�GOS;E�M�VNY Or��[�JiD�� 7}p�m�Q��È�Nn�W���k��:o<��S�(G�j�R��ܮ��
���"b�� v���5������ �/����f�oF]P9��12A�"S.�/�����@P��͘��al�t|�q�z�	;S�w�#��$~C� B�9?���W�g1��޴�����tO� U%�&ny�ac���)��/�d�5+�ܶZ��LQ|o!%��?2L;q��~�pŲwJ�ơ)W��ʸ�e*��,i�UJ~��7�������wz�V2�Վ�ω˕C4ȃZR�S��Ȇ�aJ�w�O$,�R30R*���6MA*�	��3�g�ae�wMF8 ����7���FΟ�Ë���G�PǏ�d;e�)�b�C��f.&�)��~�)TnKX����I�����Zn�������&ܞD���؜n�D��s�\��^c��_�E3E����\$K�n�3pq(�KK5G˻\o ;%��{��v�y|�9G ���%�4R"�;Z-��a��w�~a=�_ ���FX3���JD�E�1�iU~�8�|0�_�Z��<*���IY��xt9p��.��ga�Ԩ��"a�ǭ�N���$W�eK�i�F����gTʳ�k���\b5�����u^ǔc�|�	�]�NE%y��m<�~���a�S}�����/e�/��*��ءK�[+�
-���_�XϦ�7@�_��7�haR���r`�\�p�U��m}��c]��%4Ggڵ�nAF�<#��J�M&��*�u���"��̹5���~
��p��j^�ċ.T��iK��H�m@'��3��/�~���%�J��y,�Ac���5L��T��J)���t�˙�=M��ڙ�-�v��A�.�ë�4K���$35��	��u�>�82*��kE4�m�uD���2h��%ƼsI�M�*��-=N*";F��[#f��ř<��Z1�-�L�o~1b�)��a҄!?	L�u����nF�����K��� Zlc�H��?j~|!_�C��5��U=�Ƭ��Y�]�Ϧ�8jJ��3�O�z�R߇ �������*�")is7mr�U���:��z�*��x���l&���<sNX3���j7�����v�9T���9���@x����Z)�R���1Q�E�RV*ϖ��07_F�VV��*ADɼ(fqZ�i��=K⪡�6��m[Ձt�s%ԇ�o ���^�&��^v����d�������L��j8��~�]�'�7���� �cm>UCD��L����T�Az��w����D�����d�Ƈ~:��i�sd��{����z���!���!vm
ޖ�\F�cC�� 0g?��r����~A�+�i����F��a�v�/��Xڨm�e�����E �8.�3n���\7Q̿}��US�\�"Ǹ���o
~�Lh����;3$n���Ɓ;�㾱�6L���W�LF�k������6]?�Օ�s�^�"S���A�I�� �m�]?�k�O*��H(������q�y_y���=��P-���O��9lʉ?����=Y�1������-���K�n������w��N�IGUU�V��z*ES*L��D)�����WDơ���陃���!�N9Kͧ��'�:Xz�u�M�
���^鷄`cCfmJG��g>�L-HC����@`f���^�|\�/�C��{�]���] �v?��<�&�+ʄ3N�О�vG�A��7@D�AT��۴��]2D&�,g��
���4'���y�cb��$�c����7��Ηknl�JG��i�+��C��:�s���L�]-A0)T�|�/E��Kɀ]�e��\�tyH�����KTr!w��X�m���f�:���ץX	#��3�LV��N%�MO.Nj�:r~��r��Ez�=��/oTxW�_{Jo_d���(��a&s�!��\����T}[Y>q��V��#=L�^j"��Nє����}�4� �X �������l�bL��քi3�n퍕��OX�*w�K��L��)j�=�}�߷�w?�O��؅��M�>���$|i��0�����ނ-(8�K���6���lds*t�|/����s��ۋ�phn���0W�;1��ˏԪ&W��3r�뼓�W^�]2o�i`��i��sm�2��ذD��f�fǐ�h����t��w�`58�Ǚh��u�븢/1���b
������EX�A�+z1����y�|��y~m�߼s:L����i���`��췸m|�]'\��^��t�.�X��eqL8憣�9&�,�Ԕ�`%��4:�1YG��9��ۣ�1�Ot%��Q:�c�|R|�o��H������Sq�r�<��Rj~a
������!u[㱬)N��Y���>m�.�.��e�g!w�%��5�_���^�OR5[E{�,}�;yW{Xaֳʖbv��<�~��G�t���K`�`/� �k�r��lt�-`5Dҟ�6���!�h�&@@��R����)s��G�+d��GDECù���G��dcF����"���Z��To����¿�r�F���*d�7�Y�ͿFzO�섕O��״
+zџ�`������t �&�93��ݖ�7��h�����*�P�߳d�^�~�{��� �QVs���	�d)������Xˍ�����ݙ����i�g��� �i���5�H�Ө��u�mȋ�&��޺��?�Z;D�q�\cd	�-ش���+�
1��z�u�Xz&���X��~�W?��k�����]Z�>�Bap�J{�0��L�!�_ՠ��ڲ��uPe�m��'�ǹX?��|N�eL
� /l�y��e\��k �Xl���Q�a��+�	L�zFC}w#C�A�L�e��k���퍍S�j����!�,�[8�P҃c�
cT�L���{��_�����=965�F�XA�w5"O�]�� ��]����A��A�,Ib���-���]&D��~_�ݩ�����|P�����bl߻�R�&-9C�\%�aǃ��f����	w��|`{�UTz��j�z(R�ᦸz�����@� ���t1��#�.;�@�@�$�*W�Px뻂M��_g��q��{Z�RK5%��n��%�.l�c���$ؗ}Ζ���4!���_
(�5���P�Xp��V����(�Ӊ7-6; ;�s+`���ܘF<�AN՟r>}e�$�1�ͶӢ͈��-=���"�q�QN���-�D�l$Uf#.u�.#��A��]�w~�0�|lw_�kG���_=�f��v�2q#[�V���:��
we>\���_c�oG߽R�~s*����-���U]v8�G��R�qָx߉��#-��䰍��|Ļ�Mɱ7cq���ϳ��'d�M���)@ֿ6�r~���_"^��ֶ��ͭ��guq!�n�;�<Y����'��5��� �@RKAu�kuhw�RYg*AfQ��s��S�����Լw�6�I����2E��f(e�	
<�'yw-�\�vGZ�/��EO�m�"��(�T�ږ�k��:U���l�)��J춇�<��d�0	<k�-��;��ִ{u6�u�ƌu����b��[\I#4��w�7c�Z�������Yٴ_��ͩ�pAs� �Ŏ�x7���y�wS�Եe�� �-�*c��@r�V�Z!Q����r0Y�J���|;�4�R�M{;�����_>�?u��<Q9� �=a���"��{G{C�%i,�u�N�ω���5���]1��)��W�9U� Y��g���l.���lQ�F(�D�s��0��q�n1�k�������O«�S�B�ǽuf�UU������3֪/��>����v�}Y�_ǿ��ǋ�𾡭���<?u�ܮ����5��o�`J��B�$6H�7�|q�h��Zx����$k���?e60ltܝ�J�ڻp@�/�J׼�[xro���̂{][M� KMJ2�2��C�98�w�;י|8�G�|A��� _��?Z�3C,�3��|���H���[;p�+�Zǟ�֥F�斝����a��'��uyu{�V�Z[��H��Ȉ$���}��YwF@��
�o�<K��]i�������-���3����N��[xUn<E�U�|1����S�ö�%���գ6�g�x�
��O���Uς���k� �֙��Z��m� ��P7�H����ڢ@�T��cy'��֦�u��IK����٫[w{.��!����#��е8���h�+a��@�G\���}�e?b�1���� �+�ώ��ߴƑ���z"��;�9>�q_X����X[�a^wD�+IK�Ȧ���q�U{��W;���B��s�S֡~�d�U�c�ŝ��V�<���o�7.�05�\)�۶���r=�r�)�t���yu9kl� ����|F�v��P�����
�z�A��{n=>���Ģ������� 	=�A� |W��0MBC�y��[�V�7«P���� ���{� �^(��iڇ�-��˫x�Z�w�klI@G����'
�p2����ytf�͞�%�h�&�-��W� ��X�@���ǎnkд?�7����j�v��v�e�����\\+D��M�7�ю��F}/Yז��w�ھ�a{��p���@=KU��������ҔT����BP\�v����|U�N���@��K\�ψ����{�}BG��v�gh`�GF �}E��9���<q���χ~�tPf���%���F(≭���ݑ�]d�䉰@����<��+�������4�{�ꏆ� o�f�O�ӥ��/�d���oS&�����FU��G8���L4_��� 5}�xꭦ~�6򋗷����3&I��m�`~PGl����7� ��� ߋ��Z��}~���6$��I.JF�Ȼ[Dpp��H�&����ke4k.J�̑�?�0\�7\���M\�C�F�ZC=�{�s@��~��%A�RW �j	#�Tq��ۢ��A�f�0C&�Y[q�:��w�R��7`�Y�0M��򳜬j�c.9�#;�#򢷗��p$X�6k��{|�U9��������H�L>e�A�o9-�=�r30�A�v����I�;(��c3�U�>d�~\�vV�a�n*H��2�8lb2K����l�d���0R�h�\nwp�'�!�#������O*Y��&w�h����Ҿa��{eD��℀Z��;�
��Ĝ�� /8�}1��Mn�<�y���gq@��v��9%��zc5ψ�<L���ھ��G��~Ϻů�������:t3�v�0���;�H#R�嶖~I���/Ο>�^	�zm��{�O��������r�*�$��n��s_I���π4��~�MOU�i��/&�S3ym$���P�Gd c�3�ǋ�Ή����n��(-�⼎�����#6�hӀd|�`��p9#u+&tP�Q�T�ӷ����E���,�m�.a%g����6��sǸ�4����uلXͪL�����ϑ��Nd'���u~(���όZ��O2����M-�������/  {㚏�?|w�k�6�!�u�صh"{}�B��F�nFV�	U� �A���tZ�����ǎ<I��:�Ƒ8T[�l��w#����(P�ya��'���Κ����?����u���T�&"=�������04�-��|Y�Z�R��7�?��T�*9Fu�a��68�_L�+^�����֚����"�/�Ou��Q�(A;�w
��Y<��m]�yupէ78Ui>���&�/������V�<-u��J�����@�hb��I�F&4=�1��x������f�ת����q�k�"e�ЗD����u$�k�g�ޱ�۝GA���p��}��Zj���O�X<�tP"AT|m�.~�9�>"=狠���t�Դɧ[��]��`�1M"B�����a�6k�N�����ny�J���	� w^�_3��^�Լ5�%�ћ|@��1�I9;�>��y�m-o4�m��DdMҁ�u�~0sZ$b�A�E"Y!@�X�8lnq�q�]-��kqjٝ��K6\��NI����d��~�N�N[�Guu������S%��۶A1H��0�2�� ����><���W�|}i^�X�u��!�c]�mV�*D���C`��|������*�m,U�	n�r�K��3��^ya�sھ�h<Gc��=;F�TًY�5?�J�-w$V�Cop������[�b��JIX�sם�M?+k���i����Z� �d�4�Ym��g��	 �H���P��ۙ�gv����?�ɪ�wI��.����ަm&��[�w���[c�.��N����:G�}2�T��/.�+inm�Yu(���8$$�^D"1*YAS�=rZ�,|-�����ޥ��6���%��7j�?uxF;�
1ɬ���?=�R�<\�N/�[G�� #����*��:n�֚����#��]FSh��d)�pfV(c*� s7�hj�.�ե���5�[Nm/Rt�U�jSr/��]����a�Z}���Z�G36��m���,Z=>3�XX�>� ?�����mU�~��.�����a��O�l#�4򑕆�78,I8s1&�u����Y�j�EA9=4�7<%�����Ѯ-l�ou�o%`��4��J�}�l��- 	���;y��+����4�__.��{�sG�ɂ�������z
���x����(	w��i!X�wM���om��r �$t�0 P�?�T�=Ů�i<��+���m��w���ג?B��2�8T�Es���wZ����%���Okjo��oor�7��p�H%�9�p�<�Ak����� ��S<0_��kg�߆q�E'�hT���C���D�U�f1�0�I�eܤd������^]�G|q��O���D���$���F���f
��>���3�E$��$kk+�ړQ՞'�O�F�Ɓk��> I���t�M��Q�$KX�"��̀`�m'm�W!�x2��j�a𧉯��%��^����(a�p�i���m��1��	�Zf�]�e�V�����c��^G"Y>B�FY�.9U}���x9-���q�o��n[�'ɲ�b�������f��!p6��� k���|�D|t���1oƚ��m��ly��/ �;�>���4�if�_Zϧ.����H�գ\�B[��|��.H�4�F��_d��ah��U�( ��` 1_����a�_�w����櫫�[��Ig"A<ӸP�	3J� �\� }�����mF_�6���3p�L,��
�T�9 �1�T"��G��ҧJ�Qwww}w��jD�d$]Iu��4�g�H���W��P���h.�涚N�;<lY�O8@L���7�c�7u���:�3�M�^j���X��-��oF�c�T�@��DerXȿ:� ��+��6x��V8�F��z����l��5�ǐ\ b�2烴�I�&���V3�ZR�U�=�➫�Ox�_���t�ė��Dq�$�jWQ.Qlm�J���/�ˆ�v�9ajK�mu��6���j�4�+}WI6C���$�q�@zv2x'�ڋj�1��gy�^��T�ג:ȎA0��:�/�����������Ɗ��x��h�@�\�+q��U��\��S{S��8����Omm��5�SF��:W��Ka�y�a}s��-��d;�g1�emBe�7����|R��>2��g�i�?l����t��XA�AQ��aw�$8�P�����X�/.��������4�&�X\�_&%g
�s��*���|�蟴����z~��լk?���C�n1�������J���,MEzq�����/�u�^��^3�a�O�p��}n��T�����;X���<(v`@a�I�V�o:��� x�ps�A�K������i}��5����n�4��>)�.Q����� ��E}mq��Q�y
�9�5�(8���sT�8F�Z�`�z-�w��+/y�!K	bY��Q�v���Z�1�V�Oz�r�P�uc�i��]�,/[��8��IPOj�n]*��d�)�6�%kD2.v�f�#��jI�i:��rϦ���Y��u�.��Ƕw�>��I��Y�.2H�G�J�տk_�Z%��� o�JG��=�:�ޮ�y�����z6���K�	^��A�]6��Q���v�lG*�6����W�jM"�JF���ֿ?���v��?X_xCD���U��Mo5��du��οB�k�FI��[�)S��7��>��c��W��oip��嬓,�.�0��JWixd�#�*ÆW?'ÿ\Z� g���~mbZ��k�ty�����ڱ�h�1|���4�ox�Y�ǥhv�J ��Am���^I f����/���5=�����Ρu��%�kE�aI'�����~S]�RQn/C���q �e���h��e����}����C-���Ǜ4��p
��Z�f_Lב����~1[G�t�</�M��Z�X����2WwT�������s���3ͫ	�N3��ޯ�o�!e�Mթ>�]��G6�0��F:�;W�_ڟ���Wo� �W�_�PF���������̏�D'�*ͷ,�_�%�z�ξt� ��H� �����յ}�Q?@����˞6[xg��&�6��qrH� #b�r2� ���I���E0΁Q��p�.û`by�FA4�%���V-��5�_9V';��
ry�S�aq漆b ���S����v������w�/�n�K���b�thH%�ݜ!$��s��Mh�տu�n������dy���~f�s� �85f����$�sN������Њ܆$��8�K��[�P���yR�) ʃ%s���2q��&���Y[��QhCM�
F�;J���}+�o�FH�uk+���-��sp�1+�t�YNI�a�9�M�XUe�N��7O2<�sb9��|��~���,彳��� �n5W1�2�1�G̒#�'5����[XI8�������}���k>
�5)m��u�ᆻ�fk���6�U^92������Oƿ4�/��q��=ޣv6�drY�2�q�.�䌟{���?�Ӵo�����\Gw��ۤ�}?ڝdo09��QX�;�'�Oڟ�>��s�Y��<m�Etح�L��I�G������d|��$�4V�/vnz�� ����
�>5�<+�_�]���|��:i%�@�H;��N�T��	��W���
i�����H�����A���c!�
p $� k�����i$2��V-�]X)����*���G�B/��;�͉��?/�����S���>��w��g�6�<qg��s�\}���}	h��f 	��8=�ߚ��������Ꭹ4�e�����vY�H؄$a�>��+����=���%�wU�Р�o��F�E��fR�wM�Y�?�'�}Q���><��.�k\?4� xrX���y���3��.Dʇ�G�T�w(�0HÖ���V�P�IT��l��U�/��4�3�> �� �|�Kf֓�aiQ���U�갷�w+K��^�^��3�ee� ��o��G$�zt�V�gb���G��FV��a��3�ڟ����7�q�Z����{�N����I-��v��i?��I��z=k�5��^:�׭|H~3x��:O�5�ߛ!� �C�L�vn)���⹥8sZM�|��Oi�^��4��K��ks�?��I��%��m��y�vC�W�s����x�d��y���]��b��l�A���]o�5��C�zTw]��;ى=H����Zߴ����pd�3eI�#�?��k����}�b���<3�����Q�����E�BP��v�`��ˎI�1_RK������jv�Y��_������8�8�8����F���v~\��p��$.X��� �� 0�<W��W�ߊz���A�� ���Kkb�swР�vQ��vy�X� �p\dgQs���G��a�T���&����ohV>���|=���P��Л�nb���ɶ<
"b���
w�G�t����U�͹hf���K�$L.W��[�溿�{RѮm��j�6���>���A��d%b�M%w!�seRJ�k���`Ҡ����n�Դ�A�䌶���%�@�Ը�.2y�3��=%ʏ��t1�7&��f��<5=���Ӵ�˭*6���G�g�,���Uޤ�#�R�Vl�_W| ���[��\M⩠������_�ܐ3����@��V�/�no<~&�W�n�`�y)��m��@���y�S�9�|�{"�6��ZF6>�'�~�N51����&��fA�]e�M�2�F�펝��_~�� ����x�����N�n?�5?٫�3��g�G�1R�,r���7Ȍ=�q\׍�]��6��׈u�������g���G^Fc�Pr��tѦՓ>�Zjϔ� e_�ߴօ�3�>+K]SPY(�5	f�Ȑa�(�;.U�
ׇ��>�CּU���equn4	�L�-༂_6����v�A,�xp9\���Ş*��<]�^[��G�]��,�W/�bȇ�'�5�=��p����w��L�`��)�g����*������?T<�¾.�5[��:�Lo]�zu�2[B��i�gF�<cv���&�?�Z=��2�����(4�;y5Vh�]'�����G�PK�q�쓓�_�Z���U�Ko���]kR{pM��Ԧ����P���:z
n��-E�[�j�r�G��P�$Pr��$�x�_*�g,i�s����<�м��j1ʞ{�R�X.Q����h�����-#A%O���_�~��6��Ū�#Q�n"����ZJ$Ky�ѭ����B�MyO�� ���_��C��b��������=@BۚB�C��ǀw(9�� ~Ҟ;O�zj��Ք~�;�6;���h�`ť.Рc�]q�N9�\������02���'f�ﶿ#�_��c��ߴ�.0]�Zv�|�xz��H���
��B�1��@&�A�UߋtKR����N��V�r_\C���G��Iu��Sv�˷��<s��]��w�7ڃ*�I�pB� )U v�f���� x�^!𾏫�m�x��MRŭ!�.]�#�.�����94r�=y`�J��G�Mv��g��v:��|iuh/-�5�6�K�g���z�Cz�1�d(�C�_ym��ڃ�W� 4��/���#ʾԭ�E�1�;��0��@��^O��_��X�%���r���^c[D��18t��\� � 0 W�h� �/��|Z�u�[�6�k�P��Fۄ�%����eq��0Ζ
p�����})c�������;K��� զ��+Ĳ����gg��/�e���g������|I���CL��|-c��M�vmgo�%�Ӥ���d[������#rpp��?�r�Z�ߟM��uԭu�F�ur<FIv��Ն�<�t�^[�7��|�V�V��m����im���j��7�i�we�b�&X�݌( ��y���<��ԧ&�������� j��e��B�<M��8`2Ǿz{W����MQI� ��_�_��M���� ��`�in�.�+ F���_`�%Ω�& �z1�^^�9Z\Ђ�a4)"|�ӥe_i��FU���
�J�٘���Y��wdr)��g����\ӷD�}��k��q�;o"_ܨ9��k�u(�մ�.zF~�k�񕉒�S�#<�c'��S��V��x����&�U$o��с����_�36/�'����� ���`�(۷�zq�{	�k�{���� �>c�s]0�4�N���=�y���S�a֮� ������J����l�;����d�$�
�cwz/5!�������7�P�f����
��NA?1���O x���O���=�ub�n��Cw�I�~�{ir�n#_�i#p�F���SA�����4Ӿ!îCn���Z%ܗ3?�!13�$��8l�5���Aǐ�<�K��g�}��^���k��"��׺N�ýţ�+!���v��8� �^����:�+�~x+�:ǋ"���(}�W��};@�Z_6M6�^{��߿tB�;C9'q��- cǷ_¸+˚m����U�7����T��,P������.�G�ʽ�8ba��G-���y�ط� ���� ��� �U�O��7ǫA$�o�#Z{End�+ �2FpK2+�_"���� �E�{4?��0_���9�����d6߆�H�n�K1�prW:���Kh��X�i�+�	l����w�� $��\[޴pA-��&+$;^6�"|�9#�%OR��~M�}���rH@_�gwmV8 ���A�x�v3��w�9�k�ؙn�!#p �;�
�<) n ��/�4�Em�	,MT��7���wM���O�F��X��&�a�H$��#s1 g�W�+�j���7�%�ڣH2�+�
������OY�'�-�>���[��Ǹ�0]�B�$2������c��P��d-.�o,���0�o�a��e� �s_*�[-��Ֆ;�\�O<��8
{�9U,	lA_T��2��1�\iC^jhX��1m9�9�a\���M���'*x)�;�~g���ƭ�;-kCҴ	��i�nt����{��^�I�X������g����i>�ÿ�?�x�D�BҬ�,�eK��$���bb�N�����r��C'�|Y��'�ڦ����	O��-��ZE#y8�F.
�>vgm��t�����%αa�^x�9B�h��Z[|�Q
�6�lc��߆5!)��p���E���_[�W�|4��5������	�*�L��l`������8Լi���B֮<7�Y�O��Q��0�l)lB�3Ҽ}uH|;o=���0e�*��ۺgr1֩�jV���0ڑ��.	� 㝽q۵v��k�� :�ϳ�	[I��io�-[[�ne��O���D��j�I���b�°�u��4��]���.���r��0����}��
�(�6���(Ƿ$�A�|�@�캤ς|D�{X��cY�'d���*�I# �}���r�񎓮k���}:�.b���2$�x��o��N8�YT�efϟ��Yu
ΝWiu��'G�kz���Oa����,���2j�uҵ�YV7S�2!DDۻ.�0ܒm}}�J���L���(�u�jq],��� �+=1��Rf�I� 9��[i����<A��i|e���3��;�fh�K �i�I'��G�H�V-��ei��s��~v�J��_�E��fV�ҧ���st���8}�[q'nT��ݛ�-�
�V���v�}/���>�?L��nb�ڳ�f�|��v��S���+��X�a�V��I_`�,7g,s��<v�9
�.;����2�$�/n���� ��sN��U� ��rJ�������%�������J�o-o<Q��,ծ �0ڹ|nx<�@k�1����qx��Ż%�J����܉�;e a�J�aT��~{xWឌu++f�R�k��5�i��,0���X���o�?f�uMTh��(X�B^6tI��#bʢa�J�CI<�ܧ1$���#j���7/N�q��,��;+�_𶕣j��N����pw��I.��3���dg�@_t���� f��|@�� h���	����KV" p��q�C�[�����[?xjM�C��Ӥ��]J�Ģ��*JґF>]�U�m�{��xp�UΗk�=?r�f��M����R�2�^[5k_usd�US�����rrb�NsJэ��=�Edx��w��3�뺳��M��{�� /�s�9'�z��}vȃ�2�<	���oZ��z}������*"��P2�������U�����n9lb�c����l��G`H{�3���������[�o��tk������L�����-�}�L� ���L��,%���?O%����t�'�M��궗�g}80,�1�4 ��32�S@!�H=k*�r�V��gڵ�*T]����]����K��,�����qN���.|�]�#��?Z�`�l�7�RGV#�H8${f��#]� �3����l}�?�z��8���ϥO4rC�>� 	l`���>�fK�ͮ������27C�=���QM�ɜ,�6�d��v�6>���f]�v��WT�5:[k�Ka�/(�͎�;���<�8�0��>i_h�#P����m�k���1+� 
�<���Jܯ��t�˩��p3�O�Ҽ�
)0?����ݶ��/���Y?!�1��|�$���?/B3�ۊ�#�߻9 �2i�T�,��1QI"ڱ-�n���9�:�^�&����;[*03�������⮀�+��'�6�s��~<b�8f�bU��0�'���8������R���يf 	��~�3mE�^e.\V�3�sP���*�n�ѡ��&��3�B�nN:ׁ�/S�<?�S��Ν6��iwCL�_�~�i,�cO(���f!r(�{䖫�p�Xف�`��޹�gö�.泍��J�=�Q^_3���~�a]V�I��t��+����ik�5_���N�-o!���O�(c���b����7Bg�ŕ��{�x="�9���]xN�8d��-�M��hT�:
_�E�w%�C�b^O��ꗲ�_��~�E����'�!�Ye(����]�����Ǟx>���E'�!�FH�o|?���� 2�e�Ik�ȿ�&�Q P�|$�� +��</�5y�;��C��m� c�������<nZ��˫9ۏ�_.[sx���X�U�K`�q�e�2_�_/!+7��0qi.-7�;�^��f��F�¿�(��t�xN��#YB��Ȋ���{ԯf�Ɍq�'$���͞[�+⯉|q�j�}*y�'��խr�[��#`��Y՟qFl}܌l?���<�� ����x+��L�W���m�=�Cn�e]jebTP���6�v���=k��h~�n�/Ý����n'�*�L|���:xzN)�}���Bms������ZƓ<�2���L ��c����Z����H?ښg��M�L�YrT�3�0���k嘭�OYm�1�Գ?x���8^X��
�
��H�T5��#}�"���[8>j#|�u	�RkO�R�uga���cM��>&�E���Jr�b�W�H8G� WY��ٞ*m�:���{k;xķo��$�I�ڙ峜r�rI�|�iIy���%�����-�7�w��Î���ȫ��N�KǷ�R�l�q��;@8�(l`�偃��}��C��7}�=3�G�mC�o�#ֵ�a�崷[8?��<�X�9	#g#̏h�@��5�y�� �1k�� �z�qy��2xc��t�9��R��W�$n^�0���h��~O����R��B1��4d��7b��l҂���1*�ޤaCd7q�r)�f���Ũ3� �+'�����dez��9I�y��_c�ˊH�D��xެ �8��*�Ьd�_��L��p ez.U98���4��n�D�֗��Dp&���F{�э����*��f�`X��DPm�c`Hɴ�������Ʋ�C<YO{#�d�� Kǀ2J��玝H�%������Ջ(���h����.Uv�\�2p:T��wn���R�-�~�0�����X����}[�$r��#�t�����1_���	's־T����QK��c�(�*I\�� 8Nrx���3� H����Y7jz���w��I<����a\��zmx��T���l�ej�x&՘��N������ �*����:���T�I-��e]̣p�Ǳ<Z��i��� g{���/�bF� y�7�$!w��2~�8���lu�Bk�]D\O}$Ф@. .W�l͉Lp�0?����[�h��
wu"���s���_�b�-��zw���X���l���c���|��G�ԅ�]�l�������|/'�m�,��p`�gܓ|�0�9��=��<k�]GC�薒��
��=�� ��ϝ��11�.���Q���}��w�c%�����J� 	�Z|4��M�Ĳ�5ē�&�ߌ&��m5��L�+����t��u��t������� �3�a��M~���� ���d���R|�wo���_��t5�WR]BБo6�p�������#�\(ɯ��Mα��e�Z�fd�O���e��(
<8�D�kmei
���nR�h���.�M�VI��n�*S�*�#T�;�\`�K�>���4��,muy/.5MP�|��L�qi�y%�vH�O�c
���>�C1��UҾ���s����^���g�F1�d��z���?�mG��ir4��9��X�����>��i�[i֑[���y,�%�d��� �*s�<�ݮ���
-�;(ff݌�=wn���;{�	sX�*��r�Ksc�K)C$/$�*�r����G#�����/W����ן>#��l�P��Kr7��0s��2��p��~]�5-.�ĺ:�$V���+<���|�'�y�k�/�� ����������Z_�{j֑On��F�"3�,�1��X�r���Q��<��5��웲��ߪ+xB�����-W\���([X�k��<�geg�^8�1q��C�p��χ7��o��ڞO?�����m��-4��.ү�k��_@V1[�)`�7�Xg��껈�W�� ��-���k��ɳ-��<��>����\�F5�ůݾ��t�E�M��pk�?h������G�K���+ֽ%���Y��ʌח��z��?�cc%�%��T��m#�$��KBr�dd����dT��~����|+�(~˪�����\>�-��[͚��Y���b�)�`6.�Mp��+u���ܛ�~I�]y1���`�ki�򙔁č��f
��z������=$���1� �r�f�xvY�%��+{��R��PPZC��N��6U\�>I����Z1�����L�`��58I):��)�V��g$rq�ߧ�h0���O�^��?���;����c�I�DV�y�mF��̒H�ي�^<���ж+զ��?e8f`ڗ���'k������c=6?N��UhƧt~u\kQ]Z�22D��$���J#n�#�0G_N��4~����6���3���zz��{~��?�?��P���|�N������ ���'�t�� �W��_�|m|-g���T�-��#�)�1��G ��5�G�OV����5;9fD�����H-�h�~�o��o�5��kM{\�����O��x��8Z/-b�cUتF�'�\D?|�J�~𾙬]�S��k�����E8	5Ǚ�W�N�G5����)�R�(Uļ4�N�h|���m9_A�Kr�qn#�&*`h$E�����	#���?L~�I� ��{��F��7��U$�K� ��u��1,C����^Ǻ�?7`�yf��˩����߳� ?,`iU.�FH��c%���k�� ��>u�렁�ib�_4��<�_�� ���v���[�iṻ������"��H9<�ʥ������V��`��h��$���OÚ^�p���f1��ڠMĦ��l>` �9Q�A����ƦheM�<�@ϧ8������0ry��^l}�v~-C5�S�}��_�mc��"��'��3+�9�c��cn��ʐFy�mI��a��)��bnnݛ�+�^��0�9'5n
^_N�
63��D޹V'�1�=�Zǟ@��T�z��>O)���ա�#)nd���)zG�[����·�ƴ��S�鶿��a?��Kjk�������1��ΰ˵�yl+�E_�#����Ү�!����U��~lV����L.6;2�6��h<����(퍶�g����ܐ�>B�l�1��ܞI��OkY�f�fWxI�������,�({NeK�����hzf�q��#��Xl�1��Q #I���*���9~����mf]7L�֥��^�I���%����аRY��7zZw>��#W{D�d��#1۲ gY�Fʬ8>�{W�7C�K�5+k��΍�$a]YY��)��銴ڒn&�R���P�o�|ϟ� o.;x<%��q<wz��TeN�"��D�y
CpI�xɯ�~�m3nu���I*��ם��<t}p>����[[�����n!M[����$��;�sҾ\�e����l緒Ya�=������d<� ױM�c������ӚV��L�ky?��@(k���ۆP#$��Q�5�b��y�fU��������b�<�7)�����kC�)�M�a���8�����0�3�Fj�ݺAe-�m\�H.d�DNr����Rr>^�z���
�Z�[�ż�	�K�t��9GBF@�8���U���{�V��s:�IcL�J�X�d�vd��;Բ[L�[����֭skq��L�yFD$grg��v��s�����%�
cv�
(~@�
ۆ��F�j���]��hl��4k�W���	&��`\�s��H=s����� ��a� ���7X�����H�I������jȥ�D@���c%q��+� έ� A_���� ��dcHe��/:b�1��G|�&OO�Ha���K��.��pe��`��1u��|�NNH�r��80��k�;��S� �u�N�ʜ�A�-�q˗���f���az�$���$|���4��j�=����Ō�3I���m�.�d��<To-�Ȏֳʅ�g�x� !�v���.Hl61�ݷ"O��Cu2�&Q2����\��@ʒ��� 
�[X>�"8�,�m�ݤ$2]U��J���G�@�P���&��q\�*J��cb�+�ʌ?l�$�}y�I$�ӛ�X�mgV)"}�ʹ<����k��܂��X�F`R�/���N6m|d����M��{#$iΨƣnִ���	�k�������'����
�|a7��B�mm��2B��o:�I���n'��m|A�� 
��N��]�k�f[�����8."W
eߐ�Ic�ȣ �Q]�� Y�C�����5�.�>�m�ǧ��������q�!a-ۄ## Տړ�X�ׂ�^��j�'����[���W�E��fd1��)瑃��-�ݏ/��]F��l�]�k��8�V����߄�/V��!m��y,XrҺ��- eF� W�p�g�MR�,��茖�����GٙGǡ#��z�����A����Gǯ=j���ӣ	�Y#^�����֮J� ���Or�M:�R�E�� �>��M�̑�<I�2 � �Xu�Lyu�����r].��Y M���=>C���e�{��W���C8*��A�z��z_�� �χ��w�/<}�^�wJ}1c���7��sq*�#r>o/2I��3�J��O�7m4�߫;MS�^:����� Q���R�WE�1�?pF�5�ꟳ��p���|#
+���ZB��LC9���]����M�5� ;��O"i��W���G
�l��	 �KtS����'�5/��m֧u-��ҳ�O#9I�+��J�)��;t2�R��7;]� ����7|:���ԼY�iڈ�t3B+�F�|�1���
�>~�����<S��2i�[y�<?�je��#�2F��	�F�a��s� �[]S�[KYn��9d�KF0s�ε�}�����;���k؅{Vz�Z���'�嵏q�>��Q�4V�mե��"O�/�o�i����+�J϶3@wϚ����?��5-�>�m�-�Q۴[��M<��΀� c�`9�5�_��P!�y�-���^���@��F��u�pC��zt�].���ʴi&{���^����Y���VLs M@��g�|d���w�^��e,���c��mQl���X�U�W���?j��|��Kt�~k���'�Q���[�Udh�m��J��澋���7��Nm]&���nm��Q��lddu�iP�6��i� �+�p�^�܏���[�u��5���I�:�����qe��*,Wf4IO�� r;��\���闿	�W�Oaks����0���
4�$�<�G��j����_�Q�W�yc�� ��Z��������#9�̋���;V�Ư��5�;�:�>!��]9�a�$
�;��M�@f`�n9�QU*I6����5MJ�MY^"��5L�ߟRsǦ�nq��|?�S�5X�)�1����׌c�Qx���j:ē���W���8�ukrO �c��=9��p������QK�8^.�HZ[���'Kц�#d`pq\R�G�r�(���<s�
�e�5�o��A:;C��ڼ�g�"���H�6�
�d��>��o��.��<qH�-���YK#dy�C������~Z�/�������g��j�/�����>�&��:hv�ɴ��.B��������6jM�����9� �����:�0n�����iR��im��>8�����ȇI�D6A|pK6����3Ҙ��x��� ���0O~s	�M}�ďپ�\.��ԉ���y�U�_�v��%���a擳͍���烎���o����������� ɿ�#��/�q\iy�<;�6��t�^����V8�v��9�s�>�DzR��Z��g������+%�&��s4o+<*c�d���׭�px�QmR� L�m�K�*�U����I��[Im��v��o9r��0�}������2վ��x��~"�t�?�\��H��[����y���o�@�$�+O�c��a���{5�{sY��Vy�֣��Nd�6���݉5�d9��q�N}�Z�|4��>�g�s�l2\neB���B�=q_e��Y�k�>O�K����d,@�ϔO�S?��bG��&VN��&'�.���ϳyK��y���[e�I49���X��}9�9p ������݃�ޅ�kt95/��Z�HV;�F�^����,��� p �}['��D��<Wfs���&a� ����s���� <yu�xs[�S�l�-nlcKci����30ێ�A�z&��i�vi��:���.���6�ic'��xc����Ӭ�Iy�M$���#p�E=��Qb�fE�f�^�1�R�T��۩FS�u8}�;v���������>�M�P��j� }��G�i�_��u�������C����VT�1��Υ��Ƅ�dR�� ,l������U�8�u�;�[+J�I|��K�Q�a�����tW]�Ԛ|��[�w���C����|�v@^�匿�G�0��u]�N�.�m�iL�nVX�Hߝ�[-����I&}
���#.U��� �_s�<'k{�؄դ���K��W��f�.�|�����K����]��m	�	#���3��9ag$Ƿ 1�w1G���/þ��ωn'���9,Q�����D�� �R�������c5��x"�Kց���᷼�7���%�@r���'���� �T�-O/�x���-K^��LÛ���_iم`�y�tw3J��b;~@
���sڸ���Y�u;��[h��R8��mD*�n��p�'�{W���a���>���9��+e�$��͍����q�+�k�����>��>���v��l��]w,� +�AN� ��,��4�Q��6�5ewkv�y���k���ռ?���eH�ΥF�m\l]��ePI���U��$�[Iyy�VD��T.�����F�98������?/UY�-KPyDK!����G#�W�l>����	�h�ktX#b�ǚ	W�w����+^�/���3%�GО�J�+[8��[Kۋ�\[���	,�dc��V �%H'�Bֶ��@Iy|�4L�!(Ő�P-�2)\�`pE5�����K�{�2)Y�ʅC��v��7�9 '8b+MR� ˸/b.�)._̀�_<���C�i@J�PG������α����	�d�
��X?$��/�@o��:f{�RK�R�Vim�E��v
R�˸ ��HN�M��c��D�4]�̒A"-�?p8s�*i�9 2�_f��Y�$��=���W�K)�J��+�q�z�鳵���.#�hu�AT;8nӌ
�����-�P� �v�,o��y<����EB�lʰ�s.�R����s����� n���� �"�� ��35����m�}�6����$&s����1�0ڬ�\]5�� ����ܡL�d\���G�`4􉘪CfLR6�~� ,�� �3��*Fr$`�E�,,�0��42=����<���o�� �H�^K�����QQ�� 6v�9'��03�^e�
Z7m69T��`%1�ԑ�ND����7�X�[q�T*K2��m��c
��H�2ܐ�����&�c�3�Y�#���w7���V�n�F�hw4�dl��V`�W%�y<(]��~�������3ʖ5�R2"�W�<� �S�_#j=��}sx.^Q��A��9RXWx.x��_[~Ō�������段�U@�֐r ����g���T�~h�;�_�ǎ|;��� i�N�Fp8�^��g<R|�*�+3��Ky�v�<��x��S�`�V���iVEط�5�߸Ԉ$zQ�^��nh:e��;�J��̻���β��.�b�G ���C�)� s�� �O���l����P�����$�YY�F�';v�?ƙy�7V�g`UUF�ׯ֞�e��+��F��کn{���'�e�-���Ff0U�=H�z¿�Z�ğkZv�����]+ΚO���� J�����-��i���y�b��I<�	�|��98�9�/��U���ڙ����˫i�e=�fn�\Lc�]��B�p=*�Vh½�));+ĝ�o��y�9.��
̐i�Z��Z@��l��c�|�ⅸ����H�=��Y>�"���n<]�]�2���|MQ�l�+r9�'�#0�'<�0Ѧ��dix����c�$���v�}�x�ܕ�j�|�SΕx�{����Z		YZF$�<�T�������}K�S���1��x�� i���ͳq��z���
ض�4PF��<g������+%�|�k�`�����&���� d�������� ~j_5'���Q%ŷ�<�6ءRN7�`����4�ٛ@��.�t-gJ�-���ou�.���"�s 	��+��e����U*%-?���]<=Z��t>��ǋmn�t���(h�g>���s_d|��-sO��+g����n�ܕ�ON½G�L��]�u�}Z�$��a�[J7"$d�����`q��5��߇���G�f�]Acy�*�!�T���c �k���UG�õu��#��e��W�C�o���[Xd��i�&ght��a$�?.+�u����kS��:�7ZbM��2�U��&� a�w������ؿ�f�csm�KD���Hd���۱�Z"��1_=h[ύ��H�:O��op���VM���=��p�����kVN���[��[�P�,u�v^#�V�⿅�Ƚ���ye�KK�Z�}�cN%n�VS���x���A���b{[Y��0�[چG�m��h#��@y�L�Hk�z�F��V��׍��L��k?���L��%��x��EV�8��� y_�n�?ej���� kh��W���R�j�Z+�XȎ�v<�@�_�R�)��N�gV�Ӧ�w�  ������[���s$��d߀$a�s��##�c�lO r?ƍsi�����(��[���qoy�
X*�ݣ$�1�޻��VG�4��"��]k�����M����ccg�\�s�W?%�I�Pq�,��+~�A)��ar� ���9+ҫ_-�ބ�{���j~�� �-u�KT�o��k˫��lo ��Y�wXb�؈�I�x��1��Tk�< O�,F�r��M8b��3@N3�8��K;Y�O�����h$D�}�k����@�S�m_���|����x�j^�-tgŒ_L8�ry9�i�����|� ��=;�*?$1�#��X�XطF�*
�4W"4`��k��/#M�IFl/����$O�z��y�͹��s�]���?4�V����BO�:�S�Y��_��?�� #�X�v]�*�)�ڪ,�F�3��R�.�.���+=O�ob���+,W��|���������h��I��.�w;y�OӊX�s�J�g�uW����H�[f������o4���Hpca�W>��N]tG^��.~^U}Y�]����0^ķvWQ�W0�r$Fe'��y�fx2��M&KB�ot{��$���q)2y��h؟R��x���.,e� 6�Mf�㐂���Ib��zu�\F�Ox�(6�) �6��*�qI�]&*�t��]+;������X��?���kǒ3x.� %�"ǀĝ��t�<�k�ە�A�kǻ�Z�, �;��ֈ���ɵ�៷\��K{D_�˪�yg E���321\OOz�RK�k}F�g�m:�?&�9�f*�H��(��Kp�h��F+�?�[M�w������6�2Gu7$?حN2Ug-��־N�+��Ħ��ڶ�yL�s8�����sD�F8s^�/�#�l��E�}H�X|�$M�,p�n�+2�FCK+�r1Qۦ�$q���Ύ4��r��ƾj��e d�,��xm���tn�2D����r"�	6�F�X0m�	�s��ײ��n� oY��D�7(�X���i��<�k]Osr�m�ݴ�t_h���Ll���؄h���� )����������7�{�a��� ���.�MF{�%��Aff���r�  �g�cS��<pz�|�Y��mɅ������d��>M���޲~��-3X�4[&�����2�T�ḿ��1��!�M�n8#����������P����m9�>X��C���e;�BF �u'0�~ק��u� ���x��*����T�ۀ��� �sQ��/ّ���e��M����	�#f~N��n-�|ǚI�i[�,�!�BW*p>�
���c��][O����F9����ܽbH�(�Y�����ٲ�H�$@IP0��BIۃ���kG)���^��ʳėH������a��N��6$�1Kna�eb�YQʜ��� �Ad�G�Rk�F�m�� �(\�1���n2	犁��a�|�n� 0wx��$�,<��2�1��@���c%�<�3�AmoVR�%�Ksϡ'$z����#��7$�a#�٦����n6��@������D>��%ڍ�d(�a��Ks�~����
G��4�/��������i^-��i���Ԟ�7�{y���(>b��m��w���W�����c�E���x��ڬ� i�����o<�N�£�G$������W�pK}�鷗\\D��B��w�h,3���=��>!|�E�XCck�E���t�c���z�HN�g��=�M����� ����	��� ��Sjֲ()yla`FպU9ϱ�V�!kvAw �w��������S�y��?�WD�״�1w�m��@��T�ݠa�����KLbZ95K��*.�&�f6� ��柵���� ���k�Z����$�(cY��}I'���~�W�<L|q�]#�v6�?�z�V����h�a�F�㌊�neke��N���o`�>����u�������j�7���ƒ%�$��T�K ' {`�u���\�	����gI����X�_UXn�4۫���A�OmqG4P�#,�@;����kϼe�5Ŗ��]�I1�7 ���/��Ҵ�&��-8���O��n�(璮�������Q�n��6�� �W9B�.����a�TqiʌyOn����xn-]�h������ Ǳ�� �@�X�"H��sϵ`|!��m������C����u�9�����z��=��h� ��N�x�"���ű�kuڂ[<�� �a�)8�-��6I�J�bӴ�M�%�<���BΪY���
XЂk�?��R�ۗ���ψ�2�
�꬧�+�t���]�_c�c�Q�O�XY�(,9��8<��b2���ʴ,�w��=*�B��菪�
�Y�ͯ�|C��-?O�W��G�'lr#�\�3��Gpk��í>�䶾�4�{̛�{+�!�?x���'�^����ۦ�Se�UX)�9�#���>��V��f��饄.��Ι�=:V8�T�{���J�o�����^�ܪ�4>8|��u΋u��ukg������� S;T�uށ@��ϥx����� ���\����J+4P���̏���z��Oڊ��:�ּ?%�L����A��V��׊�[�4ψ���i��6�7Sf[���Ac6I�5�lg��ӟ�nw�]��+
�⤹��J�F�J�}��k�:=q�u})���i�&T�Đ�� �Ԕ*�����R>bEy�<?�^���Z5���Ky��R@5�o�6�>^l��2�^����O�h5�l��K�-��#�8,� '��>�`��^3�}&��~�ut�����;�D\��%-YRE��Tw���Ȉ)U 
�k��p�UZp���|����� �+	��`�fm�������Q�d+s��<u�)>�;�_�4=@�>����dh5	,�-��w�I9j� d�s���q${o	�p#򘞼��ʽ-l~����Y��\�7v���o
�bEw�RF1�~UoŖw��>(�5_��� g]N�kq&1�n��c#8�oZ��u���
��Z�v+�����*�'��=�k��ؿ��ǻ����F�o�����b���� �����q�x�^y�y|l���?E?����]E/7��F䪮:�1\����� ���Z�[���[;�hg�L���2v��$¸�v����|v�������鱹V�J��s;nr�'m�:�~i:��
8�L��ir~'��Y���S*�������;��!�+��x�C�����rKmʫ4������77ß���Ɵ���CÚ��,�TY/䱄?�Y� �'!������@���F������j_��9ФL)�d1��g��^p�4�Y&n2XG��3^�g��;�M����io�j����"��0x�|��ʬ��8�=iJ.�6&�(N+�k�>��{X�/�&S,[�a�F:��ʏQ��Xz�g��U�� 6�o��yf�̉Q0FC8�NּS�+=q��-WR�֏�"{]�C�[lGs��,F8#�"�>��=7[���_����zU��o-�o#�fi�U��˵Td��+ɕr���R�jԗ���������� i�O���is�1�ǨZ�xe��HK����g�x�W��j��U�M�kc[�!��(J	\)8��N+��(����4q���7���ݏ7�;�_WxJh�R���k�z[�Ȯ?��F�8*Pijޣ�P�A������*5��)%�4�4�]�GX�0����*�2y��q��dn;�u ѩ��S�Z�Z5�����<q���`==�McTӱ-�֙csh��FS��s\߉1$�c9k�� CZ���2�/����ќ��v�K��|7�/f�|1��_e��ay��I x��18���p@Q������	>_�>���qᆆ].	ͧ��e݃+e��Ԓk�_�;x[l�}�O�_V�+�8~�#$����� ��UNSk����:���Gk���� 2�� ����� �Ŵa[���*�\3�n@Q�#�Ҽ^���1�vk�6��۶q��M���T^I��F@��+�~9�3S����*��m/D�#�Y�g���r�p�9��c`�X&x����g����z��=.�u��RY���p�B���<�u��z4�թ����
��s:��<#�O�?g����ׄ�!�\}�3ݬ�<Wv�(#%Q�`
�8�@�����<2L���I|�dx����=���i� gԌ�y����u���=����-
/ܶ���c���� 8��7�p��+��� �z���Ds���_Њ+{J.�L��9�
���|��m�&�'Ï�:.��_i�N�u����٣��!o#a�1���>��?����� �+��(M�j_	<m���pu��}"� �nS�YO�_� �%�������� ���N��w;���J�[�e���k�D���0ٖ$��Ѱ�R[.G5ZX�f�Y�kXXm�M6c�H�-�Ğ2FI9�ѫ��ढ़���&����r ]�+���:�p���^nú�B�h�Z�*�X�O��d^z^>�����������v��heRm�L	3wl]�C���ێK�n8�WL�l��GL��L!9�͓ʧp' ����|S�K�]�5���ҵ�"	�ٞxX��h,c�`qڶ4/�o�����A.�a���|A$������n�pӭ^�kٛ<��ӷ��Ű�*�-��&��
�e�G<�ܟ������ c�z.�#���Y�2�������=�׳7�S�ZYV�u�������.�-Ԍd������ �	���]3��j�p�$ښ-���7H�1%���c�a[JPh��L���Ό����O�>���:��}��N��|��5�Ӿf�c�v�*�=\�s~&�`�����5t[i�6�|V�%� ,��;3�tV����;��>;ho5+�%��=��$�'!U��� t�Z:���Z=N�}J�{�u��ss�,n̻�I����p�N\ܽO��*uUNX�{Z�﮶���xާf�x�©�x�[����� /��lM��ͼ��t�/~���J�o>�Z�}>f7�lL�R�������=c�D���f|^�}.=�V�t<�F��cu�����.�tyd�ŭ��23}���?zg�����Gծ��Q�d_������
�;���ȓ��r�����޸�x��o�|P<;���Q�5���L�������� ���猶."r���  ��-�,b/�+,���	9���_;|P�G�X�� .�?�ѯ�� i;m3�6�Z[O~�I����Ef���O�|���ūiN�r5���bƞw�)%�H�%������~G�|f���J?绒?V/�IC&O�aZ	�o��@l�3�3��=�+�+�@���Q���T����X��W��*�Б�����z��;Nm���}*���x ��&%F��=���޾��9����V��ۊ���ᮧ�iS�i�xr��˞�8�E�}��W���/�M�jw����Ax�I�������lm7ݫ^���w�0�%iZ��>L���Tx*�3�n�	)��lW���>9xÂ5�~�g� Q�9�<��I��Ҿ�����>m{Z��>��f�h������ V�h#޼K�D��x+�.���5������Ҡ��i-��Ȓ8s\Bea���T1=뚎e���8�M�e��R�����W?
���KXҮ4�4�g���Y���u�im�B<�,Sv�t*A$1�5�����O���U�Զ��i��&�"H���Q�+�u/h~ ���)��`��t�1��Oqk
�#P]�#�Ņ�0(<��íW�> e���Q��ȭ��=�ZΒ�[dv���q���8� ۆԦ����<L,y���$�Z����������	��熵+'���Csm=���'�F��2R���5�ZW���<+��5u�k+�E-���ʳ[I�m���IPƬ�h,�y8�J�6��SY�>%���7��u#𵞳�è��d�#�cN�ט
��J����_��]!�U�-������;X�E�`'��R��i%Frm���5�7,o#��f-�ҭ�wm[N��/��~��'�>%�zF��[� 6��]ݠ����!�LZE�Y��H�+��s�����w�]���7�&�v�oc�X�}�dh���UYA1�$9�	�{Ω���M�h�k�ϣ�eY�-4˨�ވ�Q%��aURF_�L��w {��|D���~x��A����i�DRy�;��ds4%�
D�Y!9��_YTҒ��zx(�*%Z��v�{z�sv?��$W�<��V�'Q��t�뻁��,�9I.�<bBFbu;��g��|��2�7�Z���7�5�R����p
�'n�����m�ᯇ�]Sᵶ�k�i-��vp���`���!2G0������6|/���~�{x�]{R���<I`.�n�I-��7?42���������Ԧ�Vy��%UZ���˛޻�� q�� �-鿵W�"E���h�eå��+d{Ȁ�����#$���Ρ㏀Z����]?E�ԯ�PMGIK�$��	e��H��zps^�K�{�� ��i�\����<����n���j�E�Ӱgh�ñ���?�� uK�C֗K�m�٪����;I�|����胖 ��2X�*+ssr�s������§�e�k)~��O�a��4�F^����[=��Y^=�J��r�y^s[���^#�5�Ma�E�D�|��&E���0 ,>�$���Oз� �/��^�MΪl�!x���Y��=~�8�K�RXY٫���1�n'��_$����wV#Oѵ6n�]麜�%�i ���ʡ~�#��  d�kz�䍏z������g��S�?���KҵmN��ΉO47m��֡j�yP����	�*�PT�H��>�'Y�>(�6�\艤$����#�&�24���fV�0 �2v����:Β�jv�_[ɦč�f���EYL[XUU*��%N�X_�����ݤ����'�h"�Tt 4+�dn<�;�\��I�4�P�JxH��7��>۟C~݁�Դ�@bF�l����������4�2�Ņ�����fx������k~��� ���З*��T`��I�}5�Kx��Ej#Qª� �b��;#ԣ�KWF2)��ֳ�1ۖ�j,���>�wl�u�h�OQ��>ة��O:����k��d�����?�U�C(�S�d6�C�oZ�.5�ː��?Q�[�n�5͈32�_���5����c&�ύ>;\ƞ��6?dq���?�}_����Y��� :� ?��Mgx����O�+�K;�(����pF3��+��T�n��H�� ��Tyk�P @+XF˕P��NPZ�����9/�Z]̗Z^�eiqy�I��Lؾˋ[{���F���\�l�U�tS�_���E%���ˆ��Q#�#�R͏����ow%�߻fS،���ck��1�ˇ���<��(�{I灜(�V��q�`{W}<C��{�,��q�<�㖦��;�n�;��^C�x��cm�Z!�/��3.T/���#��&����#��Tp�1�UA�<%�fhU��`ͽ��]�F�ܒ���1&��0��Xԛ��rb�rĻ��_�(���W¯4���.�.v��'͐���:�J���o���� ��� ���'��k�m�g�����l��Gx�$�}�+�_��[��:���j�of������>�?U�ծ$ٍ��+���� �M��9�[������f�=K�| U�4���Sض{WEv[�v\�g�j��\6�}�/7�i��M�l��m�W�`{�3���������������ka������iWN�u����7��,��VviQ�b[�žM�g��� h߀0���)�����[�;@[�쵭YD<��NHx����2��O��$��wiv�����O��������&⮭�Ѐ3�����ŷ�<0� tK3�"�`��)�Hf�T��S��޵�}�g�U�?ew�:kY�P�����I2+`� �j� <G�`O�t�A��p���k���-(��E���>�1�Ҹ���
���
F�� �����S��⢒���� 2ޘ�3����VC�}/#��J��X;6x����V�t:g���u���="W�ᕎ	� ��TW�܏\Ԏ��		�*���X��}��+r��[t:�S���� ��� jO�?�95��yQ�8
8���>�\Z���_5�����&f���Ϧ��WA�-W-��K���ᰆ�!{��iڒ�3i�m��r�*J�Ĳ��U��0c�s^�z�.�ib!��O�U��$� �� *�_�Cg�,O���I#\�`��|��'�r=���߈wZn��WJ[���b��d����2�P��JO�ݿ���;Q����=G�j�^�<��8�5���.:|�5�|4����I/Lu��?�3��u.1_WYl�^;Z G5�n�9�'�yΆB�	� �F��m�q�ҭ���O������l��$����i�T��#�U�����zǅ<]�A���2����v��p�{+���� �'�~,���i!�YY�:���Fx�=}k��G����^5�&��@x�~^:g�J�~���^P�nrW���z�*Օ5+%��~�6���?�z�N�,b�7א��-`h�2��c}��@I�!x���-B�J�m;Q��K�\C��<k,O���� ���׋����C�jwZx��X.~�!_2>>V�kտa���g����k6�&�,����o*;up#�sv���1\q�J�!O�r��Z����T�>ڿ"N�w���ᯉژn.�Kif�ޏAsoe.���	�pq��P�#]�?]�4�o�dծ�K�����E��I�\φk[i�&a����� �5�ڜ���#��E�Ht�|S}�x�������;[�,\�ۀo�8��|)�O�4�cE-��	����W�V�!K�i���$*�
0@#�OUcѝ8ԋ���<�\���#xW��x��;oZ����X��Yf�"��	auݱ�%pH;�k_�/�ӭip��5�*85]2Y.|=�mf��p-טd�M��i�yaw,;������>.��=4��-�7������ 
��.���Y�.M�v�<.O��OS�g��;����)�^�Cd���?5~4|t���?�Z��\��i~$U���`��,ۄrcr�\��(h�ubI����5��O���Q��6��xvk�k�#R���w��m�5v��	n1_��2�g�~$x�'���]:E(!� � gk����A�E|g��	�q�-j��?�z�ӥ����뗳GP(�ػ@_�ʂ�/ ��*�ytNǮ�g�:����/�O���Q񆱢ik6�����A&�i-U��&Y#.̬"ۉ<����������%�����f��I	�0��uʮ���z`����'G��u��n5=OOմ�N{k&IH59��I��À���+2���B�D����b!Y��f�ٱv�<5̝
���k��j���9�|~)e�f�N���������|U��_\XiZDMc�x���������d7.@l��C��S��3�M�S���%Ѽ'����mc��1r� |Km�̦6��Pҙ��w�E{ǃ<i����ӭtk�{6s�!9����&�w<�-�^�x��$��x�s:�Z�X�V>mμ����+lI*�5�8���>����y.z�y=����ɾ֮�	�R�>(����Y\�cs7��Cw�6$D����� ��9R3�Wi�|L�����yᨵ+X-�ķoj=���\�lǹI���$�FE<i��������[^Z�ڤ�p�]ɤ�u�%���DR�5$��'��x �#��� go������h��~���Ŋ�xjH#����\])�l]���r����j��+>jN2z�4�_�W���<�^���Kp����H���g�����g�9�h�q�3ĺW�u�� L�J�d6���zM�o��i$� 3�"��Y"���I#D����_ ��t�#C�dK=J�P�_x�缊q(�$(�1#�8����+�->#|f������T����g��Af�r�@�l2K|������HAAۡ�W�bJ�4֗Z_�U���� !�%��/-�H���F�?��۷�~b���
�x_�+b�I�
�rH�4}Os_3~�>���\*����<��㢾��ش}�6� #N�Mݎ-�J򹜠�>v�G*�ٜ�ú q�(�d�.l���2^9���oQ�Fz�u��1)��j���ʧ��b�SǔS���ŗ�-d���K$�Pb< ���wZ����$�4��ԟ��-��f>k�ip�l�\�����X6Ѡv�>_��;h�qgD+�v�}��~6���2i�|�M�	�P��{n��>8�����е�7�鶷/& �^bp=K�+�㎃~�X)��ǧҿD|?l���픝��ֱ�� x�v��5*JIjwԭ��������6|A��y�6L獼Ew����#n�=�t��F'�d����=���o#^�������
�H���H��2m��8���°�:ק�Wֺ�=�-{S��mk������'�n�|q)���9�W�x}�XЧ�����)��N�����^Q��G �흤��k�����\��)B�ׯ�����z��ύz'�� kz����|C��$w	v	V��E��wP�T�q��ײ���l��9p�Բ���]�D�_��j�j�ed�I�Pyd޼|��zF��j�,[t�IN�����F1��S���ӥQJ
�>X� ���]�xw��YL��	��"N�b�#�?7$��}+�?�]���ߍJ��� ��#\x�$���Qa%�E� [����+�o��� �1�߉��oC�q=<
� f����{�3��y������Տ*0+$n����T����nY~�.y%��b��Y�]7�>���V�,m@\(^Y�'	j>� ��5�rݟ��;Gr�������]�xp[����i���^
��*U�?(l
ӱд]/�ڧ�-�� 3Ě�Z����p#LacA�� }z���i���}�i�������.�/�u37T�������>(x_ĺ���0x:-%��8W��VM����rTg��9\��#�T�����y`s
X~T�����!��]������i�����j1B��>�b�7�� }잕``C��=k�h��� �c��_GѴm?T[�)���Ed+0L �<W-��c�O���ǳGo��K��t>^FZڼӴ��خQN�;���8�ھ:ӿj\J���r9,n'�0��4�m��v��̧��y6��<�}���7�Vկ���e���-���,ӄ�� m'�ҹx�7308;N@�\�>>�<c��i�iv�O�n�Y�#a��Z���(�X��q�o�M��dܺ�qp�� �r>�G��^˨��w�cX��UTA@T��y������q�� �E|��J�e�߁�.E�h��4Cki#�m"�rU�,����N�%7h�N�*���M��ԋ�ď�~2�|�dq�<�G�9d<v��9��_��U��Yl��Oc�^��\���@�>�t�� ��8���8o���( �����?ߨ� �_��[� gG��g��2�/���:~&����&����8�����5�x&% w<��|r�db�#9���{�Il����8{s^�b�쉃��k��;�d�0q^���l�)8�z��fz� �?�xWG�$Q�)ֵ(��oq���	o���'�l^ �V�����?���ю�)�r��QҾA�my���f�������'��y��1�3��\�� �=k�XzQ�����݆�6����3��m� ر��&ba�9�k���|I�{y���W� �[V���# �a��`��/������e6�<6V����C�\��'#��1^��$��zU�Ƌ�I���(��F���g�Q��׏W��^iUNj�_����L=ju�Rqj.�gu�ٴ��W���uv��~ �R��Ռe�Ŀ���X���x �LW��3��:�4�5=k^D#D�Ӣ��G�wB�gku�]�<�� n�����������M�T�]Wc�Y30�GN��^b�Z=Þ���j�P��7�Mb��vI���^#q*�J��Vƥ��rq��8�{���l����H��'��M��V����wy�� ^K�g8^�-z���'�g�v�>���^�%Uݱ�0ʝ�����yoį�W�����MJg���=�w:�C|H��5ܥ��۸r�z0�7���� �>�9�׍t+�Ҧ�<�@-��~�hch��]c,���6�r3]4�yn�.��.{�{o�uusob"��{��Q"��1b P��$�5��������� i����c�r.���b\I���.�V���S~�6�c�:W���v��x�M�m.��F�2���NFY�3!8���`�����־~�q��g�Ū�j�����Й�@bN��#Wv���@R1�Q)&�Q��ŬUY`��v�C�n5��tI�?�h/<M8����d�fpd�ɱ�Sb��H�30-_�߳_��4˧��Ҵ�X��D��I�|�NpK�0�1����0� W�� |3�xcǚ֭q�"��~2�����T����G1�v�x0�#9�S��o��Ե�?a��mtkk�wj/ux^v�!bh! ���y��\��3OtNO������Ri�����>���K���<q�V|�!�O���	����kj�&kTԆ���ll�IU`�_����p # 79׮����>�kqq�jP������i&TX����s������hk�|A���h?f��F.�,۔ ��ˍ���=[��ii'��1�a`��vH�ό�<9�]�{i����;�fb�.��;I�e�]�|�[���r#w��8ԣ��D�C,���h5{����~�Tq��=ԭ�������TQ�jzŮ��MgNѢ�'��V���ei|�*ҳp�n@�;(B��7�'±j���<S�+�7÷�\����Q�4�"��cU;N_1�A##�\��������g<�u�`��������`�Övz�u7��RҢѭ�7���4��,�W�e�8��N[#&����m��)�cG�ះ� �"���H��O@�t(.Zᧆ�.<��~��w�w�5���6֐\_YĈ��`�bx��%����m���W���\�i� o��>�v�cq"26J2�8bAV5�&ߺ�>'Ī5�.X�߮��ߴ��������6��N��E��0+J�H��0FM{�m����,�V/ogʤ�R%F#�FT��w�5X��h�a?uuQ����[��E��5{w/����^_�8���u�u�����aꤽ��ɟڪMʤ�� �򨮬����M|	'���FQ?��]m����P���]i�o ���vk��.2���z��{��XJڧ�ϵ�Ehٵ�2�ڡ���⳼U��-�#f�����/�]�$ ]O1�/�xs�Q��5֧=��Q�M��׷ꌽ�\��}S��D}J�������㕚� �1���������q�}�����1ڊl�����a_���5K?��^���m��u5�8��Y�k}�c+�`�g9�E`�K�W��9[���:�������Q�J�.�ך见�/�z�2YJ��4�� �~�����|H� ӯ��t�����z֞G�t��`��+/pB��<k�B�O���;�ԭ�m^��|B-╉Pʝ�m2l��z���/ڋ��RE_���Q)�K��Hܹ#��'ֶ���~.��П��,���M����g�H���c�ㅯh��r�f.����/«�?�Zo��]ycw��k ѴM-��t�����p�����W'���<I�'��q��~YY��VH�x��9(#�[��
P��%s�grGJ��_���sK�x���@�m��F��Ѩ?*�8w�'+��sY�U�NI����I��� �L/a����x�V}B��7^#�����dq�����V� ���� ^��ǟ��m���}/Oi���<L�Cʬ��G�'x%�W#���/���� zo� ��Xy�
'���ԡF4���I����{�?��ͧC�O�	��Me����
Ǽ�<Q����]��5%��'�y�y��5��j9,��˪i��	nдBB�`�������)��?4�TT�����:�7��ڵ8�-��m����	E��pσ�#�>���� i�Z�����ui��gu���7i��E7(^�����O5�jߴ߈�YeOxF�N�s�Hm��u+K����n"Wܸ#��Ȯ+T��g��M%��I�O�M��ǧ^�&��΍�/5�)���ɯn�zn��&y�Nx�������Ty�-��}k��=譬x�Q��=�R3��7@���+د/���l��A^m�b�9�m���+��1a�n�|����1�I�D� ��|?�;_7�J��@+��� [-Dc*d#=?�����ņk��"ai�q��� �Ҏ��c*�OXO
�v��W��i|�d)Z���x�͚֯��3�<+j�8>z���+��ڳMKψ���� g[��ƾ��˸�A���� ���?�f�y�x�Ͷ���� ��0$�c���(���ߗ�Ƶم�W��|I�}��Ou#} C���>/�lO�;�� �W�~Ԫ�|F� u5����6'~ݿ:��M���V�!��5x��~P�Q��G� 	���Y� �Il�?g_�S\��@y �k��~��]4m��,���r~:
$�������\�a�����8��V�c���߷j�5��O�Cs�L��P�G��<1�;B��tƇL�.<45{�H�x$��
+c�@�u'��jh�U�
�cU���n�-k�mi��&b����X�>����v��*��~���߷M�=%�N�3���/�oX���Io�J��X�L�s�rÃ�r1�׵}{�^�xSC��xv�Gѡ8e�M�>^q�:�q��ꖺ���9{��,���Ku�;W�0��Z�.�]�'�o�������F�-g�Q�v<����k���V�*v�v��������om�6���&��N�F��e��Y�.Ծ;�+�9|��D�'�6�������̊[}f	&��K)rIp�C�z� �!��:׈�;s�ri�D�ydO��h�� uAc�U��<E&���!}!��"B�F�%�NG�y�m
1�F�>+k���|֧��8��<��j{�h}7�~�>"��_�u;�+�sM�X��mA��n$h�_ty��A��|�Oᧈ.o�n<-�YŢ�3���\J����"4���_����}���~���@�I`��Lחk��B�ǕV�� u�ǯlg�}���E4~H��4������ 3_��� �2</�������񡽒�O�-��$7fK�U���` Q�6@<Uxz[���.��6���][�-���L�ȫ<��R0�˄l�	�������Ə��>.�%�[��n���j�{	Z71yM�PZ4|��s늮� �'Ĩnur�+�W�/g���#(JŜ�,B�1ڽ6�I-ձ8z��/���[ݭ� ���{��>h_��u��K�6�����K����d 6⯴%�5�|!���ߵ��/��uM
;]
�K��l්d����GX0�	]��+����>%Y|6��m�'��ΐ�=�v�.ahܺ� �.$?3�Ns��Pi�O�}/�zG� �=�����,��&x��#h��2���H��D�R��	��z-�����w���L���}�@�5m/TԤ�2E*0�(�٤(T08�#�+�O��8���m(�5��_���H��9fD!��dn�2���S�� ��{�x��k3x�!�hʬp%�2F�ʇ�]� �Y>9������^��c���̖�Df�#EC��Tl�;����yWS�iԖ;����Uo7w�~K��ӿ�� �]{��'��� ���xs^����ɹ�i-Ɋ�m�Eߵ%8R�r={�/��7�v~�4�_L��Ȏ�E�D�D�{T��~V�ds�a&H��_�����d����B@WD���O����O8�ǦO�G���������V�;o��M���u:ۘ������8�Mh��g�b0��V���z��>�t��]�j�E힕&�z>�,֍q�Uĭ
(2�#(e�[ �$����� ^��ÿ6k��H�j��w�Ŵe6�|�m�c�=�|?y�L��T���m{W�\+��j�!���)��;g�Z�%���k��C�z]ޝk��iwQ]Mq�]\-��D�pʹ�$z�K�IhqR�֣��E>Wm���EY�ⶍa[Y��8��@�x�XZ��������r1�t�Σo��Z��Bx����xՈ�Wr�8�ӊ̸�8�>⸴G�,��:��wW��g�p͋��9�j�֏�t���� Z�	l�r%?��>�&�db1��9�J�%����ٙCbY:����ҩ�V���x��T�\�����k�%ۯ�fja��Vb�S�����KR������'�-~̿��cj:
��ٴ7�[�[�5�d�hG�	ݍ��\��)-��}7C����<Gn��Z�		��@9=Eu�ٗ8�T q�u�������G�$�G9���SN�Ԩ�іɞ]�HE��4IZT1��f��J�,��M��W�t�[��fX��Fm�򲜌���� �b����mq�ߧ�{iU��0&������G?1g�"�]���P�G� ��F���T8$�8�S��������%��p��� ����`;B������#;�Q�H#v1�N����١y-'):I&U�Uu �rA��U�V�m㴕��ȎH\݁��\� T�!R���r�ъ�gpַq�ME���q	-FK�t������n��Op~�m�YX��X"�p�#+�r�P��  ��[6I�X4����q�I1#%�0w��rۈ*j���9�3%��vȡ�"Uն�9Vr�����aa�#�+gv�ڏ>���	
��P$-�$ 0HP��$��Q����l��ĭ�,�[d��8���R� ����'q� �6��E-ݵ����cW�\�y2�I����|��d_� �� �O�;A:���~޾>�����=&�90۽�����$�FO=POۿⅬ�2���7�m?�;��{��` ��9'��K)�[>��b�ـcì���~�����?�R۔󿳰��}��q� �B�-ج���Eد� ���ER�� ���T�C�>���������V��Rw9''r�a{������7��.xa�͎��O��W�E� ga?����������6����GӔ�'�5v?�G���V��֗�j�1n���8M�E%\�
~a�ӵ|�ўz�����o��vK�H���ć�篭eSG��(��`pq�&�+z�g�sx��F١��������iM� ���|?�����f\6q�=j����!j?m�<G�-v��� ���95Ӊ.�1ܐ���v�󏤗����h��O������8�<F������E}�)�XY.of�>m?���]��P� Y� ��d���0O�����q��W�&���
�d���_��S�̥���A��$<G����rt���W���<q��G�XҼE����n*�z:0!���g��Z�$V���#��&�G� ����m)�E�#�����Xq��a���!�{WN�R?A��r�_�2��^�5-;J��:p�i-m���ٞYDm1�哖��᭬m5�����4�3��q��+*rq�����E�nD5��J꒱��� �A�O�5�me�`���$%� 9�zU�+}�Iٛ@W��k��>^�*4M��r�!���E[�B�׮8<����W-*p����h���8,7,�Ϡ>�?���pv��;Ǎ�����|=qo�1��Y�k���-u�k߆�Sc�~�I��t�;]Z�t�J�����\�}����;�c�)'+��Q�E�����k �Ŵ�{�KF����o�X���?�k�������q���� (���(ú���׽���������׹��w���gare���6�r'������>,h������A��# ��� Z�=>��vF1_HZI�÷9 񂸫���L_�(�O�6��*�\��#�����ڄm�mJ�W催����9��|qt��\*\G� ��q�W>-D�x��m�������!�k�.��˟%T��?�n��P�઼\j��-� �x�5u����:~����7�+O~�&���O�y�<W�x���Zٻ��r��pQ��3��ʿ�3^��dx������}�� \W�kJF�`�"P��$����'����L��M/��}�7�J_����>&�4�2�Z���8#'�u���������w�Z�e-�+m\݌�<t�kJ4�he˸u� W���E{��Q���B�}��1���K30^3��K�ƿ2��ǯ�OΛ,P,���<��J�{�� ?��ɴl�N}�ێ��ձ����D�P����6����_�2���`�~S��l��8���\��׀h���������x�0FQ���w|�+�� ������28����Hՙ�q�Z�C1i�ws���0	��J$U�����s�O$�������9Oھ�%c��R2p��Z��`q��~S�}k���׈����Lt�Ƿ�'�͊��S��G�D�Q�6{�B�����U9�nA�N6�~U�Ʋ��v�1���@����Үd7���Gx����wD����Ŷ�s��X�l.�5K�R���o�,�V���M"��L�( s�U<S������#�1I}���}�$#s�A�6鞻�8��8������^����t�x�8����ٔ�(�m(�ߓ=	��y��?W�����*��"��kn���z�#/Ŀ
�'���(}d��T�%k����e��������+`tt8��k�����c�ȴ_����Đ��bG
�h�')�G�%��4�l�;����:=��':��㜲<x̞VrA^I��@�H#i�����/�������ێ�}#䯏֯o�9�7Q��,z�kyB�et���9Q���_,=�"����"�~_td�2/ ��n��C������R7쿥�a�e���������?8 �c����a�E���Ha�k�x�����VC��� 3�U����J�����r�_?�)��a��"i"�;��������(0Sk� |�kbK�f�5	�rϽ���!��RZN�� Fr�i�9��M.؉a#TdfUvV@\s�*��c)��M[x�-�̷+9V�Q૝�2q3cvq��r:Q��'��o,1�k%�R,Fף+	"-�ۋ)����Q�04c���|�Iw<ae����ͽF���"�4���j4Y�����>�<�$H���  �I�l#9TQҥ��=՜3�Ebm����Y���n(ь1^Q��X�!���h�mm#�s"�
``B�p�7#���N
�q���ž� �B� ߋ?�.���u8 ��G�3J���,���;�N�� �/�?�
_��� ����XC�IXof�1�'9�]*	X̋����nܞ�=p>��u_p`aII��1�d�y�Ң��{w?�d�߹ǰ�Tg;@��534�,Ͳ0>���@����T"�̐.d!W%�t����OCZ72�#�J�PG�\�A�c�*	,I�U���hi#<�2s�?\Pa�f�& P��I>��<3� 	%����0��o����RV�����$zW�\0����JU�����:�J����R�Ѵ�j6�N�$�²�*�,�8>��3��c[�g:Q�����G�� ���-���nt������K��eY�E������yb��q��}X�|O��꺵�����k��,�I=}�����ù?k/��Z�l��jńr�\C��;�+4�23(V��ڿ|w�Mᯈ��i�i�%����|�z������mF��~#j�G���l����g�����&<���p��⾱� ��xL�
�k�.�E��5�{�����g%ͳ���O����g��<w�	��0x��?,>!_�I�� I����R#��� ����`+�� l�_L�Ѽ!��;A��%�5��^�k��Cgk��J1�7<�($|��3���ʳ�h�S�'�I�cI�ԼS���H��{�B�j�n�a�HG�$q��g���3÷����lEŭ�-�[��?uU@۞�df������ |�k�I�~������9nF��_��#6�0#9��ڣ�Tӡ�/�Kk�3O�x��d��<Q,s���d�p���lyq�6�D���᪹ek�k�cͼ&�u	�`�b�]������$�>�
��W��t+��9�����ܤ��d�$;W-�x�d���\?��l~\V�zsX�6���%)aT^�>��}<���A��-�5����D�\����?�}>�+XYDq�/��'�j��sۊ�cdqJ�Nǰh�"�9$q��l�oonH�Ny��-~)][�1�^�kN/�Z����2m;�ZwW1tg��s�g��?Z�Me�4�>�rK+L��澍Ҽ+��ᗻ�J����7���V\�p��5��m�����|-�]R�M���D��I\|���^����)v����)�.c���i>���n����v�^%Lf*N^Ξ��%�ݞ�,=8%��d�����^� ������-ɖ�ʀ��2W;��q�1�_?x^	�����<>lʛ����}q^�����D�'�,ń�X<6��(�B���s 3�p3��i����N��J��TE�'+�	�Dx�gS�<����"�7�I>��'ĔiR��N/��u�|��A�?|p>\��x�� ��^_�(�-����R�����nO�;�	�i�%���b�ӥ#�^� �Wu�y*����+G'FR0�~����-�y_����1Qì4峋�����I*�+�-�K��|��v�2(�^+�>��~���s���խ���U�T��	*[Gƶ�eJ�Js�2���_O�� �/|4�95��U�P�����W�	.T@�'�Js��l�ϡ�E.�"*�I�J`���k4W����޿H��վ�Aּ`}v�����d��J��R�ߌ3љ.a$t��SR�c���,�ۡHfa��g�>^O�Q��ϊ�[��e^F�毣>%~��~)x�ú}���2���]�3yo�T H%� �q�k�<{����W63\�e,�	7���"�)�8� ��j�X�f� #��fTg�Z�ow��e�y۰ O#4� �c����=�1Ҿ�� �\_۱����ɇ�v]7������	m��x��+�n�I#���~��s#�Z�cTR|¿.��+���^&�p�X�"o_VB=�?�}Z��J�I�<�_��[��w��/��1|�4��x�m^xuH���[�\�v�͓�l��9n�T�K���̪Ɔ�Y����t 7�q�¦F\�?�������w#��w,ɕRNW�9>���^_��I6쿯�z���� �l��AߓcywW���[��'����t@q���ĺ�"����yY5(�/��u� �P�[��ɶ��N�h��C#Z��� ��y�Ϟ�����{����=�.�ʯ*s����]ߟe�}/�?�F���E���ɱ�=�M��U�չ�$�Q���rMy'�S�6�k�o|8�h�� ��u]Mm�Qy4�8�1,��Y
����?��$��Z�u�[�p�ZI;	�mXm��>S"�Q�ӯ�E� ���ώ�����-{O�j:$�v���pD/'˜�e�+��R�3�W��B�WBpw�_^�������"E�}��rG�u�j�m� �h|Tռi�S:�?n׼={��B$��HD����wM���IP�����о�K��M���ēj�J�`mU�:}��* r	v�}����M��O��a4]nhg�&�rڞ�<s2l���X�P�%�AZ���Э�|�� 	�S�4�"#�[\x��h�ڱ$r�^3�G? 2�u�1������DѤ/V�b���I�y�FP@30$�<Z�o��񥇏��^!��[J���mD�w�K{ń�9��0v�|E�kD�I!Լ���s�`��7nޣ�  3��A�K�G��N�L;���V� ��LʷW6� f����L�H�²e��
�`�\T��~]ū��2���ʵ��Z<;�;�AÍ��K��	�K.#�G!�7��eu�NB;:���wvb�k�mJ�V[�w`�F���P�06ȬF�"��k���#X��C�Coo��L���,�&T��<^�U�,ǧ��BY�̐+39A!�a�9H�"���p �J�'ۢ��5�o�G�r�1F�4���Iv\3D��C @e6�&��Iqq�#���Y!uiSk+Fɂ���(9� �Uk�&���͑?vm�G.��|��I��������D� ��R�5m��\�1���;�t��P���Ʉb��s�~^���}����� ���8���D/0wE;�X��(�U�C��ҪF�FZ�t�;Z3�_�$�=oδZ�9���C�L��c���V=w�ZK�da<Ne�1ܪ��U���z�ΠeT��d�g���.-�R��ŗ�����#��&����������y`Oʹ��<rs�T�ݢG���3o#�O%���01���$���'H59Qs<��w�����ʀ(3���	"c|Q�2>2ۺd��� g8�� �x7H�U�x������X��|��ׅ��ʹp:�D�xP�w8'wL�i��5�?�#Լb.v����e�d�*,���=s�?��;��ut�=�m����f��Vs�J�is���Dl�R�2G�F>d$�p$�|7�A�_���xw\��a�]���٭���v�@99U t�5����iZ��x�����%��k
�Bg�\�E*�L`�p�� |p>��g��^-�U��=�_܀�K����a.yiKϹ@��)�9�ZR�[�X]y�V���k�gw��^h���� ����C|�k��8�� p�㢂w/�����>#���'Q�uHb�c���#��2vƣh��$�I��G�>�{O�}/����h���Zg����9-5ē�qE�~l��%�-=��дy������f%KT,XF��9 � �,pc��i;8�[��8�,UI�tgZ-���h�F���t_�K�eӭ$���D�^��I�\��\[�Q��v6
�<���ֹ����O��7���ē\jJ�Qe�Y��~cE�$2�30F�#ms�i�z����9�A��Z�N��Ot�`V�_%Xl�� þ2�׭<~��x7G�4�ikwy�yڒIo����y�c�T.�N�#m��P������|��|��W�U�Q�j�s��8~��q�P�pH�9=������4�OM1�ȗ,߼��[K"�:e�V� ��]^�Q�6�X�J�R}�9dT.v���o ��F{�_�Z^��O�t��+���HŤ����}A>�p�b0��f�q_?���/��ϫY��͞�7�5դK,�eA���PA#��[����O�:�V�ZE-���+�I��[���& eOpyC�G��Yuk׍Ֆ� �-դ),�����A��5���;������7/u�mOM�	Ķ7+ �V���2��AФ��Ҝ��d����.�u����D���ߠ��q�	d�<����������[Q�}�i:�������:yxnm��Q*Q��?#�{�+W�>��.�w���7�B�O�P����`�L�'~HY+��m�����Ƿ���>&�L��n4�MM�7�?*���A B��<�9�qJ��y��{� ]F������e��$��� ښ��|��yxr"9's(_�89�j�����03O1��>$�;��Y��ڵ�֚��V7p��(Hc����
��6;W/k���*z���5�3[3��bf��h� _3gD�[�\Hi�pA�,c>�{��<%�/�P�Xi^�r�q���w�g��ڼwD�W��q�Yn;|����5�zW�}\��ͤh��~��I�ǳapn+���Z�|�>�įgZ�&�^ߝX���}3��������t�:oّ5gx܋��$/��8 �z�e�|h�Ε�P:��'���|��_��m7K��l���o�ϳ���+q�
@ �ܬc?5r�>�	.��#k�%�����R��g����]:>�6iw���Z�?ę��m#TѼ6dDIM�����2���F2fh�>#iwks.���i2KC�_�ug���|�?Z�O�k����O�0��SRyIaѲ�y�oNް�� 
<iw��/|-���%�̌�t4j�=x=kXJ)$���� �0��Уt�4����w��W�/�w	B�Z�Կ�tO>�������qm�|3��;��NK�yV��D��į���!���Q,=2|��[� x��]�m�Q ��	�yz~��������_ڕ� �6��� ɛ�:gĽNey�O�c�!X�@Qp�$�rI$�NI�3x#�܈Ϭ�Q$����.�ٔ��;dTᯌ��F7>[�[ۂ�q� �=9�y&�� 
��M�5
�� ��&f\�*
c#'ۧj�\�׺������u�[�R����~� β�R����&վ-=��va���\gp!!D\�瞢�Mg�g�a~$����[�r�a$���N���mǉ4KÂ��ܻ	�����G#��/��Z����Lg q�3��+w(� :������Z�� ~��?�LޛH��,	?�!���р珕����V�����KE.��[K�����3\<Me]�b�юrN�3Ҹy�x�{1h�#����zc�S�n>�����)/�^�eV�r�d��BD<��c�����}�5��MҞ.���N;� ��\4O��><]��8뱏���Ӛ4� x�;�%�5�x�' Gk�\M�l�����Ïj�b�G�X�rk~	V |�Hǎ��zsW�O�:Ι,�_�xZYlIy,�$'<���I?]�ڢ
��� �#OOZS�($��s���er?y��ی(��
 �p �=��'���C{�uGPm��$�$`^zV� Z���� 9h�z����*zg qǡ��\|8��#E�<� �F�xY � �8Ǧx%ќ
��Zz��� +�I����-��|%g$2����]�%�A�mc�����0�����w��ĝGDmYb���j_���*-�,�s�C�A$��/>j�6R[Aq�8��7��.p��u�]�+�|6��R��>��6�=v�W��;���C�>:4_)�6/~�;CF}O���t1T�5��6}d���4�"��Z�0��Vw�B��pP3Ҿ}���r����Դ�+E�L7�w���ѓ�ǵWl�FTe�pX�����g�cK��_
��W=ji��w��v g�x����j[�?�|;��>��5��&��㧖A��q�s���\�>�:�*B�/֡�+����;f��r�(䳸�_M��Tm��#A{X�,��
�� y(��K~_Y�$D�ve�Y&+�(L�7ʌ���T��l<����3-�ܐ�zb#����s��S�p�x�k�{���X!mB��UT�ʻ��9�\�B1%w
����,���K�����Y�OԱi�_Yʷ�
���+1Ec�m�A!��e#�ku䭻y����r�n����H�2��F!�~�!��,bM`�pQ����e�7��,p�6��Jz��c���Ӆߛ+�Fg��c<�ݣ�0(˃�z�&փ7ye2E(cl#d�T��ѓq�� R�8r�k������巗�Agbf�B�� *	<��l�$��}�^C4)h���D��(�)$�+Ӌ2jI�� ��	���;N�.DaT�$��#s�Hc���]�f�X��iX�^O*]���.P�Շb:��&�틯��� �z� �a�hSb���+0\�8d��֐ά�x��g$���� �L����j���PK   t~�X���!R  R  /   images/38c30459-3482-47ee-9b33-edd591009797.png Y@���PNG

   IHDR   d   �   �\95   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  Q�IDATx��}`\U��o,3q�&i�TRWjP�[�-���Ylaa�]X`qv�����k��Q�H�4�2�q��9��d&I�I�)��wwK�7�ݹ��{����kN�̋�����yA����/��Z4�����~�`��z�~���xNC��5�h58�����t�5�/ӵ�}��1a&�6blb+:7*;b��!GM�3���J������l3�9�^�9�1d�E�1	�����\k0۱uw�����*�4-~��%FDE80-�9�2ߢ�loJ������b�?Mچ���6����w�$�jI��w��h�v�'��E^Z�����Ȯ�)�1oJ2�~�h2!mJ�,hh��=csq��yH��b��&<��.������f�h���D׬�N�u�`3-��];x�����3cfF�N�V�W�<]6c�8,��+�nƿ��ASW$��F��<�۫P�GIމ:<��D�3�1���F��H;�Q%���
bz0��� &ƀ'.��3��{��pރ�an.G���z����2��JB\r.�:2��{�_V�k_܊�N��{M\x^4?�N�HK�ƿp�,.]��y�:R�-`�%�l�����b|�>��i�&ZO�.��8�O>e�YL�� flk��
n㛨���m�S"���]�/�'#X,�������1B|1GG(��DFj$�$.��-AL��aһ0�D�������4&&7+	$���(|s�\؜Zw��Z7��Zddء���[���-���u��73�ĕs��Cq�QE�ioE�Ѓ'%c|N,��a+�_G}{PR��qS#�l.ڹIp�d�-N��ю#r*@��ť�~^�d���ߦ�H�M�yokL���0���b1�;�����\z4X�x{=�ֹ/�ئו�q�Iy��V]�Յ+O�h0�Gĉ�r�̽a)f��ǰd^����uό�eF��6M���U�N+-�G�	�}ɉF�t���Rn�/~�3Fm��<��9�WK}�&^f��N�M"��W�{.?V��w�2����'�xg̛��?���?W��c���w�£����Bimn;sZ��)��$">ڀU�7cLB+��Ez��z� <�HZ�Lc��Q�}�i���7��w�	t,J4i'�-����Wo�t`���cQ�bC=1aw�S�!]v76��㚓󰭼�vN��1)<��%�pŔ-�18�I��㰤2�/�|�ӫ��@U�w��5.��	&�na����t���{���(�!�\�v�ty�Vzf=��S7��׮����Z#}k����ˉ�(=ƑDx�r�����h\��F��6��-�����D��^��K���p
�+'�]�����im�
C�A�����8�,�����03�!��:�'��;	b|��g�	�Ņ�76���/�����j<>	��LÖ��}Ϗ��>]t��Fى���v����p�q�Q�q0)�#����߄xbO�&����\I�\��������w:s��st�4~�����$,yx!�:<��T�kj4��V;�~�Pv����>YM�����]���L!c��W[�E�6�A���ID?��=�[lm����+���J���L2����y��:�l1��N��i:�=,f~a�Nߺ��)q#0*3�}^��"t]O�"h`�?݅��`WM��s�Js*���Iw�:<G�Q���+��x�&d��eg3֐<>���H��Q��$�%m$���XM��w}K�m?;޴������Ǉ�kD·�KHd- �1����7�1sTlČZ�g��"������u/m��qIX��U���W�ٜ�Z��>���v��4������O�$���b�J2����qմMH��\@��<64I�G0!��9%��ˊ��%��6��U�V�5]67)^7�N\��&�ӣX{h{4�� �LKEZB$~\��i�I_e��Юm��<���'�}���D,�=|/b����ӈ��نNE�.�H�!TO�}��N$��=k��YB�a=���d���Qx��]0�9�-($�FLm�G\���v��i�28�1�ˮ+�U[O���^k����!|a79+�^3��T�c�%�QC[�}���D�C����e)ki��5��Վhq����x	V�J#�愃Ұ�،$M9b�n1hu�L;�xD\;��e��[���-7?�=�7�&���=��v��4���$�1�XH�t-�P��=��1�c��bk�-��(Un"3X����͊Y�n?��/�E,�]žH$�D�_Hg����K����>h%K���|���~�լZ��0�{�H�k�b��J����-��7���G�Pm�-�3|�?{��D�ѳiu���\�k]Q��)�6��ǎ�y�=͛i�ڷ��a�q���e�׹��`�%�4��hR�	F�4u�d���VZYe$�q�������k��e����H侸ϴ�t��A[[��|t�9�>�lz��~��l8Z�N��~z�E�#YVN�7�Q�n�g�Y��rI�����4�>�@���H��Fq�덏6�ҬW�_㍍�z�,o���[p�m���]��L���+3���>,N=�O�[B>����B�kp���C�-�<h���Y��R-��~a�����*%;>?'���t���G�x�CJҢ,��e�v�<~�#�4�èO�-9�n��>4�ʄ̘NdDwI��]�6R�=#�A�^&��ѻp��
��r#{�~�`\������&���ⵏ�ɳ��kD�+��_��;&��G��_o|��g�3��7a;�-w_����t�>!	O|V��՘�L�s�H�ݤD>��?���ei^P�{���3�qҨ61;��%:h�uHV��V.�m&�.�j}y�ȧV	m{�J�2H6�/�0&��,H�~����D$�磬�#����_�=9|�u�8�&��`��=��[���[�H�M�;�㮧���^��Č|K2�������H\ߜU�V�V�� ��I�K�/�ۍOn��nZ�?���.��ß@�=�1d�67����CM6�~Q������))Ϋ�d|R˂�Ȏ���8�v"���QѨl������E�bw��� :R/���B�mt��΢ZO�M���.|��7�1�=�W%nU"����@��r�i���� ���u���8���t����ݣp�5����[c��b���hDnZ
�;���İ�H�G��!����d�I����Nq�ٍD3��/��vG�h�-,J;�I�~E4OYK>U9����h�$� ǭh"Ou��HL2���-N��D�SS����9.	�;K͸���x���8vF��L����8��l4�;��ttX��������o�1ի�
���ly�L�~�*n�)ckX����������Ʒ!/�,	�Rs��>�A��@?O�k<�ϊ�I�F�����zw03����/�Fb{E�Ds���B<�?���N�EWF���y4�L�C$1���6a
ьh�1�D�-L]Q��I)�ki�?M��bڗ��"��})g��V��b.yû�k�٣�RA��"�?:/.::GBͻv�!mXbhe�hE���&�M+$��(	�G?)��ъ�2��$(|�]RUӅ�<���nN�����#N]'awj��N9��]�h��R�M�ſ�*�i<�L:�ěWLƟ� }vw�J�7J~��a��A��_�1�p�t|���zun%F}�����YGtM+��b��8���Lk�J{_�3���{k�G�y���&A���ƣ�C��n�r�[�H�NY͚�����o�̢C�d�:4K��;+�te�J|��J� l&�;?V '5��>�>i�K�����eȈqH,�&6ʫ�
U�f�uF��]#1<�P|�����נ���^U�"��K��Eb�AbW���lN4w8G"z�����������M>�Z U�cy�Dc���Qi��7�r����X��j3��Y�(�e��B�y����a�݃�F�8>ZY��F��rx����[�T����U�nfp�FK;g��8�	���:<�N!�I�x�T|�&O�����dJZeP�^�SK&z$�7��b��ϟ�S���7㕯ʤ��i��<�3����K>H�Ӓ_c@Bj&�t�Rb�2�g�mu�0�L��A�~���7w�_~�����.a�oV��~�0���K�����ud�<C~ȍWO�d��6�v��M4���qu��#��&�Xz��r�#k������~��D����|����s�Y�R~��F;�/�DT<r�D|s��XQ0߭����Fr�$**
y�Sq�����tf]�+vr �v�^��z�liĵ'�£�(ji��x����6Z��S_���咝"y �F��4[B�;jxE�q	Ѵ�z��H�#Ls�}��ޕU�0�NYƎa�VM�r��;U�:�.<�NtZ��Jba����>Y�A�hcq���)�����DН4�E�\��:�9,��LOMbU��E�F}���sǛ[���Uy޸o ��f�����欣9�e���f�
V䰖�����~W���M��"�KGV�D���~]FF�~��|���d$�2gYlvD�E�%�|΋D9G��M_T�O��	Q��kCQ�"��{�I��y͍����yR�W�]M�o�nZ\�~}� ~�t��l��'"���9>#I�GE��rx�~��L��"��W�蕍�0w8���Rc�B"{����!���.���>#�}5�CݼJ�����F�3xՕ�UD�&x�y9��^�J_n���ە|��Y�{}+V�j2O����r3){��꫽�D=SC�k��^�O@Tr�������DQ���D���*$҅���)d�9]^��]9��.`�w\8�Z���z!4\}�XR���~C>Y^=��"#�$|}oY���#jg$�p��x��R��;�p�073��<�E�� �~��t��O�=��u�c(t�]l�f�L��:d_FCDa�������<v�$���6�J��K�LEe����y�x�ϓq��������8�aR����b�����X2��'����ILAU'N8(��[$�[C�����P.�y��]�2*W���K�؄�N��5'��#��ԋ��I�q���F�P�!a�[�����_�x�!^��q!YYٱ�ie�,Lc��7�v{�c�o�a��ft��1����Q��B�r"�ŬȲa�q6YTϐ��ΜqIX��Q�{�{E(#����:�@���3��sR"QN�i9W����+�9�r�Q�-�񝤑i>m\�(��?/�EG��������hv$є�Z�e+�j +��q0=@~�x�d#���1��.��Cǅ¯o�z,��&�U��Q+�LZ������4�MJ�D$y�\�y�ÿ�X����zl���?�;�Թ��8�@N3��rK	{��tAw��]�*"�p��g`8�sɓ�d�I���[��ъ|~��'�h�[��[�L��~+u�ۣ-��̄�漱I-R���F��\L����B�n�K�����W�(�s�i�6���:���d����U�O�F�d�1��Z���a����k|v�x��Fד��=���챸��Ѳ�ɟ������P�`��N���d���"���ٱ8�vWr��m/l�a��q�cpny��rzn�<Z$}�
����"��Y�E+�S?�?�'�8)�Đ�Ş��Ds]aK�X_�����\h;1�e���l"m�s��nY�t뮏�z>�;�Fa�4C(�V�0cLz�Hz�K"hB���u�T
�� ��^���s���+��,�V�h�O$����Go�!^�_H/0���.�7�CXO�Br�AV,��w+�]bT��q���A�[xC55Ut�;���K1ӌ<Ӑiyn�N�����ã�J4����Kv�=�Y\���W4�8<:Q<\ g��f��{]$��u��H7PR���h�MH�?A��HQ���ݒ�""ъ��[�/R�,�y'|Hb��86�a�NR�,�_�n�\[��w��/�>6>ZQ��â��$qQ��oze;��zҋ�$�D����Ƈz�|^�m�
��~1N��)��v�Xq_��ǅG�HH�������q̢�5%Qŧ�>���4d���(.8WJb��.LI�"�F�_�Y��6�KaW�����m!k��V��#�&t5�T=��D����8�px���9�3��>�hTk�+���0�f"�I��� ]�͍�V;t&.\�At��:��ir�ju�^ـD2x��~փ�Ifo5��p(�W�_��69��F����7��gfZ�x�^�N���w*��>��A�7�EҒ�0�y�	)�1#;-R
N���(����v''�XEM�ӿ*>�����!M���5*�B�F��6ʹ��m.��3�����]NCR\���z�����xT��)��4U�`o&�f����Ǣ3�u�����z�i�.�y�yo.K��#���������B8"g(-6W�j�kLȊK��I�~����tk��>�n���8\��
�a<�t���R%ʋ���q�)����;�a#��ri�h��F��M�d"�A��7g�:w�RΈ9��f)Ĵ��%%�)��s9��B���n��s�$�6�]��йp���,���Db Z��nk�3$��Ҡ/�����R���Ӝ���ѝ��J�4�{0%���}ހ���^�*�}�^�{��Ճ����3�A�c�����;K�1!'�''#->��\MD��N?xv��'C��lŖ���j�����G�#	��(�sK�|,×��3�7����+�:��3���U���-�U'\� ����c�BX�֑x��E�s��K7���(V�k�6��m�)Fp{��.6�9u�����;��8j�n_֭S8�'w��M!���|�q�o~�O5q2�~?�,�Tқ�=��"�C���As{�<z�q�/�����D<��ϓ��n��t�Z�G
&�����l����@��֐�9_�ɏ��}U�N���Q�/w����,�V+�x��2Q�l�|��^�#�y�`b�X@��P�쀱��ɊA%�]��6�Þ���i��ndK�+������������ǎ�tQ���U}���6b^͇	p�Z|�����9S��2G�(}Ģ\?���j<E��+�Mn�7F������s^�,�Μ?����_�<u�uY}1�7p��#�m�Qɀ8������$fp�=���&��M2��/�p��x�b8�q�T���XT�v9�&N��6����	�p�Q�X����b*�M�b�V�Fw�|4�����2M���"k]Q+n'��uȚ�V|���$��t�4|�EC�����Ȉ�яv�z0jp�^�t}~Fz�«�S�V��K���&	�9�J�摏�Sf2+ه��Ԩ.����A�&>�L�΀�5�;26.;g�Ÿ;n%��`�)2�O�ج��~U#:6�6bD��ܯ��%K���W��]S�FV�]]ʼ� ��CR�le9�JD���ŗ�Y���������)Lck���>��KN%�Y����{\3a�>\���H��u;I�8���݈�O���O��"�V�Gg3��-e�n�9#�Q߇��M�ӣx�/p/S�V4�)s�HF�E~�~�pX�Q+]ҫ��Ʊ.����S��|�sc���}�z��<���������ҍ]]V444��L!NWЈ�Xmm�D�FÄ�t�a�js�����C�3M� ���ͭp��;���:�{��?AS��o�� :��q`��M$���J9&�J��T{�D��x�7�f[��6�hI9�D�<6�����\S�7���b�%)Q�a��l�0���>��M����.u�gOˤ{N�����6�[n���b��x=R'�`߳�L�<��z�
!���F&��J�!+K��E�eļa5b��B~ʾ2���:���t�����HC�K�roU{"�d��m%������GВqF�Ʈ'��I�7�5f=���G̩���ht�N�)6yG�u�pvFI֔�z8����)V!-,������Z��sd���CxE2���b�[\�׉���p:�C�S��+0���?�uwǮ��G������!�l�N�ev71��U�6س�㇊<�����ᯨ�$`eK}�����X����I���ߐ3��!�Qt��A}i�]y��@�p ��bt�3�+F1���f:9��i���U�B��\b9�v��pY�ӆ�!�s=��B�����a��h/M�#��{�\�o��v\���_��í�D�N[��1y��8��l1�8��������))r
���*0>'5-v�Tw�Vn���hF�z���jAL�29ch
���K�����?�z���i�V��ɬ��,��8r�8�X�J�S�;B��l����9u�b��>$:�T��X2��,�����\���#1�v>�΋���h}QUGl*�<�i��|?2���H�.�� 5lA�>$���䜸�ד����:T���4�0{�w�U g�O�A�G뱩�%���C�r`�
���m�	�z�vh4Jĵ�łTM������+�v���^
��m'����N���7����.�qw�����1:�~�X|��<��n2>	���C~v6�7?�t��J臾:3�Jh�y�z?�i�Z� ~!ొ�b��Rri|�;����%W|��^�����ƒ*;#?mjDc��s�V̍���j�ٸ?��E���DKO���E���¢���-���Խ߆����l$�R�0'�
���l2C�eT�xjCis,��D귴�A�Cț>~D>+�(�;^PL\�w�x9Lĉ,���F(�ώ!	��爴(�vp�$��,�[I���P`4L�.��:0Z������(�?3RM���� f�d�d������2k`&q��[${w��c���	�řz��'%�*��e9��ȫ�l��#F�Y�`��J��A���7-�{B�_eu��� ��n$=�I�Q}j1$X�0�3�0v����t�$��,��!��:�Fڃ���������������;���\P�e���_�����W7]��ت'Z^�Cb:�		�+����t���t���53�n]�Շ�E�I=�;ZR�óÉ��q��T7�$��(�]0�GJ���KBݧ�J���f䆢6Yin�\t��֧�Ч����S.79��Y98��K��VZ�:��+���B`�݁��8�^5�Oǰ�t->{Kq��JLL�>H�4"�d?��h�3�Pb9�W �n��(��qc⧓~���W1�����7�6��+�<��%�!s3�8�vY�52��x-3�ipNZ_�!�.��""恇6-�a�Q�}�7H�\��LA���[$�22B+�T�����q���[K;���Iβ5����V^e�LdU����� �9��^�ֵ����!l����)�u�H�x��zD|b@vz�#�ZC~Q����`�����-M�k�a\v��
N�=�(FJ���	B��V��_��~�d%W�{�f�m��C�;��;Y��3��}�1�(Ǭ݌��&��@��s��K+DzP<\H�)z_�a��:5�$u��T/�x�2D��=�Z7�깈bY��an��_^�g{h=V�:�\v��)F_���=�}���։��ޢo1��W���TY�)��D��QN��/�r��^�wy�Z~�U��S�N�_=�s�tF��~1}L������<�!��>���j��*z���1�� ��WD���Γt�Gd�v�!��	0�42�Z�{h5����n��(�1��ɽ�.i�9���q�\#�q*w%��/z���f8me����ڨS ��42�p�a*3Ct��|����|HpA����|���6$�?8����uy�k�uñ1Vd�^޷;Zig��՝4�K&
$ޞ2�%m	R,]oK���T���^%/����ȫ���XYg����~�N�ᅣ�|��� )�ʇ�J��ܶ1���G(ǋ7UkU�_���#��x�⧬,��K�b�Y,�T
kuЛb`��I��k_�!����R��A��J=�����Y��cLHMI����Y��5�Ɉ�H��8��x�9����� ���W )sn���ElK��J�,�G�h�W/��?�����H1K�s��[���1a�مLʹYҋH#���؃k	4C���9J᜻G�W=áDC5J���T��V���*T*�M��E�r��ah��_~]�'<�t8��`0��f�3777W�j<v�v(A��餱�)"�CR�^�bi�8J=l@�\4���qz�E�L .�g{<35R�9-�0���ɩ��r<��vF/����斥�*%R�iI�V|w�W��lBx����S9�ƌ����'��iA�^���fB��88��B�fk���\
�S��ds#��-�>6��W4Y���S
���<:�U��^.���ڊFn��h<�a1�Z4�w:17V��IGLI0e@��������R�3��z3\�U��x%�\.a�Od11�)>Q6���x<�����5�6��$-6�9���CL��|�c�����s���fZh��u�h e+��5^=ocN�{Պb.��K>\3{l�����K*�9|�ty�1��"l�7���Y��zt83��k�T�[���/��U<�".g�z,X�@��H�@\j���j�!N<�n�S�! )�y�1�L^F��lr]�	���~ e7g� ۔�+v�����|��i�rƂKMz�@
��
������`�;J0E�w������=���Od1�"""�Y����=vbVDcu{�`ū�! )#�rJ����@k'1�O��Ȍ��p)Wf�3h�����SH\4����}�[���8D���޾ϭ?H��i�]$�P�:��o�
TD�c��
���˖�
'�b.�]'�]/�ʲ2��2$ eF�xW��]����.�z����ܚDO����isKu"�V��g�����C$_yW��i��B��Mˮ����(�9y�]�ht9����6��F�Q}v�w34)9��τ����]����1ljLF�H���K�}w�`�F�[�I��փif e�oiR��i��vu�.S�3�z�U��>
ƈ!\�{��-�C�\٪��2y�:G�_��/:$��C�t:�̙�h�y:o�H�Cb�U$��s�!hg�_��)�<?�{�D�uʓaR��Gb�z�
��$�'��z�Dw����1Դ�V�Y,)�f(���ƌ.++%�0�|��$UuG��B�z� �H R�k}���@����M7�S�E���U��k������ֈ�e31F�?�`�����@ʼB��땸F��N?�ӧ]9��V}��N�RLu�WD֔)S`0�0'�^-{�D�Zin��,�Á�:M e�Ka�c:X���e4;��Z�6�X��/aa7V�J��@5�Kf��S��<��B'��X e޾��n^�@��h��k�ڨ���/a�Z��)�56{W�Z)���	p���z�(	�8���ؗv�)+F��*��΄׈Q`ml�����f�.���䇴%z�`�E��)sn�y:��!��H��K�*������N�͸u�1{۝�B9�MEkK�{�	�v��DN�7Ҡ�$�k��N�Z[���G��? e�=�/>D@�.��؈= )3G�� 7%� �|~�����eYU���E����s[H�8æ?|�k�����N���8���x��{@��J%�F�s�a��6�)��R�=B*o>�@ ����̍�]2^�͍�����G��i�2q�KV��d�f���#�#\f/됥K�Kc�o��	/u�:18�Ds(@��<�y�!�p���~��^��{)c��!R&�$5E9ʫ)%5
GLN�wP��8���W����2���,�W	��g����{$�+�������Т1a~b+<:[w�D����L9��gJ@��\3�'$!�v�ڢVl,i��'�r�� )ˋ�3=Q&��3<un�T'��� '�Gh0���`��&���)�?��1��G�d(�!�g�Ett$��.�^�X[�N��J��|����{�#�\N�G�o?{�|v|:l@ʫj2%Tpؤ|��A�� 7=J�"�7�@/KQ�l�_3�V�#<�C.�ֶ�V�)졓��]:�׏��	���42h4J	P�BH��U8�H2�w'�x'���vPF�����f =ɀ5�-���̫e{y����)�K8y3z5j!kmgS����A���������:ٺe�#6��&���ʖ�U'! )3��l.��L雴S<'��ebIEK���i2����|[�G�y��J�����o8���:�!��OY\IB΁�s��\y
������N�N���	���� �}�T�p��	�)H�#��~�Hy[6#�/?�r`}k��j!�j3;��bI'���р��О����,	k�$''G_������ms[������\S+��{�W )��N���P	�g��������K�{�d���bf���Nj�Ɛ��7ʽ7BTɆ�@ʾ�=���ig��L���Qk1�R]K4̡3��Z;��n8u^	���zx}�k�8K:�,��7 �F[5;ތ�[��NÔ�!}�}�447����Ἴ���hh"&q��q5:�w�<��:�����O���ب_��_��$��Ay�JƐt��N�=���--�ˍW�:����.ή��!��Ӂ����&Y�������.�'��;^%wv?�N8c�'�!qJ���w�d_��8�$��S,�O4�W�.]̑��}g!��|fovVYBF$ŵ��w���آ��=��'�Ԯ�O���~R��^��#�R��B+���匟͝���Ix�#GiV6��ް��g̜	���Ǣ�N��x5���
���G�W/��;Jx�$�� ���tt�U_l){\q�H�
��]R�3��V�hg �1���+��BeŨ��=4M`�XT�;��'��m�*;�*b&��ĥ�;������G�D�"p�)�ʐCF��<���7�d˳�����eRT��s���o�Td?��F�)� ǃyp��F9�˯���x���#
����	��(jQ?��ŭ����	[�:),*�)a�\u���4��F'8�l�q�S�l��G���k�mR�ΟO���c��_��k2��2':=M�v�g��%�R~��d�)�lͫf�<e�D{;��*!4��Cs�9���O�j�Θ1FY'��y�`�[.<�e**|ǷKH(��1�����Uh�ZNL������ɍ�xǌЋ�����K���*e�5��u���z��L:���*oIH�r������1a�ҹqߩ��R���Rubu*c��HW,��F��	OP�^<A*�9�K42;p�����8�2���nl��H��,��
���w�V�뒉�pu]�U�$R��:�s�!�;��H�����]Z�	<E�n��Mlqh鯿���mQ�����[�����֠q0T��O��yVI�~�M��*�_��/����"��<�����2��ؚaq���t��i���6&�!��įY�� e��H��J���<���!�.�v��Z8��� .D�$q�1L4)�68������:q�[%�Q�j�dFg��G�I�-g���_���h4R> e-ցzSy�)��ʮ���F:$+�w�[E�̀vg|f�{�t46���?6�����?BD�A�Bcng�&z�p��yr�5��b��K��$kR�k!�h�;0㙮aR�K��﷩�:'g4��X��1�BgoF{}u�ҷܸo��)�Nm��(f�(VnH�[�^�T�L��/�o��� )E�����K_=�V�ٻ�����f��Y�|�d��^F��o� �u�$����^)�kcG���[.�=�;Z�Թ�$��丩غ}��|����\h�1��H|���]���ɸa��p0e ��5��J#e�GC$&2Uی�5���9(PC'C�K|~���3��	Ǳ�C�Z	�pPSW��J�H��8tB��Nf/# �ƻ�C'�a-_*N.�6��;�����KW�۶l��`Be�,)�cRn.v�Ue;T�R����t���e�^q8�%RB+���IcQo��l��Qzxw������%_�ǩ�{<�_�R�6�5 &!%ɤ?���Q5��!�:�/@���@�[��P���vW_�Z��Yt�A=�L
���3�v���B�e\��q�)��4��2�իk�am��6���j1/��.�T0���R���Il��!�
�,���\~ e�ϡD@�8i$~�؈Rr�F����2��_�C�I�6�v���Z�
���`=��%FR�.L�0#-ʺǗ�Tv����id�90'�EvdϦ���`�⃢�~���o%�,�����.�TZ���el*��3�p�Dux��"����ޣ�����i�lYC�������^��z�D�NqHeiu��0�����~�9���;�kw���a��t�0���o?k.{j��]���7��%U�3�
��U����7�%Ԝ���>+�m�縗ln�z�w� )5���A��#v�wA!3Ybz�3ǂ�S�;E����<���I�)	@��x]h�l�u�WH����9:A��-��FU߅Hy�����n��yE�SSL�K��rKa��^2�U�<u��0D��X?��q[���yG{�q	�5�t��b��䗼t��@�n��:O{´c�4JbWQ��ʋc�:i`H���yq2�<ìGE�z�Y�F �႕5���o){�B��˸��'&	�3��pdN��|B����SPP@�yL0f.1��+"X'\��9���7o1��Br6�b~������f����ժ<�_H��&<AR�����ߑ���+rD7�HY^9gp�;cۜ,>����R9I���WJ�ͅA5Nj9mx��G��ֻ�=Ҩ��ÎKF�ס��o��^/+��D^V4�����1��K/��RR���q�9��{?ř!)��wt:$���#�Ϛ����dyF��Xjу489t�xQ�J�� �H=�37Y&;�]�G�]tKk�W<�����%�!c���N�Ջ��'�%2| �<$ e5�l�+�v�)� �b�+E߻�>��|j��=��8sm�p��åú���S�$6.wkq�a[S�  p�B�O�kFM�؞;җ�#xW��,�{��@R��X�F�mґ�~�-o<��1��ە�S���5j�1��a�2<ڨU�R�1i�ZWW�8�0݋!s���H �=6"��f�7��{�����򸫋Ģ&Z�5wt ��;v�
���
��&q1n.�M|��ǋ^�H���6s@�w��H�W�j�(���h���d��{#<8ut1^)NGy�߅Օξ_�Ҍ����d�\;rd%`mFE��;���)�v���<X�ڰ��R�=Z�^�;�*�E��>�����Q�,�ĉ�dHz���Rik��s�F 6ѣ��,�1Cc�P+�v�)�1bA����7Cod5�"��}��ϥ�M�:w�H\y�u��O,m�啵�q����+�BT�p���� ���3�6�.���9��t� �|���}�4�D@iʫ&:��S�y�r��e�����s�Iߘ���
̕0C:�*���+�)��i��"N&YV�W�I������L�o	?��q���c��t�R�^_/?�.+��z~+l�V��ѳ�Ń]ˡ����D���h�z�_N�MG��a�W��%��k����a`G;���Z��G8����Ig'��̌A )s�����m~ e�7�6�5��:<������H�{˪q��H���1l�/��tO�p2kb���gZm P�z/�
���->��ފY���ݯ����9BR��1l=iv:���p%�e����H��͎)#���������d���j�$o���FK���warn��]���ܯ�fV���=� �ƿ��#��%��lת��}��ІbY� ����M չX��E�Q��ЄHY!/�7e2�	c����v�a�`�\�1g�`��>��i��|ԡ��_���M�L�孓��/R2�~���r�%4���E'D�1! )sq5;9$ϋS��u�/�2)ܛO-��K�4I��ω��	�q΂,,��"�FF4`�m~�_�'LN�T�ǡ��Q_�RԜ��o�.�k 1ѠV^��o�-D ��IdO$��YT���)�J4�ho���5��A��0Lʍ�c���
W{19Y���%E����V6�$a�|jQQ�7�{H��BR.k�y��x�������ާ��76���r�J-�d�w�y�2���p����x�)ʩ렢������0zd����ln2��[���_l4����m ��>@�CмJ}��i9������i��ځA9�S;`�����(�0/3
;ww '=
SG�a#�����w�	Φ8�;��!���8�Hy��|����1r,�����������m����;Zp�9cų��>��G�@���i���"B��m0�{5Y�;����ۚq��d4&������zx�q[]�*0���2ʣЅ	����]ON!Gw�V)t�bR^�x��5J��p%�Ұ�6{X�8�h�m����eg��S���-�y�h�I�i����"/�ٗ�= �2��>1?)� Gxu�Hy�p���\K4I����x�@�z#F8��I]�MJ/�@�ٯ��=�C�_o��qb��w�g;�� 	�����dÜiQx���{-�BR���o�Ac�QN�������ƃQ�(���!c�V3�|� ��&A<���SĨ)#�$��
1%�<��X2p�fބ$!㎋��/�$�����H���t_�B@��];YɑX�i	�ȋ7c�&+�@�Z�������g���2�nw�1a����Ԍ�Ȇ��0<�F#/�LizӒ�5�B~�#�S�[+Nn��y��*�+nC6����DS�-�5M\H�1{�r�qOxAJ��F'xc�R�ן�'ɘ�W��+&��_�p��t�{������������Q�i���I�I�/���wh|��ͮ�9�ɬU�L��J��RM)�KH�w/����I2��٫���#9�H���qɻn�N&'�Z�q]�Lx�Dp����8a�@�lQ򛝹���o?;�D�UD�r�G�Q��}�ǫ J0�$�ρ?��i�}D�k7����
�23�s_�ϑ4�z����Y��b=d|^_RIc
7�2�G�[���H�����<����O�K�M�o���TH@�f���������!G،�Iz���ʜ�>�N_$�ȏV�
�͉�c !�	�c1�|F��E�:��;W���KƑn;|J������S�w�|mZ;�������RO�q�O � �6(_�W�����ɠ[�'����c&���K��!��;9[���⪅#PT�):�K{�?e�T�/���i��Q�W��ig
�X��(���Eĉ%~c���}oЪv��Vv�R���r��4��c�)ʨ��J&%�ϟ�#qy�!��&)nf��K'�G� c��2L�o����5���5|��b&��s�9�-��e��1
*;�[��n�cM�9����k,n���y�g"���*��h��4Q���+g�]�d��}��^��/L����wm$�UDʝ_���v3�2]�m��/�󼖌���y�qڡ���R�S#B2Z���̘�|�æ��]D-��R�`��M_��Y��ZI^���k����t��v3+.ʀs˖�ُ`H�+�@qu�|��dT8�
] �=4�?r����ݔ�j�~V�j�F������&��)}�� ;��.��SbW��>!'���k,�d�^�^U+�*h�)�pE��2�rM�t{80*�)�����'��,���*ӫp�.���fXm J�T��A����b��R�	 ���>O��cwc<�G.���㒱��LVQJ�a�(���QQ���cgf��G�hj�M�َ��Fk㾃�{����s|K7�@�^rM�z�F��luF:`ej#y�GK���}��L���K��z����tM#��"���܈�1D�)��8�����c�p�q�r�t�[|�%�ci޾��P���O��o;|����rU�8Yg��C������g���1�S���G�E��$��:9D̸�|�;��K�܈��e���2d�8D{��'�b�dĶ�af�u���7����C�ʵӑ��)�]-"3R�h/��k�Sg����WԅH����bkeMa���l�o,i�c�a��,\qB.9[�8��,��[x%/��s�����S�]���q��:�֏]B=�"�E���x�h����GJ���-�7���>>��<T����5���G�`\N�$�؊{��d�ՆH��������������Z-��^����'�NG=���g��w�^N��ˡ��̕Sp��[c^�Ec�dB�h�ѿŴ�7��7���w�Ǔ$u͠��@���ǩ���gEK���k��fT�Y<��L@�op����������/��@�:�)���/�Dv~����<!'f��v�E|��6}K���s�aݮNlڴWM���
M�h��.�^�j��x�9�:M~e�����}����3�Ecj����W�>/}���fB R���<�wf��y�W�A:Cx��n�讧iK��B�� �g�n�+����t����<�`7�h�:/�=�
'�(�Q�N$f�D���QJ�y�}�����݊��.1գ��Ȫ�"�,�g���m�[��;3��:��.	t܂����y�d��d�|X�E#%�V e)p�{%�Þ-�ǫh�������S+xYn�t�g���Y��*tC����ŉ��B��b�eQ�O]��ۅ��W��D�c���/��������<�aј�Ȅ�?2������ ��z���&�w�6����U%RH@�$�""����Jښ#[t�R��Jr�y�Ҫ���_M����cU퍩y��	����b�K�5��k�p���O��ٿ��8�y쯴�8g�y�V�|��ZF}�1	aH 3F�lg���8��a�l�ObJ�@��9�>:(���,�{�G�M��2C����m�.�F&M@5m�4��lp4���Ok�Bj���]��z��3��*�T��w0���#˗N��gc���(�%��}��bR��s�����oSs*,�]63�|%�D�6�>��_�����.��mFz������j�O�[��-�!�� ��gJ;U[���>C�~8`��jr�䠁d<S'b %n�b�h�3~~����ҧ��5��3�X�^=��$5}��~���i�� )��$DF�a)1��6��E��`#iLu�>|n���~��{X_��гL�̸O~�/���lb><éke^����= ����@�5Z���?hl�Z�����G��=�ƴ*������[oy�������u(k�cz:_㉗w$��scI�2Q�p9�$֢�����Hy�ƀ�5�Oǎ���\t���Ė�Η���BQkb1�$|�F�|�A�>��M�7� ��0�l�K���vZ���c���Ayp�^ӿ�Ą�5��1x��aR&ϭ{�i3WrPg�WV������W�h&�b��s'a���8at+������䬶�9�_+� 7�B1��ބ(��u"6?��*3p��I��>W�l���Y�{$�ćR�@�p�\�����-'l9t�ъZl-nł�i8��{��}�JԒSȱ�	91���"v�z�M��}��٫����1�}	2b����!/��4�Ռ6���7���N�\��y��T���Fئ��zv���D�74 ���t��r��)���=)�t\T���{�)�2�_O��g��$z��<j��:�l���*��ܧ���.��c��ѽ���5���/�8���U��G[p٤H0��"�j�x�[]z>2�5�]"� Fѵ�4��H��Tz�Y8O�x(�F�S���B R�Y��H����t�b�&��rg�@���	H�����z�G�*����3R�ӦF46X�
�IF?���0��^�꾌�E�mĪG�ݗ/�/�pF�&J�2UOR�5�����%
�N�=���$=�ݴ����Z@�'��s����pܡä������,��:�Ӯ~~����~�X�*h\C����MN�O����V������V;��m%��{.^��T\�lY@�b�Ef���f��u�5���*����msa2xp��}�m�l  e���ѱ��~�W�x�î�)����ٚ�=8��(�]0�GJ����~ZS��2�G0C&`5��y7-��w�I�{�]Rsy9�-��+���e�ٕ���\�uZ>Κ����UI
��ӹ�Y���Y4sU��珓(�q3����F�D4�. �fK41݃{��\P� ��?^ۉ���\�񱸨�A����K0�����iq�G~��ߕ�o��߼y>�փQRkQ=(�xTF��X��	��sVmiR�����$ e>\�i��_�.@;cGj�B�0)C
Ֆ��PzP�ǹ@�Vޚ�V����:$g}���5㴭��H�Ĭ�	�ĥ��
�Z�ܗXGV[y2���9$4 �2͙_Gۤ�P4����G��/��J���|b��V�X^�/[���"��:���Ղ�^���Rދ���#��w-T ���S�0P9��    IEND�B`�PK   t~�X\��䓝 Wt /   images/4809d2c9-d031-4e44-9b5c-1a8b0048f1c9.png�	4�k?��)�RB�SȔ�M��(B��"2g��ls�Hl�D�L;��"2�����d�f��:u�����}k}��ֱN�y�羯�w���~��sAI~�=�0�ֳgdT1��Y�N���O���j�~�;u�����*�{��-;���gͻ���w��jګY����cp8�uKs;�+���V���d�=�~�Y��#F�ͭ۩n��J�5ǆ]��_*^-	�w�s���b�_����v���O�oԽjV�kw&X�]g���_}��z�X�C��Cї�J��EBxU~?X�<q��8�][�����[Zvۿ��C:P�}`_���)�V�,i�)G몁�{k1Зs�-�9oo����׌�i'؅c���u�_���rO�������9�n�ž�#������HbgO��l4��7���N�/R�
�PSHJ�M�+j�g=Q}�O0���+�j��nvl� ���4�3E�w��|`K*�t/f�ש�P��n��p]C+{�QY`:o�|�'|�݉��	z�g�����vL�ݮ2�	�$��86ױ7�x���-mk��\���9��晭��`�~^Uj<K�7�?�Rw�8!��f����s�v��U��E]��,�Ε�m��O��]�7���:b��c)x<�L�Ѝ^083ٔW���;v�<]<RUL��8#\����IY��+o7����촷�!Nf�O�Ń���2U�7Y�9����?�O祣��R]�G�ǎX�6�\�O������BA:/U���1?�z��^D��ޛ���������\�A�:X�����e�}y2����}ǩ;�n���:ś���|��j
��.T5�Xv�@~y!l���z5��8.� �� cdC�q��m����F�3��F|p��(�tm�~� ?�(����A0>�^�<C��Q:�R��j�P�iN7W�����9}�n��8w,[ ��s�Uˎ����b'c�����l������s�8�>e����<�=��\Y��N������/���ԥ��j�ɚ����V5�螟�qF:&��t=;�3�%>_ �S�Ҝ��!;�6Mn��%3�;�=D+/ک��d�G��Ar2��v7��gځ��n�J����O혳h���4��&�ڲ�i��^�gj��z-��G��Kh����RH���ak硲9��
z9wM�Aj'��A��v"o�_�-�
1�m�}�����<Š���!$H��X��^���1�ZJ��T�I�m;��x6�~�c�5�����)QI:k?XS��RK�#��	Zu�0չjY�u�!*�Bn0v,\�1�5^����	)K2
Cx<�-�p�c��ˉ�	�4*Y1��E�e=���;U��`�h(��+c�f7�LI�{qB�ez_%l�²��"k��ǋ$̦Bٻ8��pt�P���M�#��Y�"w��1xYYr���� Hs��\Z���X�< Lu\pY� ,F�$�����Ǻ���<*���(�ZMUAY�hZ^��vB״�*lާ�����Mv�]��* w4�I��*�H�RG[�L�:��Y�QmY�J�s���gy��e���A3= @� �ϑ�#I���� 6�����S2)�i�8�ɧ챓��������y�^$���v#1u�vf�3w��(٢�l��,Y{�I�G�~���+���_��&5e��H���p `��k�k���E��v���H�V �~9`���Saq�?�q�l�2�总�>K�Aj��j�֭����d��M��u� �:2�:)��q/��H��	 	l *��?^���uލ�ݽ�:r�,�W�w�t$o��^�ޖւ��B.�#����<�V��zd��Mr!���M�H���wl�5�p��3:�k��-���W��M���룔-T*u�AfA#[ǳuz*��G6pw� "��j.�R��L�$6z�XyFuܱ�pg'w���:6�x��̾M=�����c[�7�r�\��S�,rW�Q1�A���K'Ɍ�\�l)�v٧ᵜ	(��s_p4��$�/iC��X��ZH�^m�{�QCt	�Oի���NS <�eb���ʸB�V�!Z�8!sp�6&<4$��BH_A_br4��������I��i�
�;���8��͈�ğ%ƾA�J
[�z�j$�7B��7�_�"Mf��nkӭ����ddd��4���ݝ���L9ONM�lٲE|��R�=<<,�R[�1���o�+,���������m~����\�v��CV���Q���"���6�<"�����!NΞ�G<�Ǐ�jL1��ٚ=��������E[��������������1 Y����+ Gz�E�<��;PE�)��ƙ��H�5��=z�С��b?�'vk��>>0���]�>`/��k��X�?I'S��]Ix/�_����h�꣌bL��e$�\�x��@�k$�q�s���v>�4!'^���n���F��@US���Eg�p�W�fA����go6�H�J� �9jq�4��fWm�� �k,aNԶ!�e������y�`���Z�$�%ͼ19���bt��3Uԡ1hРq@����Ψ�)�d�  ^���Al�Ν;k-3�8o>V�hN?H.�'gQ
�Eqs.��i��Ғ�p�jG�X��N�g���8U��\#	���KJz����9��;�#���@�E�TiY����U^�i8
y>�i�$/�����0���� I�PyzUM��	<��Fm�E���e��i;�S��cRl�bσ�Q�������8���6�|2*���ZQ�n�`�0l�����	,I��=y�M��3._�R�Ԍ=�g�^t9PXI������*�IYj�>��Ǖ�;M�;vݢ�Χ��<����`bbR]"�4�����c�)����)�ec���/�w<�%I���ݽ�dJq>�#��ґ�<�F���b���}'҉\�F�i|8Ŕ0!�C>�ȮZ��X������V������f(Ɏ��i�p\���ܭ��X���3�$g�BlF��D�.�jm;������H	�)
�W��DŇ��T�V�W�!	�F {7��t��6��f�8�-,�FHyH�6�\A$9�TL�u�ac� ����Di;=��Z!R�rc4 �G:v�\#jg�e�㎝	��6�<<.&������D�$y���#�/�)1�Z��f��J�$9o��t��h ��ǌ�sFFF��s�k3�\�@ �� #�$��jdO�#""LQ�=� ��b�g��ʹH2���>�TU�ep�J�� QwY�8�U���g����˙�R3���?�"3����X,Բ-�DH����	QQ�a+�-D�����A����qN����Xl8�k�'��E�9Ոv���3�m�D/�� ,xq���a�
�ny;�}Fss�L�ԒQ�4+������P�	܍��ϴv��b���}�I�xgr�%1+�R����nSBb�e	S��W�m�989Du�C�V�aB*v����[)�}<6�-Ķ݉�cccg>�0(**f��4��I���,͉�O� t�vѳ��J*X�J)���ik��>Y/�1HbZ��o)�*5u�j%Z)5C�����ȃr��z~)�S	�B���[A� P��2[=�h~܏������F�̍ёX��5#ښޫ5
��w�n0#F�|� ́��{�T��d`�eU� ~>��L��P�b�gڙ�kn_^���7ؔ���X~�Ƈ�\���T��-sVf��!W�:(ks>����q�d����¨ց�6[�fT�$17�j��W�;?=�+p�����g�n03���J4@�G�����v��� q>D������h}=:���,��;D���U��d �L��m�=F�ə�/�>����~x��3磹���[�NQڲ'�Y�&kIa�a1���*1��k�T���Q����6��=�,;J�E�N=~ <r��s�{|8#g� f�����!@R*�ut��/{��|�ȶS���g�<9�$#3��\���;5wy��K��~�B��Bv��x�N�����.O��&k��SV�zJ3[�u�j�=���Z]�,�ϫX�^a��<�:����v�I��Q=�Qu2_�b ���g�v��ܩF�\�fPɫ��F����'��ë����gff(�ε�E�l�"�`;�5�����&ȁ�� ��[�	t�9a�繓l�S^6XX8��X�W.miI7.ϴjϙ*�='~4����+ęS:F4��ɿ�ʽ0�㢢����;�O_$���I�ւGORKlrE�1����W���<˰WĲ�P{�rJVX絅S'�tA��	$d�ѐ�dAJ��8��I#I]�#n �n-�	�����$YC�L�\�~����e�8�u�#��ܟs�z����yd�'$�R���bm9k��*�E�.�i'���Ea[=�Y�
Q*��\�m����X��rFm�ER�:ݨ}J�
��B\����N������]J0�dF@^Z��<�ӵc��__�~Q����X�B�`cx�2�^<��	d!i���PNM����sʀ��^�l�)�.
K����x�%B9�i���@���D�Dzm\R�O���ag�e�>@CߩOCM�M�g����)����3y��m������G�{����s����0�4����h�
���G$%�
��T����ܜ���O:����Ú
ܒ���N�/
'���r��V����1��C1O�+� ��&v=	�{'M޺eKխ�:;��F'1ya�-[���&����ß��'�K�:q�s/]f�D�X��S�v�s~�\vr�|;%p�B�­7� ���m�O,���"�s�ԛ7o	�������+���4d�ڨ555fm�9�c��J�G��֯_�M��E�:^�vtϾ}����A��`7#�TF@Q��S����y���=�ss챗��o>�Nz�$�C'Ӳ����0�Ķ��-����m�z7._��@v)�#9�<kЪA<�B�Q �s">˅H&��L��e/q�؞�R�����p��T���$� 9����u�@�d��(2�5/Bsꌱ�:{�����4G'��ƹ�)]���)5{6n2œ8��"�m9Cj>�Jgj3��DvT�Z<��	n�'�l�[X�ȑ#ۣ���#]�o7�޻�O�c���(�S�|WWן ����ҖM��J�UEؐ����tۥ��l����0?������nU��r���A��,����F�\�u���Q?<��-q��ݻw?�j˪@Y��;���:sۓ��C��$��V�'���}O�h)����Y]���qJ~6o�����=)�Ao��,7�z3���2 A���[�:��Z�p��H�TEIy$��;U:�0	����d&n3��ff����
Od{&�2���98��`3s�J��K�y��U�.�H��͈�1���v�5:�����`�T�չ����mqP�ggԌ̖m� ׉o0�5Nr��gzק�����i<^;)��q�-l_�"��fc�8�N��M���)Ԑ�����gTK���(U�	n�aq��ԟ)U��.�����`������4�Q���aWb��+�J-x|ُJ:d��*`��kwp򕗗��m����Ec��<�iJ'���Q���'�Gӝ�l�+¢�I�V��Y�(��0��-W�g�fc_����Mg9�@����1���E�������i��6 .�����tcE����W!:���(��B�D@������k�=�w����#P�rM8yU�3.�|(b�YX*	u�)X��qC���>̯�s,G��FI�:��Dȉ��Q�ns:�=�:Y�l�O^�ڎ�����^���jh�w��A++�P�kj.�#nB��y;S^���d�"��D�x�GJ�I:Y��IU�>��`v\تc�ÇUB���)�=�����ŋ݀u���,P�(�d�$���\�/���1K��l-E �q� � ��l/�R�q�"���!��Z�>.�NP�v�j�����T�������SM mGZ�<P��8���S���l���M������FID8:5��p�2.Xlx��*�a��M��O��
�V�[� ���PԱ1�c��p �$��q&��q��&��h!���=���3�>dP������P#ܔ�0���Es��S���y' �I�\���.)�c224d��`-		G�}��Ճ"m7�a>\�f�cg	�bb-i�^|R�_-W$��3���Z:�ej�CV���Q1\��o4Wt�E��v��@��%��?�4�T��ͪN��-$$�cU]X(����I�� �������;�߁�Ѫ/{����og�E�=	�{z*�"y�`Uh�G<�66��mV [�9o\�b�>|x����aaZ��Qb��h�����@�F�+q3�E���lA���l����,�*�DG�bo��h���nŽ����J@U�>r�B�w����,�M=������7ɘ͡211]��]����Χ�%�Ǩ�L}����'j�|�II L����(���[��C������{{��zP��)��v����ph]��t?������e�� 	//o�ҁ� !�|����q�N&�?y�j �4�9��9h��a51솢�¤3�ŠY[�m�]?|�g�柵׊B�tr��X�U����h*��`��3�{q^P��R�k���Z�z�p�l��y���Z��r��pe�3,�����NV��)UT@C{�W	�R)cmED�O���Y=7撮�ˠ�A��K��j��e޽��6n�7h����	#�'��4Fv,i�4zm��&�j-�n�˩�,�Ï�B��\��ʌ����?{�������N@�px�ʝ1!�>}���=_������=�Ү��۶�'�����)���p�\'��I�P�	k��8�:5���E�ha!o�_F��{ �P����g�Z!�=E����l������\
�]�KӁ��������oߞ"���x����LLm)!�ϐ����}dT.t�c���:�� Z���M�n�v-~@�銥%?99�4O�����~ļ���(��)̈S����N{���hǉ8���� \T���/N�^��y�_�����nC��N�[�1��JК��J�� �w6_?�O�LF�?PO.����'��V��8%F��9>�1�Ɋ�B�pc�<(Z�rnٺ���ֽ��I�J^𖃠*#����C�ub�j/�������e�(����G%$X��yp��L�����f�Cx�8<��ӓG,�M��y��e/Ī�ܿĿ�dm{K��7@M�ww����p2{'y>���#���=d���Y j>�\��'���Ă�K��Ǐ�It�MT�i� �>�A`�i��[.��;� ��$���X8l�d#��SVUAPT�����iYY� 0-5�r�BuB� x8�j�n �QX$C���K o ٴ��+*+��f�Z��`I�����׎��?`����W��MR��+�~l̚�趶��!3���Y�] ;�N��ʼb$?��Ag�����Г��l��?�z�T_�F}�Oi��'�'�Ų�Qg��� F�}$���4;�d�SP���" �����Sw@z(F�O�<[�!qMH2@]�����0��ʣ�K�x8p��h�3��k�,}�rT*A��Y���w�\�_or����xb�J�B�� ��J?���k���Y����lL-Xt��FTpD�&׀tz�& ��'UQ�qh;�	h�JJ�@,YP<���s�ű��e�rvs��,Ǚ��T�����)x������}������������=���rg����3����G�3����;��D
b�U��	 ]!=�JH��7�������X3D� ��~8s7�cqH��J��!��`���a?�-$(#S���Ufk��F��ƭ-�S9']���i@\
@��I���9�)�f� ��-�B�)�.�� +�h'�|�ce��.�4�Z�=o��u)�!Z=�����kI��tx`Gyz�f�$�9�q��O��烍w����'<�"g��(t�~��bB`�K�Z!�f�eW+�6�,1f�H��c����l�\@�*�>���R�Н
$���T��J<�}�:�>M��##SV��a2�#�Y/%c�M���JW)6�b�t����=�^-���%D�"�»<@�j��}F!6]\�4�P�d�5�l@bdd�3�7�O<�r�HPsIU���"35��l><ߣǎ]���3+�Ft����H`%ϣ����Դ��[�c��r�m���PPa��S.���v��%t$]�#��[�faf0jm4.����x�A��̌����cj>WE��)@Z�]�b�r��1�j	�.z����+Ϡ#Ц4#�a�۵[�5s�ym���7+��V3�<PdT�;6�0���NP6�F�2�,���� g8ņښ�?��"2�r�ږjd�s��ʊr �#�� q�\#�\;����� �+�k5�h�`�f��B�'i�v+7L�]��P}gn�H����}�e�xG:����i����?f��`N���X�^sy@AP��d���*����0(�>1�A阮Q�د[��.��q���TP��H�gE*�A��@h�ĽF��{��2�'6T���]sV��*��~��H�0����NZ�;������U����2M����ΫW� ���p��.E�i5B+ְ]%4��T_i'�!�b��]7 (0���\>� �󮬟i�W��qi=g�E�^�q�F���( �!h�Y���$�\��O#E�*�̰>R�[74�@����r�Yf+|�~��E�C �֤��yތk�xߜa�*rګW�XxWO���?��Z�m���2�z!�;�ǀ��qD�$Q�%W�p��F5c\Y?��[�d�������YQwKWk��������Ⱥ�$w	���Yf�LV���gavR�m;�[>��"�'�ycw[���� =D�[x
Wn�ViH��y�Z�<��h^Y���/;4���V�R��E��I� @�>d�~9`坹�t^v�����::@����l�㡆�=Nx�{�V���r�Y��/5����-2j{�7h��=���x<����ͥ/� �,��m���	�M�����W�3�o]+�S�����m�Ė�I�I&�ϙ�m�D<�y�5�����(IO�����@ 'u
��r�	�+x����A8Y7{�P���~�=��+�3�B~ et#xǩ;T��qǔ���e�MPCt�|1p��"0��HS�ф�z�[U~���D̢�_���.?�l@*7���|��[1䩄�h��88QQ[�n���y�|*�c��XYEq��nP�	�|��w���9x�1Q
���H}�Q	���k��/--� 'N](x3�x'@>��UTTMN�C�"..�{��fl9��*ׇC#��vniYm��l��8y��zfz�)߇?�2��;A9�I����Lgq֞�E����-�/)u�BCC��9o���I�z��n�Kݞ�_�|�|
�?�7$�]�Az̺.]YX�X�<_'6�F�L ����<~q�B8���Ig�,�-`$ɨ�ŉ��iQJqq����@�؎��)Gq�����Ԗ���t^��րw��8�7Q��6��>MY��W�d$�[�8䦵[66��>w�ꞯ_�3�Zn�[~�߉����ǝ�:*L��?p���-��O�s����d�ۈl^�	�ݔF��	)�1��q7�*T�LdR\�B�wg����ygɊ�>HډH]�v��q�����N)@��b>�VM��y��F�q-��@͌|����UϠ&C���G1�����w�7�w�7�w�7�w�7�w�7�w�7�w�7�w�7�mÏ���+���_��/o葆�ʵ�o~F��|�ESV�V:o�XsH�=�t���B9�=�����6lHz�v�'�D����{~���)����=�v��RG��e��î�:{�]��f-�0��%;�����e��3%|�*��6K������"֦�A���A�+����f�g���҂mn����*)�`3|QPSW7�aq���B۲��͛�ʒ�k��y�-��L��v-jc0Vִ��Z���)uCA�	S�^��%�kfff���i���/߸r�GP@�bu]��]m�F̘��,	���-..�222.u*���,Y���^rñ����@���?._��[�YXl�{'���;�ܪa����*����H�pC���k������u�p��`���-~�V�,�I,v�oWHn�pȀ+4�"]����� �q}A���ۅ���i=��I����c��sh<�A�:�\����+k����=� �Hc��?Jv�����*����yt��n��
���ޖ�?lC	-�Ǯ	����v!(x؋��θ��(��R���:��NP��'~��!�`-&��L�$h��ӋU�;X�쾵���3g�A(��8va�)����N�/�@�O�%j ���2�޽�Qq�QK��1E���1���)��驩�SH�s}��2E��񟹛�j0S$H�x�Cg�V�����#R��d�z��d���L;�M����ۺ`���跉m�R9<�e��^�-ߡ�:i�4�?��4W��|5�A*�˸��K�?���rER��ݱ~c�*QUJ8S���ERػ�}��U���ޖ�G�M瘯�|�ʍ��y2��y�E��LV���#�����:u��I��ډ�i�s����EDJy���Y�QuC!�g�Wֽx=:�\�*�i��0I_�#	����V���o���5>_�81��p��4�!?�S��c9X��u�٦�������ee���l�2a��gN�="�i�Y�mF��ڪlV�b��}C|�;�9�A����J����zV�/A�/LM���&$�i.`�����]d}��%�k_tH� S�o�ݧ6�����eF�U��0�t��t�Mf�uq����l}rfh
v
.\w06C�~by����D����v!��.���ɭ���t��o�i��N�<r�R�d�6$"E?�ABfTf��ej��͸%H������KVD���<�)g@��lw֞�C��_������fi�0c��4s�)x1g�;��o|�O���ĝDov����F��]�Ѓ��>��Q`ő�lwמ�EWT����g�Z�����u��'{��y	���U�]=�؉�I��=�Hi�*=�I`�
4��]�=!��Hr���.Խ�5��5;����#-��� ����.��|K��\�dD�[�Ǝ��U���pڢ��0~n!]|9������}��D� bM$�]�G���=�=�^3�ۉ%��+�'sǻ-O��-6��߉�{8�b�h�9M��]���EȈ��D����ח���WO�hz_��-@�?�>5 �/���-7ڞ�R��A%����y��o�7�	��3��7[�}��^?|�e���H� �|��Yki'��E�_q�,��>L��Vi��AL��0k���y��h��?���|����0�Bj���Ō�Y����k�:�Өb���t�+6���aRR��h�G\��%���"=���;����ͪ?��޼yiO�݊��Ҋ�-��E�g6���f��C������փ�c�!z�d��5���bXc������׈Ý��	��M�F��d��gZ�)� �D����Gz���5��]w�A_���e�����b|�!$�n��Gi���U������Ⱦʚ|���n\�`?5�m�Y?�f-}��ҫ\S����]�(���[¿4�����ٴ�8�0!ˏ����CBC�/�V���-�@��_��Q��';��d��^N���$c�IM����AC/������Z�n����h�
�`�v}�|��zV�0�1Ӌ��O2�"X�/�o�j})X�=E�
�R�4Z�v �ێ t���[���������@�^xL����6�з!r=�� ��I���`?"��R~�،�@��yet��� 3WA��X��7��4���8�yZ!G��W'N{�ox��ߒ�#4
���l*.M瘪���E9�0�y�S{/,l�K�PU��>q�g7b�B뿒�K���Z,Ɠ�o�CƢ�v8����"�%^;��\HA���NV��8�E���U8�$la�^EP������Ѿa%$g����F�K��&4<��3���{I�`�����x�e{�
^>�-PN��nf� �E�����f������Bl�kKِ���Y�i03P���@+w�-ETr;�����C����"�}Z\(�'�S�*���|=�8���8��1�S0O-`#hm�C�h���2�=����<d�B ?@��˒��!Q����ьO����_��N"�3�xF��N@����]�8#J�!Ǽ��a��&u�M���&�a�,�ؽ���8����+���g�x(��� Z;��m_��ɰ�E�s���T�>�u��F��.�����z~ ��L��3#d7��������/XA$��?�lTc$s\t�B��뇂�
�����l@���މ��h6�l�H���,e_� �Hl���A�z�*.!�|<<<��
X�q�3�0<��^�%qY�u>�Ve�~ڪ$�Wۉ���z�w���-�MuD���pɏv`Yu;��x	E8k��)���?��N��X���'��m�-�ۉ0�4gUq<���	r�����3Uq��F1���� c ��X� ���ԵkSa �����;;����ݳ�0k��Sؾc�´c����V���D�����xy�N^�Ի�EZ��;㌔%O)�	��N7Y���oO�U����\G���߈Y��%�	�v�*lEl�?�GE><وa�H�����W��~R��R�3��B�z���$7����
�������9$$1�9CO��J9��k]� �~v{�b�4��f~�{x]��T�(�f�&z�����Ca��h�S����Ok�7F�Q���>'�a��������WT�e���2r;�b!08މ�æ�p�̨h�����V�x�O�ڦD�Q���׉��e--O �!E�B��h-72Q��w��/�Ϯ=�� �sV�y� �e��ˌ����ՙ�ӛzC)AW���I��Y�O�L������Y��.'���3}�YP�?�Z�ztz�-�S�ML6��h�_�n�c���c
�(��iw��%)����?�*6]�t�h2wЎ�f@�����=Ok=�@��9�ݿ�?��X0���I�'@?2����Մ�b2\�l���'���O�O*4Ґ̚���j 8�z����;C:�5\�+S^E;`� c�����#���]��=�v��5|�#�(���m(W�@x�0�R��1��5�݃/�Ճ,�֞�p��$>�as�#���7�%�a�n��^���/#	'M�ȯ�t�C;����͠
V���^ج��E����<���b�6L!݊�~�˵2W�����6H��gP�@&�M9-^T��F}�
]�	.@Nd��}Z��%��܄���Z��ap�@��)C!���1�q��YSQ��*��[��?�mï�����5'��(A�i�VYPq����0�xƷ]i��WǺ'�#���E%���S5u�G؊��k ��l꿭�_�����?�%t��Ŀ�s�Z��a����������I�r�e�X+x F��z?-���}���wԕ�cl�p/6����,�	�!��8�l;Q'�h��Qv�j���Uh����2��<�M���v&��	�;s ߒQO��X��j#7���]��U����0��wOm�4=�����`i���Y֟ T}�F�/����&�� b"�8Ү�7��X'����?�;*�0F����$����b�M����^���i�$u?@�+hs
���M���0䈍Ϗ?�	3F�[�rG}�����f�<o�iVmb�����THV�Wc�9��I�+�@�MB��&*r�aRqd��3�{�H���^$0r^~�p V*7k� 	�or\ʄ��O���?es{�6���e~������Ʒ��G��Nn��뿭�=N���n�\���?�٤4e�9�\c^p�4��y�8Ū��%c����Kg��ˋ��-��;�����Bl�O�+��E�?�(�O����7�����@�|����\���`���t�k�"��B�pƟ��iB�b`������b���wi�ؒ�=���ڵt�dt�=a�b,m�ձ���6� }��t�Q- �������~���y�ٲ�t�X�
�w����ٳU�� Ԍx�ڞ�Ϧ21�����_����+`S}��*���0y����ʀ�̝�B�1T�C�H+�<(�ߝ宸9z~jd��:\�tB��c3�"���#��9&HaY��:�,37�ߺ���;v��=	�;��J�F��Q�H��V
�8�@{NA�G�J��"U�]eF��� �?^��Y�� ���E�>����˔Y�B���������6=qP� ��]6e�Ώ���T}d�݅Q�/S9�IIg���i޻W�[��0�yi��^[�سe�����e�d 8���b��>��%�nZȁ:�6  1�v�,}"��s=�hž��J5rNt��Kq� ��\!��?����� dd�I�O�ā#�ոVW�݌��6}{Ȑ�$�e��&C�d��kDm�Rȝ���ϊ�
�������QUvU��j���9�
T�;f��Z.���nnn��6櫒[䴑@��^�Ƹ �4pgn�
�*�J`>ӟ�Js�2���8 �)��1��ᰧ�"ȶ��R9��d+�@m���&�����	
\hLq/�ٓ���������jO��P?u�T�SHE���0���g�LH��[�n��sQ��ޮ�l�u֪`(��gn [�Vо�Bp����DdJ4t�1�煫�2��L�3��pUm{��.2��H�2�X��M���c�<�'1����Z�'cPu8=0���ь�Ʒw�w��L�����	D0W���!�&��ڙ$u�V�+���N  U��z8�[�tm�H��H����'�ƨ%�x5��؄���w��F�B��X�m'�B(&>^��*���P���7����J����������m'��[?���^�D(��t@z_mq*B-�YW��,`����5f�@Z�G
SFRؐ@/!8�ʭ{���Gn�WK[��fڛ,$$w �菲1�cD�����������5U�^�O��3�/D������UоO��P����iW-��	��g-`��d�;�NgR;91��,D�7��@hѤR	��(_�籽ծ�����՝+�౐����[:��#<9���0��=��G|�?p<���A0���v�}e�����|�h�D\=�8�E:tv��i;��7��'s6dp�;��1M@݌a�c���\�y���L$ᔦ@c�3mV9q�1vA�M�I��X �"b�WD$#�oli���vҎ�
�R<�n����#t�	wa���C��g��cUrW=�����ݨQ��Z#��*�h��?��J`���Z�|k0��bW�L�'0M��o�<���/;��|�k��&N�E��e�_}��ĸe���\th���d�<B�R�2�!h#��85�� �!�WH��r�W�ov�`��=�Z^�A���hU��� >L�>ubK�x�/(��+��?�X=#C���~��������=�ʓ�r������{1����>�s�yT��DtЭ��r�>^;����q/�^ϔ�q��ؚ}��3��[SY�8������N
�0���:�!�3�ƽ���}��Wδ��c�a��,����=�&݄�ak�f�w� >����-��Tsɂg�j-�l|k�J�@�Cb����ɓ��❄Jx���w�}�o�s�؆�[K�33����I��T��!VV�Í)P'?=��U�h���!#��� `�i4,"��E:�ɓ��6'Ǟ���L�b�?��ŋ�����[oͳ�GO����cos	$ݲZ�B��|�.`X�������ۂ%�9O)�~������6��8G���$�V���5�T�����G���B?|8KO���=�m������������0����`́����I�:�t���-�^Γ\��'�A>GOh��x�����Bp������_s����Ir�&��;����߅��{�<���[J�u&u����@V��f�̈O�)++��8��K[�n��ӭ���q��^�V�B�!���ʁe�8hL�����S{��{������H�����2��NDXx��z�|����s����>���5��/V~���!�l�~����S��+]k�?�w%�+�	��(}��gbbb)(�P���6�����EG]]}n)+F>�lr��>��%��Y+�@x�Λ.h�a-Ɠ���,�Nd�d�-���]�1�|GD�f�>~��#���rc�A�ׯ�y���!���NNZ�K�����{�u��rT�>~T�f��2Y��(yU%Al�;9�Jo��v�1#����37AY�r7�Ÿ��8���A�+w��r���" ۜ䆸9BE�ǹ:?&��9�!NNcu��4j�B��wM
h�N��ᚐ��-���c��~�ߟ+d���z'|���'���=o��);�[@?�^l�A��n�<��S�R���n��Md��Sԗg�{2�浓q*GCoGw-+))�O?Qu��ө���ߪ�㪳�����a\������!��t�ik�3Ǜ7����(rssy���B����(�JJer�տTs񨬪z�Գ�q�����Ruz�p������e��_0Hi4vw�gdd�z��IF&&c77�	�A�������_AZ�-,�~2�iΰ��:�#�ֈ$���x��~�x��T�^���hj2���P*��(`�)g����%��� ��?0 vt�PXD���C�)Gu�8�c�i0�Y�vi�7�n�A^[m(���?����DDD��3L���:?d�VCJ��t���cg���V�E
弲r9������\J���@_כ���g:�m�w�^��k1��e?մMdh_.��aqqq���f���#�CC�O�ͽ�8a'WE�r�)�\���
Vr(13��R=e�F��d�G�,��a��O|S�kOP2�Z�V�<�Nk�K[5�\v�Ƕ�ՃuJiP̦[�s3�t��L-BnEۉ�~��U��+�\LoF�T��@���/hFJ����x��������#Y%��A&~�{���KcC���Ѧ&;yUu�;�gf�NQ�O�g�n��M�.����F%TTW��d�k1��`�-����'<����ɹ��E��1��_r�q�Q+w�[.��E݌R!����=����$2�ZU�T 
a�∦3��2	�6��O�32:)�v��M2T^��Z�q��~���=�u�i�����`v3�c䲚2;��^�0���C��S��]O���
iY?R܉]9R�>H���8�A���S��E����/M*��<e�U��jZ��ϻ���S���{{+���Z:�����t}ӌ�`�L��i�z�ܦMOOW-�9�r��o�����LM��l�n��3
n���B�Y}���gز�c$g5٦m�w�>k%�H#E���>
}t�!ź��lfƣv`0/~��$��ݖ�b�E�:�Dzgj����z2Z���<`ဖ�~�ݓj���@�C��~>����C;(Ox>���<��R�A��������5��c����W�l�>_�I4g�G�3���{ߌ����CQr�E��B����V)��ۂy��p�H@扐t���H�N2���d��d�I�*:h�i��_�й�%;�a-<+&d���O����o
�ٚ�\�:Q)��B��I���޶l;�Ź���O.&4T�i��c��W.]w'��#�E����>(��\x�2�P+��.�	[(�Ap �������-o���P��ȳi;�t4������om��n��k��c9y0%����G%-����\�
Ni]<��A]���e[�� ֩%Q>��:t)��u�o�	ռ��(��
ְ�����Ns�ܝ/Y�Em{�y�*ɺ��@Q�wE��X�s>/�Ͽ#k�D��r�hc�ƶ��i���\OV:�ݧ��2C��]�2��i���i����a�|~~~^���N��Zv�����!����8��y�����;kY�k�jѿ�P��ᱥtH8M�aX��w��$��!A�б�7�����+`�/ �S�'Ӳ}SG��������_��w���N6 �W� ��Z-�^k�AҸN5h|���3���bf&+�:��8Q�q��TT��]䧪	S�b��J����5��i����=*"�	��7H����%%����A��c}����>+fRqɎ�1ݞ5��/5�e���`C�*R z3lv�{$�Fm�O]y��)��)s
��{�����'�u��W�p���rK2$^/�
.�i�+Sާ﷐��2�Ӗ�ҝ��$�w^,��D��^����W�2�0�k�H% ��?5�R��,'�t��,4��p�޿M������{ )�]��BY�d�*�@BH<(�9��f6̤*H�|j�Ce�Y��(�Nj�Q���{���a՞x}1%���hK%�^y�u/��@��H�ר�h~՜+�uJe��,��v����	NB֜p����3�(��7fW9����zí
�cq�ҹ����䅅힝�	�	�|��1���E��SEZ��)�̳c��Dvy�����.ԫFF1�[b�l�v�sS�G�X���5��W}�	a�VK?9�hU��$��@���@Su`,�4����M~�x|�k�@_��IƉh�u�O@�$9wƲ#�[MM��/m!�	��Y���7�҇�dd3���qcע-�8��7�����΍��Uy$��wz(w�@�VB�x��ͪ�g�����fy?ub�t� ��s�ý��S�aE��+h�w�\nll�KH)x`�q�%�P���#�.GiJt8
�Qr_�6%G�3Qh�V�#���$	9�PIr��1C�c��`0��{T[�����w���Ƕ����~�����z�.(u�|ك��)�/�NW	 k��6J��c������w=A�p�cgQ�U.���ݦ{_�;M��^-��](w}v@S.�"j�M%��� �`��Z��e���ʣb��9R���7�����������p�F	���LM݀��]�v1p�l'��2��( ���A�«��6	#�X��|����s@�+�33o���6zs�-�}_nn��'�ꩾJwU����u�ӣ�O�6�9qh�t_���(��<hmG+��d��M��8 �����6����W��$́���A��3�L��~`�+n#Ң��M7��@z�5�e��$�C�������kc9;[=_/�*�j�<(��lS@��|�v��A�я )$0Z�P���]��`�+))��5��n����� U����-?6�*5K�%����h�Wy�T�N|�� ������^rT�U�#T����Jo����_��Mml��&h͕�X�o'�X-�\����/_*�G3?3Q��SHD�F������s]�
��P=&�S�f�r�=�Z�_�1���վ�S�U��!��ʀ�9 N��C{�*�X|��2��p稽�x��ɳN>�\Nb܆������s!�W57���>
b[��yKPHzbH��+������=7��|��5`X1 >F���MuP@�.���0nM��ﺲ0)�24�_jȝ>EQ��wt�{0���±��Փk3�Ï�65�ݱ2�$i�'�F�������f�ʙQa&��� �~�^���q��O��?�H���R�P,W����|4/'⩒�(�j ��=o��-�9��K�@�W�
L���dq+��E�� Xt�$RH�<@��Kq�Æ<3��&����8�י��ك�"IӼ��}�+E@��=3����f��/'� �a;����S�����c�`i?���w3`��w����Ɩ���A(��P��
��p���>?�ذu��##e��������r@�
����C�W,�%�x��l�~X�oɅ�)�ߞ{p��U�#���"�� �e�,����<ܫ�>�M��i�'�r�q ����K�wJ���k�������4��jK=�>��m�)��o����jeB�G|,�����i���������LDc��
�z���H��*�l`��V�Kh���t�m�&�[�����j���a����r�\ ��QSS3�ճrF�^�~;�Wd��C�7>P�[�6Ƅ7��c�<����=��O?�pKꮟfHi�� F�{����3쵑�7�����
���Lܟ�|�;��U���&�������֮!��ݳ�.�B��%����^By+!!Q=�)ǒ:�h��X)�N�gx�yۯF�y3�^�OD��l�׽������ӿu� �?Nr]������G_&���%M��H���W�E�%��W�ߚo�l_F�f��p	)r��<�	�nj�u�'I'癙��/m�z����YJ_����+��l�F�����ࠇK: �U��"+'e"�p$4� ����h�j%���6*}*�kf��;s�V������|������q�������ٶ���{)�Ç���e�t���T���.�~���w� NIx��F��<j�������&����/:;?�v*m�w�fk[�f�����U����j77��t~�� 9��q|P#.��0��e�}����/��������W㱎��D��� ��y���U����:�����~[�0Q�NA�rV���#4����l"��^VF�dd��k��W��VY\,a�Z\�����s���蘘Ѐ� ѥA�(I�jC�հ}Y���{hٍ=.̖�$F'߱���Y�N�Dۣ!�Î�NrO�(������v��YϞUG��3��qp0m�RF�B-����r,i�V�����â���Ϲ> �����팭���0 �����������Ǫ������w����u�u�PKo����Zb����q]������+�n�9D��;s�� "�	 ���k&c�OI0 3�]d�X�q���U��Qᵈ���
~`x! �)��������@�ƾ�X�x@Z@ԓ��I|	�c�I��
9Q2�E~G���g��#^u�]F>�$"��P�l;Xn[+oy��q�V)��"��M�v���N ^��v����\��?�Л�ivdۙVB~^p���LY�l݅7��ͽY�L�@�����^���Bc�7R"8�\��� �^��W,-U�c�ΐ��<-~�ղfN������Q�RȶǲWwӪ���/f��>Tv�(QWW�E�b�W� �󯶯����i��a6k��+�I�f��WW+���-et�U?~�1��c����_��-����q�3O�:����7�����g�эc'����2�xڟ��e} Wn��V,O�[����c����˹�?��8�>��`��� ��b0\[�:-/�;Hs����={��i�=>L\!j�{LLL`s}� ��8{��[CY��|�.�7e[��vv>��Ѐ�G��T��X�}Tϼi/U�5������vM�B���n��IHJ��1uu���z ��8��x`��L�ĥ�=??�{�g���*������� ����u����8G~��[ /�����"��j���%���S���VJ���N��/�yzYK⪪�p>��^3ccO���۫fffՓ��%�;��۫��ҕ�Խ�[Y��o@��q�e	�]�|4����D��/#���6�����Z a�06�{��nLxF��i�������������ΤaC�E��e�nF�;�Ӧ�1zT|��9 ���\7h}|�� ��RލM����7w`jzz�@?�x��$L }O�>%-��"&�Knt]$YBL��u9~��U΋{XYYP��=����&`d��/"��I��	`�?���}�����nf[He��o���F`+Ma+v� ��]px<>Ɉ���K�<B�q`X0��#-��i��뽯|�����e�&l�����d��W#nm��Ow���ǹ����9��PW�(T[������֓��6�Ү��'mO�ʁ�- {hc�+��ve=}��*T`����{5lb�����^+ݓ�[Tص�R+�\�4��s)���h$�3��V�(U*�����E^ɫ%!'c��e je�;4���C�+�h��w�mV���>cu��D[�qkMg:�K���j�������g���_�4����8w�!N�oh�144�n�[��+s7 xP�V��6�Z�Dx�Т`Э�T�r�i����t�z��w|~��s��iƌ7;y�4�6u�0whge);=ee踻�5թ�8
���ި�+�v��U����a�k���a����i�\���=,?��0^����������vO԰��U�a��b`-�l��*��~������M8j���}�ڭ��%P�ζ>�mQ�& }\	윜����҈���"	;00���6�'V�b\Y�L7�u����$Rg�`ЋY.�_nW��g	zYՉ
>������믬?�_H=z��kȱ?�v�0p�K�12-�r��{\��QT(�`DS�N,l�O�Uz�<�C�'��g`[ȏ���jD����]�=1��E�C��U�ʬ��A�m�J�°�2I[�.Q�5��+���Ñ�? ��P�tiZ�i~��V"�K�֩gX~X*�X`3U��1C'��Wג��5��h3��_ɢ����V������x�����$t��A-֌�a�����:t�q1���2$�4�����A_Ӕ�l7Tϵ�4� �r����T�Z#I�� ��n���-'8QJ�����m�f��y �I<��m����zY�IF�@����~᳿H�L*���-�HG {?��~Z�Ն�
�2�3���)�7��"z��T1ޅ�CC!?mF�R����V()B""����.J���`��{ŁJ�J6^����M�~�n��b�/\�<T,���bfb��άI��.l��jj��l��j�&H]GҧG��1xY.)�+W<��"H������4���f��"��A��?Wn+d-�(fM[�{��.�\�25�f�E��Ti���������8�y,�@�Mx�$f�+ɈjЍ37_����bkR5>��u��m��<�
�";V��}�x���
�*�����@{�0�W�]y�c�ka�����
��bك��e��Z(�H^��;�8��ڍ�{�H�XL_mp����Kֹ���0"L�7��>6`��w|�͋��[+zc��C^����T�?v7��j�7����}�ƨ:�c�j� �܇�&~�#�*=���n������,�����s+�d���C6�u��T��<����߃�9�Z�C����{�>��.v{ &H-��+_��I#-�e����]��؈x���'�n=�<��x�^��сw^�/��b���T��4�.p4�M��ivv�����v�e]��i�&������l޿,8###�H��Hٿ[�� ��vw�y�.N��d�m�l����'"��m�D��ӳ���2A���`�&\MQn��u�����ۍt�ID�`���$���o�Y��~�����@���7.�FE�5=Uɝٰ�9�{e����N�V�4�b4Џ�9=�-�-������C�~�L���Aph�'��@�N��S��aO۟Ys�̙iXu���N�Q9�i������Y�1����x�ǚa咣c��������[��b������8�<f>���?�\¤=��/ޔ�
�����J�����W2�0Ң�:m�ߩ�����K9����?5$�U��>�E%%OK��I-�x�3,��6��mؖ����O� ��2h��T�2"����8�~����c��hn�%_��A�Ic�H2R��po	߳�Y��V֋��xds\��ZΕ�Aع�EM�y;�k ��-pѾ�G��+�����KkFA����xGx�J�c�Q����p�G����]�i�Tv�%�N��ی|�B���=W/��œb�(�߂o�e��wl��b���<�g� \q����S~ʖ[���d���3��cr2��Z�0�}V��YO�֙���O��ˢۄ,ye%��:�__��m/u��-�?��v�"+֒94�+�6Ҁo� [*�n��Z�	@�@�J��ه�R��.���S�!Qu�����������W�7??�1�-.�Yي����nR��9%mR6z����L�)��-�H��+���;"���q+՚~D^(��7߇)en�ҍOP��>����[x5Y�:�'2�.25��.��m��#wX��;�bE��0�5�&�#�*��N�.��.��5:.��;�蘹q�!w�G���7�L*s��>١�2�iԐ,-�4Y�f(���`օ�w�~ȵ��q�3Sv����;<����2K�{�:�Gh�&j�)h�����U�@�D����h{��s8C��Ʉ��&?B�K�dr|���q�ȵ5�������mx��һr#�{�k�;X�@�iv��f�����������]�Ƅ0�jc�:��z���*:�A���@~��ʱ�ӵޭ�홗��t�����f�<�+��щ��%m�G��$bJEn�U���a0ڼYj(V����T�r3���22��&ƲH+퉬s�@/ll��}.+�N�9��&*���&�<���ɂ=��V)_/��tқ��^fH
Zn:�W*B�`����7d�7�٠��;/\�ȐŶ�r~>�>߽�ǆǟ�n���`V!��[E�z��U��h��Htt��
Q�i�a�3��8BtdQQ�0zV5�1@��B��n��f~!��0|g�p[I�R��<�_9� b�BF�7��1�ӗ������c8$�0�E�t����=��mV��X��vޏ�ͲME-����ЧvX;�^D >m}s�m+����#�ye���T]n�Y�y�b�Lk%-Vu\�a�s��^��p.wp�'8��8aQ�K�1Q)��NS�0���O�踐���Q���h{�2�g��#�k��0��xهk���^)U'��ϯ5[*'�����ʣ�<�{��>�هߢ�G���P��g�>�Y��%s$�c)yB���Ǘ�8q}\	 �{"EY�Q]�(��#pw�_���@��6��K�ei��O�6����+X�e�_ȯ�!z�7��UQxݨ��c�7Û�en�<Zx�e�Y�ph(C�����D�N�&�3n�f�րi���o���!ħz�ge�`dԈ*}���'�>�݀�sK�$��m�uy����NΎm��y�>,��Wceee��_�d���\:�ٶ-95u�b�n�	I�+��iӍ��}�\3�;�ofN����l{3�D�Tٰy����ƀ�nG�$�ȓ�`�����o2G��_�y��{�_�ٔ	o����{)_O��L�ԌN4`y����u�/8S>��!�I�i�'���܀��:�VC�*%W9?p�7�gwҡ쒐q�\O�0�/��X¬�^�Y x����Ì�̹+]��������I.7��
�	����+.*��"��~HkqX��,7� �`�n����=Oڬ@����'��D���p��� ����c5���l͢R�V��S�*�Dzκ{�g&�������q=+횻��2A��;f�jO���	^.�+�2Z��}��E��)��G+%7�_v_�A-����{�����i���6l(ߢ&B�T��@�U~v�nZ��		'~���E!���5a6R�w#s@ڇ�]��1ap3�N^Xp���6B������*՞��:::��*��ܹ��[�X��;�^�E� �^����k!&-�|eHA��!h�X��ʫU��)cn�&�`$��퐻rԅ�MI|?Ha���2I��eц3���K����!}�O����0F�	��H+8H�,u�������b�sA}��Y����m�L���8�0��.����>����c�lJ��'�O���	=~���V�Y�|s�Z���;Xμ��9P;� �:^��n��l��͛7�����V�<V*ɩ�!�@rE(r���6�Ti@,=WC+oۣ��=�E,�/�~ɪekWQ �]��[���q6~	HE���tV�_m=9��p����L{��r�^� eq�9ϑ�bCa5��<��,6�lGe�Uj�{�XY�}y���$��=����jӵ��g��2���Η��Ne���f����nΐ%u1}�j죩��(�@�*݊��;��ک�
�(��s�0,���?�}�(�=��D<6Rn�aP���㉚���C�u�z��;�o��H�����M/.&v��i�����e����⟯8��+ 8/gBj��W $��:(F��.��=��:���|�%�T�ϟˋ�����#�CYv��z��)���6O^�
���0G��`���FG� �G*Nͪ��wX8q��V0�ޱ݃�ʈ�|y��Ju�H�G+pMdv�u��H�Si*�2/���2��=�o�^�?bo_��D���n��+��nQ��Ω���\��.=�Ep�C ��dF/4$i�~f�� vrDffT����������i�ϱ>|a�P3ݰF�N����{�Hn�I�7*�p(g��/�����l�n�F�X�oϟ?�02b�I����#Ms�N1}4���w�[8lk�<V���@�-�O��;.��U�����, �;JJJL��^���O[5]G��w�����(����������=�tD�H���nU&ˢS_7�G3�\r"�^��y<ձ���4Y�L)������!w���g��b�C��e�~\�0	�������>-�K��-F_ �+Q/���樫ѽ�F�׌�����A<=zT�h���prМہ=����q�.�F�<^����T���	�39�L[SЪ���^Wn�VSq�V+u�k�?:j�^�q��x׉0=�X̌�ޔ��N�xw4�%�	
�YEq���E�u�[.8%b0�CZv*5�f���R���||,o�*<edQ����ճ�.&\܌6���h�0r+SA��ڊ��V�O�y�}�?<��w~#�����s�*�"��h�=�VQ�X:�����PKK���Z0Z���jx�t�!M㴛8�0�g�koވO���u\4r�fld�>���Z��P.=��ߡ�ߚ�i쩪��
���G�役9���p�I��펜����(���"�圁�9���ۦ>��T�4t>Џ��_!�;T���X�f4=x��`��U������#!�(:�@'��"_�ǣ����|�M��b��JQ7S����5�(�� ��*�E����w'�����G�3�6�"�!>��#��<[�w��;�+J?��M��@�r�S⨧Ib����u闊���P����
�B�Ǣ�bG�� E��iSx[�ا�Ҕ�\�>G���䭘=&�^���+�b֎����
�>����JZRR�*{!!����_��!U�m��(�_��=9���q���� �k�~�^�Fss@T.����k��*��@u��k `��m,첤�X��^�r��+Q]��0��lt˩\,�>�}Db�$�ƛw�o�	� ;���uU���#zyVf���Z�e����	��t��4VzW��gn ��fKhM��t�)s���zXI��D ��P�x&�ު���+��dȢ���Z�S��<�5� �t�=��?���$\����R)7wd�tJ�ˬ�)�;U�mD��1���ۭ�W�룻j/:�[������CIT���Z>�Ϫ,j�c��M�܆P���+��Wn?����Db:K�Yy����Q�&�f�R�N��{�A�ǯ���!o�0�����@|�;���[��d2d�X�d6ڡ��q�����Q�^�&�q���<nP��-�����ĸ�].6�ژ!��˽�+���W.2��p�\&�ٜ���W=qV=�A�y~ }y�(]=i������k� 6�[��'�+��#a,�i��1�*���
�zU��PF����FA¼��4Z>�q��C�z"Cb��7�Q!��.�Zǅo��PUU��;�z�8K�q���9+��l��^psJ]���R�dB�UV���+�PG$��b���|[5�����O4�}v7�oQ��1)����?;SO�27���ӿ!�v�,Q/�u=�຾�I�QPH�)�����Ԭ%�LX~U��ϐ�S�"�o�Uy�F]Y&U�V�#�s�:�����ڬ�ʖ�� �=� ���P�G�z�b��e���?��o�lq�h7O�(�=�Ͱ���R��M�ڕ�d��I����С�Vi����8C�	.�W���SA��A�������G�v�"E�(�/v�+��pm��ۃ��M�J䌌�bcÊKn���Q���lRO&��$s/��L���VA��w���r�ƒ;���4�ϟ/�f�sgwT��8�����8ӌ�<$z(w8�m�]&��m�J��莠���3/7���4�WJ���kp疏8L�Eܳ�L+pd1�rA�.����ͨ�Y��'�7͇d��/KE,ݸ*��Z)d�)��MGG+�h������شo���Y�����1AY�����Ύ�u`�|F�k�!ON7`^�J�Ga��TC
K\�8{&�6"�[HĐ�l�jȦ�i���}0���n�I���+e�R;gg�~��Ѯ&�)༓�qZ����x�AF�D b*w�</�cr����|�L��<w�t��]�8��'i���=�Ya,��z(�r��x�R���:�
�^.&�l�Ϧ��3g�<4�a��^�|��޼�Wc���0�ԉ�)Ms�N����Z �7�[�ܽ��M**
��4&8k�.�L�`�aq\Pǁ逭��o�_9��fl~^�1Da�(�^GUu޲������D۵;������@�uB�'l]�����'�֑���fn��bΈ4��5L���w�Eov���^9YYM���������8~��X�-7rG�w�[��%8�T������A�����6�C���nd�W;�r �W��٬sY��_�KɲV��bHP���ԥ!�n��n&�[���Oϣ��I'�=�\ִ��
ك��.,���K@c�>KNUTT��݊0���´j�V+L7}�r��~L�߯!��1u��Ծ����%������d�v8
ݡr!]�� �:rL|8^ˎj��l%���� T�)dz~�mO�G>���S��ǸQ�&����<��	�#�(����SIR o��;h\����b�}r7C]nKU��a�����t����:n��
B�!�XK�@�͟B��,[q�P��3�v��*���L��X��Du&K��lrH�wG&��#�o��]���t���'�k�F�v|=��b?9�o�0�"�>��k+���**���D��Lfۦ�q��rn4���$��[��/!mmہ�|5��� �\N�B���������f�%Cc)�.O��yXT$e�̌��g�k�%��*���;�El��k���#��A vʄ�����MT���R�j*�VBb˅�vK��)=L�=υ�%s�|&~�lOdsd`/A}?-eU�v�gqH�� ~⢢��D>�������i
8��һ� ����rcGly���!�Թ�[}A�\?U�	"�Q w�����As������6g<�-+�����>;S�lB�6�S�����y(U��;.�m��W���8y*D�qM���X���ť���D�����^������ �O��9|�]�����S-P��ϡ�J:c�)&=x3^4�t�*��oq��Nĉs0��]�O��ݝ UgT#>�O����G�����̚<7K7��Ik�B�4���B�'2X0�j����z����>�4"��'
��^�#"�/����X��b|^��d+P|�ŋݟ�uw�b�6�S}�2��?s�V� ���!�"�}��ޒ����KE�<߀o@��yx�l��k{�5xR�c	Z.6Ѷ�'��鱸����7 S�f�mo0�#zY^`[�%��)h9ڏ���/����ע�K���O��hT��>��B������;�ԗ4W*j,G���?W d��`�H��Cst^-�������S[{5��q��9�+�ֆ>�X�����8��Ư������MLLJEx�.��������f�	Qt��7��b
��j~!(�����`<�tz��"$�d��fD������[����%ee����P�lbM¶�ē��p��gk�[��|		��Ç{K9I ;Ҍ���B�߽�f��R�O����͟?'�8��ݒoz^،|�n�:�I��a�4}�H
Z
>$`fZI�_�,N)�8�f.����֭c�ma�Ʀ�7�GF����ó�I��'�Y恂-Trꮷb�����6�~��,��H���_x<6kh+�kե���o�y�&��8���t�7���?�0���+A��� ���\����@�����(������+d���+����(�OK�[����<_f��� ���W۟�2rJ̗>0�$J�����@o9�Q��;jz����"����D�*�cW�+M���m6�:��Z��R@���������z"��`l�L��Y|�9*Xn/P��gn�G���<ϸbSO䉓'���-�v���ܰ�?ַ~?>g�8𨷶����d�/��� W�jb����������b� �Z�>¶X��f}���;s]��̺�!<�:r͙��~����Z����
�vS���>��	�!��3330cL�%kq̙��6C�������x���Ѱy�zu�x�����I�s1F3yZ��
�ZM-Gю�����fTdbC�5��h93���ϕ�5-7�b�㮌����U��������Ji�dhW�7i���r����ap���&����cR��}X�*z7�>tpy!<s\��ł~�a�I��H���
a���-�cd5��Bjd�cЕ�6�u�۰(J.*9'��v��_mo����FX�s�˖�#�+>k��n�a�P��#�� O/�<ŹHr��:��H�	&	7�� ���g <L��N7n<�3�A����5�S�Q=��3�&9��Ϙ�1g������/ͰK�)��$����y}4��ڼnT�e�A�&�^n��-NC2/vwW�^GG�x#��a�)a���}E�Y�a����O�GZFa�jt5�&����S*N��S�N�v�|� �@�����8���/�������]rGY���:T����]\9��kkR�,���߽��nH�Cr����c��W�C�����n�����:N̹��W�Dϵ�o��]��CNT�.�# +��� *��v���d��&:D2�c �r�6�WgF�
t�
M&=9{P\��(�RS��^<qQMDt���@8��s�q����͏D���2O�ډV��˺�5>:z,�2��^#����	�ߐ��'�x����X�a�w��.��:HnZ�Bm�ݑ���9����#UFC��wz��368��ZZ�v��b���%j����/pU��e���}�2	L����)�c�$����O��O�G(�`a:!|'SW˳u�S��%Nz�r!� �����w�HB��\�x�0�	�(��\A�����W��湐�kQ�˿l��J�x��_m��r҆��l��D���_Q�z�щ=T�!��5�c��&�I�q��7�x�pQ٨�D}*�iҙq%Ǫ�sg����۬$b��8��9��݄Z���u=�J�˗o�'�>\訂���$�;��'L����i�-\�,uö_\��Z�����
q.:�d��i��Dp� ��W�)Zfðm� ����C��_��I�jb|�==����rpL�w^�.|X/K�_|'Y��ȁ�4z��&�m`�ͨ�ɟ�%�
�2*6����qh��<�����E[
�ֱۆ�����v��TnOA��F��Efcf���	�������5�8W���]揦�c�`��R�~���M%�)�I���`9V+^�E�<�����J۞gR��<��g@����t4���5�N�[�������� -���ߟ4���y�A�œo6[Vr9P��.#<��3RX�L�E�7k��`�C��5��I%����t:�G7p��_1��X�P�������9�/���zB t>�~��A#j������ƋO�&�������"�$b���Z�9����Es�u32A;�)� �vªr��'���)��А����+���֗j_�My^=�	M��r�)Nk��
�*���+q ��V.��/�u���wA#)��!�9X&�~qqH�ԑSW��l!���.&P8(B���8��<Gw�_ǁ�
)C�t�k�?�;��7]>X$��:b1��oi0đ�I߄o4���o/Ӱ��!��#d��!-8Q���������)�ev1��~Ր��"J�[V�x��E��4���bOsg�U��뚕8�E�8Ҳ���p���XB�J����ţ��q�?�ú(Z-`��8tnK���&��G���mf_�.ĩ�}��@��m��P����r�L�lkD}�%g�}�C�_�VR%'��^+��7���n[���	�p��;�M��D���g֯�*Ӏ��ߓsz��n��`�<?��éqhP+�{k�A�_�Prf��%�T��|�l����GLu ���D�����ى.�HػYF8��!�h����R=�'�(�A�b�4J�5~vK;����;H�&�|����bcS��<Ǹ��i&�,S<��fxbe|��#����#�p��씦��ێ�1��X������������C�:IAS4�>��O���h��
��N�_��~c�ܤ�e�"�e*d��� y��#�o���U�B)����`�óS$q#����v�x��Ls��h���[86�0133���>���I�y��tHd�3��L<uIޅ���d�ȗ�촣W?l)q�������p��{���1�p8KS��#��V�b��[���t O���!h��Fs%��(
������a�s����EU��� E�ݻg|&��밸�I*�C{©�e��leVK�����K�=ٌ��x4������jW�w�ͅ��&A�J��ٻ��^�cklld��e��uSv����Q���7�^a�w�g`ڵ�H���8�8�S
gz�{e`���.���/A�e�o����h`��sku\���ZT���~YO\NNN
�,Ox��NC��u7r�(����r���9/H� �������wboųQ%�.�ة���
��h���P��#3sK��Q@�}:, 8���۴8;���e!n�S�v6���s3i۷��&M> n�[�D��}��[H��J\_Sa�_�؎\A���=��s���sr&k�}9�P�/���}.���cR��ܑ��"��	V�@��(��l5��5��CW��������V�:�l� )aӭg/�����-W����+0���n1Q[�ES[�9�u��E��������J����dl�u\l��z y�Y�ؽ{���L�E�����?�,a4�̝�#|0|n��6m�H��^|�R��4mȾ�>��V#�~jJ l*w�X��ڣ�y-���]vU�`��)������	*��ʕ+�0��"{Y~>_������7'Ͽn�L�E\l���0>��q�C[6f�5B�@x�_� [�qϿb��{@*jp�cWُ���#�fv~i�#�H ���w�G�*�&T��6�6,��3E�c���6X���ci����-��/Hv��>�s�%3�;]z_�=���E��yß��p��[�}5����K���K�k�`�9�_�aC\
 �t�Vea(^[ ���a�$<֑9�5,29P���7�a��`�훫�a{�U΍VA�F�=�m�|�����K+��?��U�5���V_ m��͛;3Z��� @��ȑx����(z�\�B��t<�%�z�iWp����<���z�|���E�����z�`^�B�V=bg2�C0���KDc5�]b(�cO�%m qy��KE`?[�����}�Fdς77�y[��Bxy+&����X� X�Z384�����oag��IK�Z�lׁC#�g�SkD�b�Kf���d�026��f3p�
Ѝ9%蟕e��7x���W��EM��Z�"L�JlA�\ZUޟV����)�8����j_El=������+0�8#΀�G9aB��'�4Di�PW�#g��{�z��3�~�Jfv��"�ɘ_�d���x7M�`a��>l�$J���6.-�hjj6}�5ð�S�:���)R:
#�u~'w$�dPKK����d���ߖ��*�<������N�������ͩ�m����:NS��OWi~9�j`y�k^Gc�qZ�z��c�B|-��̻9z���kg����s��TCNe����}���;�§zN@~�tY/�ꏀ� )b��8�H�.�<�|�1"���"�}�O��	3��{���/�X��5��Jj��2�ߘ�����y�1��S~l,�����������u���m7y�����S��I��Z5�6^�Gs����'+s��Zr7V��͉;�P�l�T���4�\���'3�i�VqqlWf�M�xbGǆ�@��T��1��o��˿�,f��as9v�_�5.���w2�I?��1� t�N�oэ�?���1�[�X��2��-JT���>:��z������9��˚�菮�?����;��Wް�����a����g�2���\-���.���p\�V�n�$_+誱��X1�����=nT�����E�;��:�އ�~���/HI�,��:��!��M˽�����<�!�<Z��g�\
����<�>��k��-�#f�݇aE2�s�k��L���	;�p�m_�9�ȹ�70Ӳ�;0�e��\�B�����x���1�%;���܁�4Ԥn�����^��n���6z�<��w�R%K���/�ֵ��*l��Gr>9��I8I�19yXSKK�q�`���/�q�ǝg���v��+ny̼ś�P%=����3 *��TV��������}zWa����6�:����9r�v��u9�o ��V(���ے��쒯wsE�U�������� 3{��N.���zi��;��/m�r>����-�9цԢ-O��&�W�c�^���7q1�>�(���^��!�g)~~�<�j�����YEXp��o�>�un�����&��H"'2�GJ*����c�o}�+`f7)���E��ξ��WV��/��� 
�5~S�o��|݃�c�MRڬNc���e�r�/��*��ψ���������mA�)n��p�]+�
_�=��E���k�jh�l��nO��(tW��9cnh8{L�0�:�C
o��Q��:2`�W�d�^ݓ��8Y�ᮞ�e`�%�mv�{�U>�)6��gΜ���e}8nk-r�{9;e�in�րɓ���>$o�s��^��d	pL�j!|@FI_�E���$eF� ~K�,%��B"K������aԂ_���c@���xHa<V�4c����� �+}{��������[�`uE[N�3�8M�"�=5�6o��*���o��7!J.����4>�w8������Sss��m�u]�H��qf��N[v��&�^ۢw�t%@&>9�y6뜥�����O��6���v#^I����T��#k��h;m�-�e��N���!���y���wㄶU�&" �#���̈�P��&~��q w�K-❿d8�\��n����0n����\�ᜨ���\���p-,�VN����S[�<���~��_pv�+�4��e���:�r��F�x��o��m.�m�I���k�y-xQ!�l�w����*g��f�0����-�CG�2?�-�������6��h!�:��| ���wB�y�c�.G�ݿ�P����e��{�ȟ���x.�C��ۻ�Ŏ��GI}��(����9&|��ѱ�)Į�u��m���t~׭�.O�څ������h�Tn�󔁯�F�j�5-v�Bil�����E�'o��4��%��cJk�*�=�@ݱ�Q���5�b�fz�͑��׾xj��0�R��F����r�[���]��p�oӑ����՚����xt۱���V��P<j�
�eJ�Ѿ�Щ����w@���,Yq�T�T؋s )-=qU"����>������:�rY�Ŗ��
�tQiZ���#�c���I x0%$�@ ���Q��^�rx/����Jn�X�Ѱ6��{�Ě�� ��ν�lI�'5�ڠ�*m��*-;�ǵ��������BD'C>��xx���:��Q���-�5���
��ߌVw�Uh;
�����P7u "���t��Z| 5���T��r��1U#c+����]��ŀ�֙�����Q��G��%}�ݏ\��T܎ak��J�������o��m�.�Z���&A7	�-k�&����1lB:.�pP�Օ������^�cgO������i�Rٵ4��e[�q��o�8�$�̾��2����co���.4��JwP�&��}wٻ��n�C�?�H|/WqD���f�'F넉'^��K��ߚ�@�(�r3џ���+9�M����q�«煋��;�����.?m��'\F߿b7}"R��6�E׀��C^��<�eq4ovxv��iH����C��PM��@��x���yzB������*�ae��VóR����®u�xi����.��ͪ�+��~�tQV���Q���zF>��9�y��ύ+6�}���!I�Z*��=Z���S\Io��Ž�֥���Z��ŗǜ�xH(�,h��Z,�6���L�d�=��TU����e�w���=��	G%%J����2��Z����@=999�*6��Y<c�>�'��n��j�Y��?.0�c��j�3�bl3��R���e��r�S��5I4ѓO}��M��et1e�
��ȕI�4�Ȝ���:9��$w&b.�,PQ���'������Rx|��#�� �[�G��E��!8 ��w�<Q�&&&���_N�=z��q�ؕa�݂w�ф3�# <��������y�>diĻ�^��kIl*�j�I�(��ڼy�3.'�^5�?k0�ie��pI*����p��q#�%��<
�B޽����qE�y�+��p��7W�&��[�>`˟�K�tM]��W��uX���CW��N˔�#є�C��o·��>���ͯ��|E�B�sx�/(6y_Zw� �w���Ʊ	o ��J����@T_W��#�~���\q���j��=M��?�)	v��"�b��&V�z@׹�-�@���N��hlR�ք���>�gZ�C����X�D�&�uVT(��9ο�Da��j����*�rO������h3��6��;s����w�8w�Ū̡ՠ���#��W7�5�D�"�U�����Es����X/����L�lC����6��?����Z��h�"����cI��E�"%�PS!����JYCҐ"I��LL�d�(f&�I�L��������=����5���6��s�����{��֥����=�H}�
��X�9/H�c�Ќ���X�
���:yg2����TeM2 ����]���S���T�,Ղ�]��M\�6���Me���X��s>�N�Y48�������W`i6���*b�>�g�$�իW�4L��8jXέ:�1R3J��"���CL�ID���[�z�a[�x�V�x@y��j8�t75��٬Ȱ_�N����G��1s���lmuuC�@ \�uZ~��HAS�r�q�i_i�K�/��8v��W'�GG�LI{:6{�ѵX����~6r�J���̞G�,�S�Ģ�	M���H<<h�*/'��]��������s�<<�=�Ōv��ݮ��^��v=�嫹ZBJve�if9t�C�T���.���t�����ڇ���]sc�:=2������ʿ�f剗����)K�Or-Mj�䂞xL��oow��.�<��J����eVcB��T��*=�hB���C�V�����=�CM�fSD�_NJ��n�j�op�Ӣa��Q�"�m@C��/�v�J�_� d� UO4i�85�5>V�A� �g�m����䖼wwŬ�䅺7�kF��5*���9@�]ųK�8���r��!W׫�bb3�ݗ��Uߨ���`!FJ��X����=r��$�U��1NU��ï׬9-�@?������a����I��ɟ@@��Iu �O�J �F�~b)����{fk�^��"����� ;+qڊAoUӛ�&B�g��+ct*�q�w[n���.𥛫�&x�< ^9��9̢���]������t�l���n}�8�h��s��CiՈV��%a͈�/[e/���9��tL��K/��P�ʢ򀠅�f�m�m
�H�p����[C$��}�:s��KVf����Mh&��c\������:z�hS�
��	n4���_�v�ӻ	��~44׊���j�=��V�z�J1�
��� iD��4�,�V��V�z�<v�)�K7�����F�*��7���c�-���M
Ǔ����(K�mxj��Gu�3� �f)^�e}���F�^�]2��Ke�g���B��Dk�Cmګ��#��Q'�=s��i�Y�h��w>b$9J�#�.,���8�Ǒf��B̊0�"�1+]ă��4BU6�t\���b7l���a��|;�Z��:Ds�zM?"i����#�m�Lz�y���}k�+�E��
r(`S������#�-��ہ��q�2f̵bBІ)� �̸LG��GFP~�=?�pu��j����a� ��W�;�!���z�	ү&���{������C�QR=�]�X���^���5� 2M|-Q���e�TGS)�Vg��Aظ~��}Ĉ+������-�c���˙t�f�,kL��ʵ̱�6y��?Bbv����GY߾�j����nZ�f@��}=��Ͻ	�zFb�ɢ�x\�������~l�g�~�������6!o��	����;��`f2���6�^����mR�#��Z|N��Ɇ����O�V���ܞu�F4���#_��G���D�B�q؟�ɛ.��7X7\��DOx��G޹_J��>̻�"b�R���\D?�M�4���9�?���^��RY:7�S/T���Ѣ�K!����)�+��H���߯v��B�
�Ŝ��)[P=Aдx擘�j�����[Ue������<f�g]��W�tH�%f�o�}iՍ&�|{�;��Kx��%��Ӕ2>�ۂ�����ĂD<OJek}
��1g�*^u��U;D$& N9>
5sƿa��$4��f=j�7���Z��ƹ��&�v#���j,"�G��̆����4�q���\���y��N��ӯ��X���ǋ�Ta���B��'�$[�N)�68xkЯɌ�\�]p�>��P�9��б5��Pd��a���=ڎ�&���"O�u;F��K���a/�9��$���/G/�f�n*)�ŕVˊ}�E��@�L��[��ľ�8�)����)�P��"�*Yqyl$@^��Ԃ�@u)����ɰ]��_4�E5�(~ͫ^@��jKs|V��l��jR�qc�ڟ;���6x4i���K�ىY��:���Q�@�������wr}O*2�Z66���M@������iuS��,h5	�	�w��뱧H�×������ϒ�wI���o�CZ3�K7�3^(Ԫ/���0� e��$��ԾֹXL�o��E�d����א 2�[)=�bq�X�z^IQfX&�uN=�#Z�mob�������C��.��3�c����\~��?rgliү;c iHO�Å���,�	���kϓE�a~@�X5�O�lY�.�(���sq�ۯ��ƿ?A4��t��|�ʑ��ʋ�0֫�7c��Ⲵѻx�滗E:�>�ɷ#aV@=�իF,:*��E%����´b,ŀ��7 �m�R�g�/5ڑ��I��G�[W��+W�L������Q �}�U���$B{2ᕇ�������x�=.��_�B�`�fu�h������%O8\ߗr[��{Ys����R����h�-z��E��[#�m
����5�`�(5i��vx|��0� ��X��g�o�G(��8��^�v i���;/�Ib|=�.��_׹0���q�w7JQ�q2���op>�S	#~RZ�%���\!��̳��|ݕ��!�c�G5�?@�e�:�W<�ϲ:Ӵ��p�U�O���e3o1r�T-�x�1�e��X}�T��ٙ�K�D��+h���̒HלK:��GT��߻��Ϙk���@gh��gdSm�U�B���a�!����ҢZ�[����:=�:�(I	�Vב�~���^��P���H"|����N�H�g��J��e���r�v�?5&���[-c��3O�_.G�?[��T�;nU��_6�pę�ݚ>�Xo�ܻ�CY��1ڤ��G���!=���́�Aʪ���Bm��;�����&/;�n��W0/p���&q�(Ȑptf��;�Ȝ176m�7���5c �Z��i�˖��YEfW��=_��y�Vm�S1���JvCz�Q�Rй��@`I�dP�)/K��rhiSss"l_%[�߇��6!�D��rx_%��J23�v��٢�Ǯ Byj�7��C�����ۀ!:r�ht+��r���2rx�=*�&7���*����bV�+?�(zdO ���jJ�#-%9�������b�)t�Q=F���uy<���C��#�Jgq��!�� �h��+�Z[��ȉ�-���8N�[u#u��A��N`�d���߽�!��g���muJ8�z�pְ�iKXl��y,��[�7�k��x"�����C�1��x���Uӑ� ��́��'�C�AT�\/�����b��-�YR��\�vlх ��#�IU:>����k ��9<��ʡ�3ԦY����^��a�Z���%��e������`���ʯBy�%S@h�d�b�G����	�iZ� aS{-�r"�-^���K��0Z�q��6!�h���7�ᗗ{5ěoT����Gd�_�����f��G��#��w�XI�!kW.A,���~��b���y�V��Y����w�a�g��v�;#�&4�e'p��]@/�.��	8a�;.�M�<K����(`K#I���I�1!ku�H@���߭���Kû�}�.�m\v<i��َb���SH��H�!�`��!ݥ[$)�k;8��ꃭ�r<.���E�NȉqYmN�+�x!">�U�j+.�}7����b}5����y�����l���ϡ_�ɏ�B�鎯VS@��tw㯥�z���TR��Aj���vh����Pql�t��B��ҹ�&H((��R�W2�R����98�owE��w�dԵ�@���h�b��E����ں���Z �����N�����W��Ș����L�BF"A�0j�v~2R֯�;������+�c�����|& ��CķY*���f_���/G�Q��J��1oJ�$P����ש����)b��� �z2u�~t׭�rk����U���_)V`:�#���%�(#5���'Hպ^g�?�y�v�R���o_8��b��3{ϼ�'�տ�'�L(���#[<�i�G�(\Ucj�J��Z�;���՜�v[�jƫ�?z���[R-X̀���l�)y�tV�j��,��
�Y��Ԫ��N1V>��9\�6@�����Z�
�;HF7�5T�q^���6^�ϙ�遂֟Z7���-�Q&J�+����K�w���8�X��}�T�?���tw���OĔ�����ϔ��*�./��T�v�t��z�tl��n���;Cb�]��[}YR\wC��*V���1ƯJ���r+mΰ6��n�������h$�z*YՄ���ܩڵORX.�'�V�?5l�
~aƫ�.����k)�L�˻���F	1k��=ǌ�i���SQHd��T��Ș��e_o&v����ŝ�M�N�-V*�[�=t��]�w�ZL�i��$�U��D��؉���S6�
��ߍ��+v������vK��i�VP4� �q��7u3�ƻ��l�����䞬�B�bp�k�˓�����K.<񖖒]-(]�U_��TavD}��|����aj��~�Ѻ�	�?�����N%�n�N̺x��>iw8��{���F�9�p�c�22V���t�'�'��H�����Y.�ŋj���v����{?��	�7������$E�S�-��嶺^�M�M�
"�#��i֣�]��Q\���B*����u�ۥ��U���Ք>�(��!�T���WR�z�a:��B
�
w�u1w���`�	�t�	��(�"E�&���m&���;�#Υ$1���L,��*&F����ݼ�rs=˺�!�����y2�-�-0�mw�?����uA��<�?�4���]pz��I��y'�1~���y�s����ս�a�%{=1t�Bb!8Y��#�n��
h�g��GO,_d��y�+;)�X��6\�����O+�8� ������%��>���*�,��J�e��g�Nt\U����V+��r8�qx~���߶g��,��b��{t�W�NɄ =,3�~��[+�Z�j�)&�9�2G ��ˬKA�����	={%�]G�?,�rM���7�P*��^���?u{��형q��T���s�ݾ�
��Q&�;|���A�̨p0�f�0�mB����x7<6�� R���(�3D�~�����B�ѣV��j�~8�����B��,�Y��b���x/�w6������i ��KM#��бF��L/S\u��W�s�*B@U�����r�i��`	%�& IK��2vY5������չ �/*%F���`����̜u���	
.�r�R���hK���+T(:� �S�����||+���NLU�9F+d
1���.�W�%߮��������%�!t���fAS-�q�|������J&-�N;�m)~[,�o�^��5{��pjD:�р�>]��~��3�����¶<y���H���J�\>)�(��r��OT�v�a��L-�jOv���'��3��ź{�'�wDsk ����k����u�K�3�l�y����V,���J�d���Ƶ��W7Z�`�5�������0-8�M��܆�S��>3$�v+�W���$��O�3\�t��������[����~
ǻ��W���y�[�k�b�oɾ�d��nh�;٫ =Q�u"сou��+�t��f��J���P ��.8k���nu������^A�8>X�z�ńr�����h���_�{_̼�cb>!~]�oG4-��%�'Dq��1P� �5#�Jh5�!�9���==lAȔ�i��� �z[�,��Ru��_�ɻ�p�3�c��f�\O]!,o�e_,H�8HC��}=�eI���0��|�Nu�1T)���ӭm��IQ��۽d_��h
ba8�a�D��dlh�� ���R$;��5�d�e�:h�Z?�-�˼�0�a����9m$�w�c���k���+��̓hM���?�D&ֽ�M{{��}�u��c���['jÖ1��?�������
�Q�{�����6,�&|{���3Ͻ���:Tҩ��Ru)�}�����i�R�L��<Sr?{*�35�'~o��g��p6<�����& ֛�JN@�)�_�t�Y?��>��9B	i�#4��~�j@L���R�g°q�N���e��,$hfv�`k�POЗ+|�>z�:�X�b�jg���(�f�8+q�����f�Ǵt��4�)��Lc�9�i�ًS�zN�Zr2w���|���v�����r��[ ��o�R�v[џq��ϊ>��R\Vq�נ��Ƀ�yv�,���$@�AP���������:�_+<�S�^oŋ�m�}R���7g$%��"u��7?uV���s�B�^7�`M0�]��B��I�{�A�k����?^�[�`�B)��^.�=g��x�?��"`���n鬼0�p�ú�*Z;�B���%8[`12��T?*�fǷu�l@�3v��5��6-���A��(�'�bJoV�b�ё f��;����T��a)[JW� ���ȳ�+3�
�BUW'���.��vo���\,@㽉�&۳r���ߞ.�����ޏ�������}�����Ѽ)���<N�I�R�a����ODb�Qx۩��e��b���%�nbCNu+������=8;,��s�T��3�M쮆�fc�7�()Q�������&�LdT�v@��6�WN�/gT@O �F��*�L'ԉ{���M��]�ő�{�Q�'��D��9v�K?��J*�_�d�B�s)��L����X|�N]j��\�c�P�/���ć$?�~��$A4�Dw�ϯ;��� �J���;^u�Eפ���5�X�;�	M��`l�*$PW�ށ�)r���ѣ�٬���
V�@ >D�J,<�	�:*���@6��f��o�Y�fo���,W6��Y��i�z2��z�q����3����E�">��<�03�ڦ�HmhQwE�;�>*t)�w:WD��:�ǧ��g��?�y�y��~���� 6.�����~�Tk��(J�*���ʧZ�Z6S%M���eB*	�Tq[�?ҁ���r��Xቬ��-7�d"&�qo"���=���**�O��su��ź}�z�B�����cCo�����Q��9#��������:��M|<=e�R�t%&ȇ[����W������K}W#�J( ���;�O�?�!��ղ���1@3goS�6�e��;kW�} �I��ZЩ8�?� ��V}�|�R?�(U�I�+�t�:'a�AiV�^i�ڏ�PIg�cjn-��/VWڥK�ﬥ��o&6����$���t�<e~�^a
��ct0���k�h#P'�%��|�h����GN������_,2�{��
eK�
��$_�n_l�{�f�ы��+��t�cg�m��s�%{��"�1���=�~+o7�s��G �!�D�g,]�{X������6k����O12�Զ~���ș}~; �ӄ�������� ��t�?h���� �Ж~9oxf��Y��?�f߃�w���s��_"��FJ(F~�Α=w}`ک6��P���©�����a �#{:�?t�D|�r��q}�s ���:�����y�B"���.x��zdb�$`� �B�*]�mj~�����ν��Łe�{�kQ�]L�����z����CtP(��Qh��;#!o�������ڝ~w��������h�lP��]��/3L�� ��ܧ��ԹS�]Z|.E�6��a~�e�����]�ɋ䲣�B?]���8�+vbJ�Gݿ?	�� ���,$	9vK��6N����b���������]5��^M����
�����@����ҝ5H`q5#�^eXؾ	���Ӥ�Ö&e�un�����j��4���),u=W�.x��o��{�k0h�(�� mH!1�֕��Y�J̐�Ke�j�|0o���B�
<��e�'�e+v#�&�H�E1�Hd�Lt{����b�vHe�q����N�j��wR���k�LXMB�h'��N13���?��=M�V� �v��0���z^�
��%�ˡ�h_tힸ�Y%˟��Ɏ:��1�A��!P:R������8�C�M3v��y6�駚��8��n�!�U���Hc�ͥ��Z��À�C
�?��w�Ub�z���#O����G�٫��{���i-E�]�K�`NO�} ��T�����=�~��q���e|y
�%����z"ӟ�!#wBO}��-�ȤIcJ��!���S ���b5r��ߍ��Hg��\�x���!=\��4#z�5��b%';�'Ǵ���:���#@�9{ŻC�q�p��lzk���d�����Ǎ���P�ݧʾ:�܋C{.!Ĩ�g��/���8�|nS��u�*� е�;2��X�+���	g>u��49Y�*ž ?l5��e.>��t�3H�쫅�_����m��E���M�S�7{asQ��&ߍ�{͛���.+y
墸���׻��)����=V@�kӉ���ׇ� �}�� f'�7�ҵ?:|G�4��U��?���\A�)�����;����u�.��V�{}DFZ;�*ҋ����w{Y�P#���>���9��5�%�;�(ܷؐ��A����cQ�t�M�?ia� ��Kf��ݰg�ٹ}���S��-p��)��t�������ϳ��X��;���k�E~Ї�1�'�N�e��J�?����v�y�}��Ld>�����h�V뉺��pq����|i�Ap�f����Ɋ[�������jL@�vx�6�t0��m<���yi�־H�Q���7�($�Q����NqT"�l��HW���� ��3������|��ļ��B�2��R������_�X�����y���(�j`Oɼu�D�6ᧁU�����פ"�� L��X�B}�R�x՟ZD�nF�Υ���y�i?~1�Ke�n�� IR�]�&5����7`Ϗ��2�����^�^��X]��>���gR�@��.���:��J�� 8=-GVE�^n�L�']��4��T'|
�?����*�	pf��ҧ��~��(�ݏ3����+��=��gjbsL�o���ǔH���Tzu�V9��XIL��a��*|��D��[�9��m�_<N�cyk"����.�3���zw�d�7�d��s#�Z�J��i�`E8H,a�c�*|���h����?5>��-���@l��yp����f�~���d�vM�F��P���xK��luM�{9yyViii�����3�&��չ���Dl����ڹ&|��=cI/����j�
��'|~O�gn��6��,�Wa=�֢P���㕋Y8�H���}����fJ���b�m�?�Q�Ҙ�����?s�u�?���Q�¡P��[�8����`�I��nI�������֔ %Z��T����������t���ks���<��lh���ˋ��.�8B���z��Ƙ��w�����V'����F�]��(��1%�̺��S����,�o���������7yҼW0[|_�������G)�,7_j~���N�)��&<"b����ŭ����)$��#b�Eі����o�pО�7o
�h�!|�*#ث{�^��xXg6*@�_	�_,�2��p>
�j��҇r����hK��#�󌠬��R$���
���dJ�&~�5�~\�6pB�xu�')�os�@���Q�3f��a4k=k��g��}��=�5k�a�Lr^�<�G5`Ệ�_�8'�lW.�&�+LYP#(//���NrPbX��L���\��v#XL�1��CU�t���2�$:>����u��so��0�#:J+�Z�)���f�v�	�U�Q(���f��پi�Ol-����:����.���~����n����=���4Ow^C�����8P]�a��^��[^��6�ΘzW^�յ4e>+{�釄ͦ08ǒ���&�Q�F �p�H-9�UWg�f7؍�纠��6���)��lzb��+�"C�-�Ո�CO��.#�zH����y�����$HS��982C��TE�z~��$�%�C�e�Cʢ7��ق�?��tDy��>j� �l�j龢^,G��{tx�o�{m�s�()KvVz�	|n�#�@><N
j���V�c�׼�<=N�er|}}����l��R��7G�g߿��{�=���������B]��>ޛRZn�ꄽ����ɦfA�vN�(��/��1�ii�y��yBI~Sv�˔��Y#v��fk�xi�rqmq�u�9/�#?���Kv�f�|��3)oҋYG��i�<�����oF�����٩�P^N�Uϭ�w��ę���졔n)�3��J��q�$ڍ�[ݛb>U`1���C�T!p,2X8nC�S@UG�:���d�n�����_C�6zN�[5�)�S�-]���#�L�`R���x���~$�������M��%og�6�ۍ#�r�R�?fpXuuu��hqU�l?�7�����,��5��7<�w�c�kf���Q���<�Ѽ��_�M���0d�/Pg]S_��H!��&���#ؽ���>xLfx��X�U'�zW3E�O�}�����Rm��
߁u?��������]�a�GD`��\w�&o�&W�&��o���p&X���#�!E�~uڶ7�롼���>)K������"y��G���*.l'}mB���������a%������87S�;��F��Gy*)���0)����9��7d�rI(FY�DP��3v6}����!��\�?���L/Yo�M\�
��p��O�
�N=6}�^z4�KKy���\��Ƒst&F�V]�;""����TL�����%a%)�¥[kki	�{�aq��8	�=�,���H9�߽��� �u٠�*{Jo)°! �]{���#@�v����	<�@�s�*(�od�CtA�\?���������Fy��sUՑ����@�ViIpvn��lGR��&2�� d��	AgB*JTN�i�S2<<�ǔ��KQa`��J�J�PD�A��%�m�/jiIx��-�ۼ}�G!]^NΈ¦{� ��^N��D�a��<n^|d���RW#�&]W@Mz�����w����F���vy�y�=��2��Mʏ�<�qk����\B�D��-_+�9D����DAsCV������UC�To�eX��R	��y70���Vu!��g�����۫ et1�����Á���@$�37���6�O�Shy
:��
�N|��W�vCV-D���R��t��vf&ZF�XIiV�������:?�$,�����dO>s�^�ܼK��G="<�c<�Qذ�������W��|-�vv�$�׉��Y�2���X�i��	!����{�m�kx����@zq<ye��)�b��(wg�O�&W�Z����>nv��#~7~b�ؒ�^F����;�{��0Û}���݃���~�^^^^`v:�C�p��<R�������E0Uy�jj�1�zd�Ei�Ztϙ��c${qZ#Ō\p�kz�����Ҝ�}b1����Bʵ��2�)��3�3*�E����������1��vY�2T ��M[d�^��~�����6)P4g$|?�^M����6��X�}�䱨4A`Is��\I��ϲt�4pU��5
<����1@�J\��8�⋄۲Έs�ۍ��N`!W��I+����t�#N�T�$�]Ҷ����=*����1��J[M�E�D� k����ҫ=���E����� ҁ������O��5T��
������MAx�H�s@_���͛�
��ԗyIs9�������m�s�k7��ͬ��r��J�9f91�Y%i)sH��	�[C]�L��� m���[�jy�#YF�|"=�W0X�u���z}��}mч�OY��I2�\�����"�Ifp��P�͎��������0)i%��eA�ǡ|=��Ip*����4��?��p��{oZ�q]��x3vX�סFΩ�SRƟK
^T�x���Р��R�Ē�>Է�o�aI�t��&7yIw���'o:h�B�W������������j�\�۔V-�rwp��o/�&�i�5�JAeef�k*Q?����iao�9�d��W�&�d�����m��d�&��2J�����۷�պJ����V�H��������� �x46�[%n�L��RU����\��a����L�� �PFr6����wUP����ѹ�����?:w
,�*���߷~	��KG_�]�'.2g׋��-%���,`��03��逄uqQbi�3Z5_4��G��y�
��g2�d����#�ы�Ǻ�=����!,9� hj����0�:,�=��f��2@���8k�s<�ܮ�0ނ�rkk���Ѣ��c[�P~����G{y��_.�N��������$��v,LV+�����FQ`��q�";���(�!.���;�|�C�lemK=��;;���d��<�]�2>�����_YXX�e�x���h_ld�[��������K�f@I
yI/
�5\�O P;w! �e�Ka�cxj����i���lҬ�p���0�p8\���Z��=��.�eغ&�o�>1 ,<<�+�Zҕ���1�ض���%s�����P9DpM�E�&u�3����PC!r���%/Ǿ�6`��8f¿�ͦ �+@�H�� ii�eO��v�I���ب6�{�s> �I�����Z�y�Hr���jcAɅ��2&Zu;xT�Oj��A���^5>g����`R�ֹGK�uu�@����F��s`C^� �%�VU{���򤏥����MnI?=�<'V���6�3���Gq�RfQ��U��Ǜ�W0�H��顰�0`��Qc�w�Vb���u�[t1���ȶ{3δ��J~�=���t�)
�jqZ�8*.���r?�-��F^^�Ƅ�GL��D�XS�#�>c�x���NN����Q�^�U�[�����3��h�g/�g��c��"��~䦽2�t�&���"@s�Fq?��L�Bs�.�)�ޯ�W@K/R�����P�(��a�\&3&�B��x�BN�O!3�S��$��$g�g��/Nkik���Z:�bL��g%��Z�﯊l��h�XF��R��f��w`�ųYLI���|㛪3�փ�Kva���R�)|MSKn��w�,Y3����c��Մ<�EXY��K�-<��ħi)��@,��Ot���r1�71eп""XN&�y����o:t0	����z��:��t ��ny9��6����?��]A�aSy=�؋W��2�>�垀Z�NMV�[U���LP�!�miqGg��Հl;Z ?�֮.--��b+++s���;o^!��P��1�
r��~v@Jgz��H��8���a������|<E�O�v���k����*���8썰���;)����/����UU	��Z�����r�3�$������-��d�k��J��G�$a�G���*u��/݁Tx�,~G�S���/ڦ�n��җ���O:]��c��(��,��>�奼�y�ɾ���*h �$�Y�e7I@�u��j#9:-BBB>���,�:"-J�
���e��is�Z�O���]�^[6�rsA��\��&�_�'�,��s���O���ԥ7
�><�M�c ��|2@��A��VP?��|�55�@ q<P���q��2��'#9���B;
(sW��I��P���t@h����s%����aP��2OvxPc�vmwװ[C*�I>�/;!�?�;���Y-��xx6qEaS$����54XQ<�,)@�feyk^�AT54$��=(:�K�+ �$#k�Ϋ��mdl�������i�" �j�4��������/�s�ߐ;�V��N��5O� ϯ00�����y�`Ag��0.߽��܃� /�i���77��l�~Ɋ�����~.�-����@�p�����3�����! �T}�f��~��^��]�!l.C����,�wK�Q�������!�lf���W~<Y��d@0�u��@�U�p��=<3�6 ?Z��.K� \�?7���g���)�����|?T�W�y,t{�$mi~#rUvF\˷���#�=��(#C���3���D��QYH�I?`S���P��誙M�,H%phf�ثcD?jR{Y�����6@�ϴ[�F�m7������G�o j��*0R�SSr�BM����Gt���~~4�>N�GIH�%^�0���m@$�� J�P!	�rKKB^�f }222�����ʥi��`F�)~߀et��} �=f���lj�Xw��C)��ko:��*����tM+�{�z��	����{U�;~�0�:ϓ&hhX�|sG��[��]j��&#L��q2%��f~?v��n�^nW��k�6�2��Ky�f��}b�~���3����5Y9#fzw�5@s����g�}!�y[��C>��в=fi�jj*
��ǿe��|��彿G3��(�&ć�*�.�E� ���o��k���G�>������S)��`+%�J����8��F#:��f�Kyϖ�4ϖƱyv�@t�&��������:4�ݶ,c������V��d�8�7�I�PZ���n?H�Ibxg�`��<罓���f��k�[6Af��f�a>H�����7��B>�{*w����Y*sC��dH����J�qSj@�qk��gE;=�1�,�ТV�($�¶K��Lxi>)Jc¤���w)�;�S�0!�֚���oY��}?��V��=�݋<(�`��+U��A6
�MG�ab�U���4����xJ5�d��4��3W��~����E����N��X��������\Z��
Cɝ;?l��>��^w J�,���:��孕y:���aBO�l� h�4d1��G���Pϭ4����tj^�+�W�Ɲ��,8.(���#����ʢ,�'�r���n/O�h�4��Ǻ���F!1�b�ė�g�_.�BD���?�	@JG��}3�#67��3���C�uo LhqPV�BNN�����hi�����H��
����*����kg�Q����6�֛���Yr��(�钣>,?�:!50�ڐ�4�1�ES���<ξs���{�VvSÖ=dp(�:�:������ӝ�8ˬ�!})ː�7��h��ԫSԓGr���c�-�I�����o�~Zҧ��֫��@=���C�X��fxh��<N���  ��#[xm� IGԒ�(3/b�� q���5���Jh�|���2d ��f�(�}���S��'Y��Ӌe��}��=As��w���Xw
#��/�Qcccp(�� P _6{D%�Q��Yba�&���X�O�3H������{��H��7J�Ez�
S�vC�r�5�ح�{P(,h1A��G�d���ϡ���	�؊��N5�ޣb*�\
��D����X�NW�oӈS��)OdT(�|ρe�ّϦ�غp�v���e@>Y���� *�fˀ%>`Q��#B�G���03-,,�?ⷧ��]$�6gط��ny���l�Ps)�S��E�8��Qm�@�E�>��oM
=f�d.�������3aXG�	�֮}
࿹��͢��G&ES�����ɓ���mX�!�ʉҰբrgM*0��Q��8!{ďf	����o�	h˰X���M�+��{�K�U����E~�F&�v,H�m�����e7o:��=��z���8�{0"�%�r>Mc�X�9�Z���:AKS���<9���YC�)K��۷�\��<�?�HE/t��M�t6�rU�^/9E���铿��J�E��b���> ��,kk�e�2K����q�.b2c�
���ҏ(	�x�Y����xY��|���:���t�
O��� $� ڙ��?<H��{�A���+�ol|�#l,K��q��(�M55�!��X��+�g��Dg&��|�����tz����~�;b"I��7o�s�������I��#�֌:�
H>Es�>��i�) �ȴ!�u9_J&[�S� ja�p���NlqB�jVנ2[�D90��b�F�e����n��yf��y�_q @5yʰ���\�G��Vn���ex��y�IZZZE��:��̯�����3�Zɴ�8�Eշ�|�W��$ ��yl�D���� 7{&�X��J���/�}��Ԭ�w�y�|�g��G_{oe{�;���b��g	#�:F��+�Y:��h�	�P3�Uw����H�I�Ll�$g'�NU�z=�4Ap�$�pxbȨ�J��V����ɓG�(�!��{>�Ds�!���YiG�a����o� �{ࢬs�Ds%',�n���W[D���)�(�_a��t��9|ԅ�f��{�E�$E.�<e����5'�g�f�O܊ᭋMs�=�Q&s��ƽ��)���u'C������7�)�?r���C.�Գ�b�gͯ���xg�؛��I���W�8��kW�y��ޚgsm��c+�K�]����ߺ�k�_����3�fF������Z���M�"�����j��>M1���n7�L/�^��5!4��	UZ�1R�_g��eETN����?�ҾM���|^˖���ՆU�z��Q�Y��U�*�]KS��b�ɫk�-��eP̂���y{n#Y�q̈́un�=���̯�v�����`�e�0�`�V଩}�ڶ2m��wʤ�k{�r�p�[\��s��N��S��-H�*Ƞ�5Ӌ%���׳>b�L} D�F�E�!N���38��?Z}���e�8?��~r�gfDs�Ϟ���Q�δك�K����K2��&ά��k;|U1K�����V�G��#�+����p��'o�ǂ��Ӻe$�G����n����xOB��X�
m����mB�c==�\gn=���?,��5��8~�u�1&�����$��$��#��6�u�6JL�^T�cg=q=k߲�$�V��KH���>�����Qٳ��r$�<����vq�����*iA�q�V��m��{,����l[d,��Z�q�h���na�#@�#޲_��Fs��O�Z�����<3%[�����2u͏2���w����6&�~��8e¯�0��~�z)�D���oM,Moi��M[]���W[�6|T{�̋vXs�m-������;�֛�����-Z׬BW�]z\|��2-1�=-��~?�,|d��E�݊���5�iS�`�e�exU ��~v�����xO|x���F���F�ZQ�l�7ُ���L��\3���Gs��Pٳ�Nt�;lP���6�
!�kx/����e���aC���G�e��~C��5%Y�O9�W5�"����Ƒ��ä��n�r�n��cͼD�x�qrw��y�F��[qqqzL6�0���l��+X���j�G1�Z�M�	��yX�����l�ph5Y�� �%D�P+!�Z+���5��@�b[Sa{^C����:��=�û��m�H�</��yգ�h�P'%+��i��G���-oUe�T����?���E[���V �+b=�%�`5}᦭ ��V���V���]J!�3���U�����(�4o��eJj�k�~CCHƷNfYD姢� ���C�)�3���;h���!Є��)��|?���Q�f�d[ۜ
w�XaV�q�zd���.�@��,x��8+�
��E�G|��M�m��1	pC V�*�XO*������5).�G@^!�~47�00�ֻ1��R^���e*���F��i`��g�)��z�D:n�=�d��ràL+�h��e�	��%ߖ�Z���|��vͷ��ֽR����Z�c��C[�hn~��pF��)S�I�u/����!�$E�pQE;0��"R������i�-���)'g�+s�?u(�'F2%.��W��H�5�	C��"N�> u1.�,���pc�Tj$��'���4�ܛ�5�{����:|��e|�����$�N���l��)���
�G<~���3��ɳ/"_�gɔ/H$Wm]ʻ��N0��ch��W`>�I@�VI�s�eU�{c����b�>�O�?���9>�b�T�fH h97G*;�G2QO�z�]nU����$`�{k�T~���	w�*i�&�YvXS.�|��`+�,\jz�'`{��F�?RHgTm
S2$�(U�M��6G4������ !����C�<�A�q��!����k�f��,�E��m�� K ��:pYb_�e@�E���H$Y�ٳ�0ؑJ�5V�0`��8�3j����[A��`��ݰh.X���j9�c�ݤhġ�.�nQ�*�3*V��s�<�:`�����J�۽�H�<$m���.﨡UlJ��,�M��c;�w�aqD��w��?��2�n:å��Wz��/�$5w�|
UUmL�X�y���ȴK��u�8�>l��8j�����D����UAo�zo��{;�bn�sr.�&3s��h�cʃ�h���-vBȉ�%.����>Xt��3Hh�W��h;w�2����57�KKƸ(u���C.�Dp�D������\ ���.�:������mUW��e{W��86�Ͳ�ƣu���Ç\�8pIop�=Մyb�]@�/���a=+���g���c��9�m�:�.f?a%O&~�J�1_�A����0#%�<_Q�TD�`cv�����?�y��~;^~�3� f?{)��=$W/�گy�6��4�D�H��յ)�/��EΟ���P-�>`ViE��?�ѳJlz�E)�����d��5I��Qu%I���Ӄ��y��7D�'2]�����Y��$θ�v�t{5�:5]�q��8A���W7��W?-�:����,7��cr�w�	F8����^`U*v�=���6��&�lN����I�7�~|=�Co��b�=ɢ$���X�Cj�m
b�<p358D*�loq�)�0������{V���Bw����2���Ϸq8��?9p,�U�1W/��^�\W��,����ph�^(�mՇ�B�� �,�������j;d3��3|��`7�- Y
��_ң�nF�"�y6z�o�����\��̞��a�/m����x)�*�lZZ&�1�]/RYc����JM�1�_H *�
�����p�V��!�w[,�$��7�6f���}\�$��nm܏M���� 'Ty�w��z��PRU�c��\�1��_TE�9ݕ�]�*��"t{�wV��I1Ͼ��s��x��!q"ab�l,�����y�y�:�)�MGX �d=���9���GL4Ͷ0Nf�)	� �F��8��\�$D��ǜ��|Sڞ��/BVW��}����К4������1��BA`K�/��.����񉯎�P?���JYv��qY���m�  �.ِc��)&��.�9`�a�w@8�Q �455�l�e�{�8ɛl�G�=�ѷb�c}��UH�C�,/{�����%v�g���	ӵ����Z��R��#�Ϸ�08������$�Ve	�!ч� �V��Z���g{�7���eSkTTT��A�G�0�4���晫�E�^��Kp���1!G�h6
I~��%��h�7ڿ�y-�"�	w��+�"�δS~c�hQ�
�U��N�h�[m~�}�>Y<�T2q]`�5�w��<ߗ�"�
Ɉ�	�	i�K��)2/wQu72r,�u6�ؑ����{?��1�޽�K)��y�o2��'�^��jn|���4H G��w��ق@��=��[Vv`�벇 �?=R|���,�P����2��E������s��P���C��D7�%�v^�1'��	a�$�F��rz]�hŅ@!ۃy��� ����{Ҁ'�`Dyﲝ����e��@~U��Mw�� �P�����j��{a83�|�ѻ�?70�.]�Q���_����'[��V��XZ����[	��t�ӏ�_��ǹ���)�f/c��y~ȅ�D�IG+�E��W�*��(+a�q""R6���\������)'��"��u���� k�����mm�J[�Bk��Vq1E�Xe([V�8^�Be(B���"RK-2#������D�����$����_W������y����8�<�g�Dݬ�p��L$�`Y<i��͹�3�e��ĺ�-uJ���<aV=���0���M��t&��V�c�w����mS�-���k��<�=���^@���WWR��\o�V�ٍr�6�R���ե���\[���6��!m!��ORZ�s4�C�o�o㒙��זe�nx|FBBB�����P�D�Ċ���|e���[F�IS0!Y�����z;r+0g�~=w���q���������P_�����
D0�X�J���ӠJIBJ"3���e#�Jj��Y�N������o���Nq-�QN"���A�?�&,��C�@����v����ɿ���#��M�b�����W�G�Z�����R�-5^�|��gC��:��X�ՙ{	�&�S9�zmɵT�2��p��}��J���:�\}���ŵ�:::�ݲ�տ���,�����8��	c[�>�{E��)�À�M>RC*5Jx�}v'��``��Z�#��j������A}�A�$�S��\4�l0��p�C���64D��fgg���CN���8�訹�[)`Ƥ��GF�\��p���"i4Cہ�؋�g<H���+��S�i �����M� ���d�C�_'B (h +:��hT�.�	8�ch�!��F^2�*LiW�!t�:?������T%�) 3�Q�C�K�B�p�?�b晝PXB�~�l֊��-|���i��03�\�s0�>��X�8����
�un�unc�H�������u���A��������Om6�Ѕُ�����\b!��>d��jF3c����M��=�L���$���"1�$��r��Z(��TN+�L�+�h-GȵO�������.g�8L���4�%��s�廂�k���-�vSB�8�Ȫ̐k���!������@Y��D8�d�r�`�y�������g���� ��%;i��Ƚ[0�J�끈	1�MTO�o(�Y�O��!q4���'8J�5�H%�7��F����)8d�� 2[�´h� T��Ӈݒ���Y`�lha������VF���0�z��t�Z����n4�����{3����K4�U`)�c��Y#�^j���/��}�Ơ��{�w�w,H�F{�,���a���c!���>���Q��GG�������Pi�.�|/&"t���k(����1:��۪�'�_����(��A��\>Og�4�"�8��ԟ7�'z��؂$��\4"R+\�����hT���"�p��|�;�q�G��X���KkGIk���i�$*�	j�n�W�� ��B�
���ә�	U�����W�l<�"�;d�)�a����Γ��m�ܱ�o�W�cAr*j�k����lnn6.�Q�nf�_��r�߿N������:8L^,��»��Hmx�
��>� �-�0>=�\��;���F5~�v[��nml0=%� 3���3��L��j���]m0O��u*r�#�c����i�����k;�q�� �Ǳ��yi��6<������0;Z��*�9���M=y�����e�i���-@l��Z��`�����D��N��_7ʷ��֤͚��tٱ�����J�k?���o4*P�}�'���]"��H���`ۓ)(��*#7����dca��b�"�>в�(7�Z��l4�����gw��>��qq3�I��v&C���0O�N�+����U����k-[�Z�5�rRg�ʣ�%��Nx�ਙ��kc�b��h=,%��69<6��;'>��ȼ���䲀���P;!�(�� ���T�l� AcŵF��77?�ܻ6���dh]����0M`ֆ���F�[�����öN����n?�\�X��c�6? O�ҙz�£�-�4����<�4�־^Z���A��n�1Vޞ�H��{��Զc|[��t�#�1�[}�z,z���	��z���|l��|�֏��wi�n@-L��<i�>1V�Y� [p��*&�Y]�>����"�/�l�r��q�섄�ڱ�m�sC���|p,+L]�W�h�P�k��h��P�C�����y7��~w4�Re}R�O;��4Q.�S�5bO�{0���*߇��k�L��0�n|��T�DSV����3kIz"����]��'����JP�#m֦��#?��>�J�g]8�8��S坤��,;�	�6�MP�ãO��E��� �2tD�~�HBp���j]m-�� 9�r�Z|���o�,�A;���&A�,fvVQ�L��8�g�a�z�t�t~��@;���Tp���Q���+n]!h�%�joEW��v^�k΂�@�;:9���74�2H�f��~��n�Q5��Dm�����|tUpp�� �Y��U��~��zL�c�� [���Z'yFʒB�~�]>hv&~]X�����7�*����}��Bs	�5�eg��Be���پ�V#y���j���ۇ*	�g���c�r�ǽ9�ǔ,vG@ȂA�wQ2�)���\������PϜ�N8s�Y3���0����������BD��j��D~>����3N�R��u����fײX�q�D���[����N?�D^\�=B�D�ƕe���oE�|���]qtZ+�h�րB�����G��v&�1$8l]5wFy�[�����Ed��T�r��u?y�_�>�����^3���l��ܰ.P�	����j�-� )���)�t��ъRP�=[��N6=C6u�`@�a��ċ��{S�r�\w?�E�	A����X�L�d�؊����<��T����&�H��!�*U��b��0z��|�z�~� k��u<�Mg/iޖSa%�-bs�B���Ձ�d2�3Y��S	`����,���F�:)�Τ�Yw�*Z6%�z,�_�"�ePX.X�H:�����p��4��@C����G}䗀q�(I�N6S��RY*<��>�������Z%K��l ��,0�ԯ��+5~(�V9ಕ�þG�ӽ}}��_�Ǔ�P���V�Mqw��Mbz�� �����O�+��u��N�b�2���x��Č�N��:;��Y5˴Q{�͐�D�$�t"~:�yQ�Q�ה۟_��j:Q�o"0���1���q�a111�બ���k���?�WYk����k1"?�(<���RBy�	�6� �r����N�wӎ�_����_����v���~A�3��(�g����=Lب�wb51���8������	x��<GM��?%�Ǌ�e��A%��,]5��7x����gѝ�&�����(�P*����@��=2����s�z���X�__��ŶHC^?����}�Z 0�ߓ�$%�-	̑�j��h o��:mc��=Lu0pj���cs�������y��~hb���?m��$G�^��`��:���T�_
|����ܶN�	R��t�Gle�B�
�QR{{x�p�LGF�B�sk::~�D{(BZ�O��4��zS�����T�\CK;�
sS��;P��-��Ix@B,E�X<����%$�f�񙗝ᔏ�wb�CP_M.R5�M+M�_���L����!�9�ܞ��~��>����\�%���ч1�D��0�$�_�M���l��zb�r@���;��7�=x�ժ�������|,���mPܚv����P��=����ĵD
��=�_α�E}SS�57غ� ��SAr8��P|3�G�b߼���aG$��?��RR��\���:�@�K��|<OC`3�"|��d�������!\���m4Т��t����C(����g`G�U�fR��0?�F�I��ml�B����5M���}�������"�hKe�^��dk�oGw-[8�
�>����ɕ�_���N(�ƻQ�>�Z�@�37,
�9�������?Cs��zEm����k�L<ܬ�n+�ut��5;4�
�4:��
�"�5!Ԃ柕������*����2�J�>��2y�����f�u���P?_ˬ�����vX��Uu�<����D8∐��� /�+�7g*~�����iT����/���)�6�x���իi�q!-�[h`R�]�6����9s��S��zKk�t�J�N����L�����
(�<�Q���/B\��h�_#y�a�����V����e趽{�Z'���&U�0r�Z�?�^�0�;�*��I�J�Ty�������"u�3�JP�<���E�|�Ǳu~K�З��D6%��κ��>���PU1qV����&��2z�y:l-q-������L$׵�Ŀ��ՒhS7�\577�)ײ�'s�0������c��fh�0������Q�W,�@�M��q�ϝ��I/�m� G!|���H,4��D���$����QPo��4:wD��������y��	��$�Q���X]��H�4��/����3�a5���!�OR��2�Yo���iႈ��*�r��p�`w�m�+n��������7?�cD�:��~�G��o�A�}~T
^C8��w1F�=-!j���7l
�K���V��H��G�C*�:��W�/B9��J�}�Y��-2RWv�R�
�żj��|��%@���N��~��	�C��7�7����7�bWd�O���i������U����"�7��=�W�~?E
��{�02��Yak�/{���<K�У��A��5w���P��qd�[�+ݑֆD�,"�9�,��N1���Ԥ@��1�zĶ ���.��Erq}k'?�x�8�_��d�{�M��m�C���o KN�W���կ�|�i&;��u��)�2I_�	��;2���J4�!�/�Pƫ�����hȳ�q����e���A#�:�xT��p����d���y��@�W(�*�"�/k����h�>��?Dʨ��bJ�T*�0R�y�c�K��E,�J�p7�l��6/�*�-��C}u�U>��N�W��Zg$��rB��)����)}&�{��Q'�ޖd���H���tt������|J'�����^il��}�Fjם�����J�0�U�־�=��Z�Y]M�m@�9�dbu�u�9xZ]U�A�)�A���!?�/�{�[*G^���J�Kk�l�)�	����\�9ad����%���̖_9�KdC��&&\�{?��Z�_O�0ݜ��8��Q�6���ֿ.g��m�UY�zaJ�'��
�V���̬�0,K�����E��-��K;�m���1[%ȅەv��O��!�H(�ђ(��o�b��BY1�r�Z�]m��մ��_p�X�[C�2S�{�Z�s�C�R����Dn~,�8,u���?�:�4�	��b�2j5��|��:�mu�"/������隣8?B���h�����BvE��x"gl�{<��/��Xݝ�+���������E�B`�Gd��սW4��H�_�^�$�Drww'��ǵ��y�
!���
�9u�Si�N�>�͌��%T�`۲�R��k�����|��#o+�(T1w������y�L;-8k��𺃶~���Ed�p��ѽQ�=7���L����Sc���	���~&':�q%��]�w��g��e�Q������0䵛U�W �T����a�K�h���`qY�I�=Uџ�o�<
-"�yf�ͮ�B����B+
�<�{#u�uA��F�a:.)����D^�[�B(�mV��|~D{4uMO�%�g�ǭT��T����\zyo��N�ߪ������!�x=�B���-��0���'�ۦ�5���'JVM���`�p�v_�Hl����hhh0�%���m t�(n!�XE�Y�^�zKQ�M���S�._�~�,z�AdT���&1�az~d��ߝV^���������X�@C;�7��\,�����3<Q��Oi�ܶ> �;�.x��a�~9ڄD?��z>�U{�t��in���ߦ7�����V��f�.�8�yv�Y&�dQT{Z����C�Z]�8q-��X!7�E�!�
�4��N�5�����D���5Jb��\i��'6zN�K�6�;5=��\�޼l]�����޾x�,wT>/�ez3s�as���ZZz�����Sn����\��c5���r���0�Z�*�NT�h*.T*��Hԃ��w��[�e��Z�%Q��hB��ʠ���������-(^Ն/��Rs���~�D���-��a�&�~8�*��[��#Ճ���ric��k��3������ @�B�̺:�2�H6Y�`(���T3$Y���'����/��*�hn7}o0���_T���چ1�m��(�#OI�슀�-��Չ�6��X��j�n3���C��꤃ϫ7�]��)�%�n7���I8ʂ*i?Tˢ-J��[eZ�Nx�5Fs��Lq��o�?��ZX�Amp�NbeY$�1Z6�:���i	ZD�A�?�ꭗ�����wsf��@���`ӛ�*�#@��23�y�]ї��o�4�2������aAs8z�7w���}p�u���H���0�������=�k��T�k���c�O��|m�o�t`��V��-��}� �������:���&t�p�B�AP>�����tz��h #�(�- �������EŠ��?��g�p��~�c������ s9pâ�����i��.�b��d���J��l�NH`Q kb�l(�TƲн����L*�����x���;���ܚѶ��OBH�)SpI��U�tUx�Ҕ��b\%�фE�&E�ɬY�@`���n���D������]6�a�����sb�h�Ƒ�p��g������?Nx�}��A� }%d+���a���u��e���.�������V��i�7�4�vw:%�����S4w���|��P�rpۊ��:��q�rS2���k�<<Z�`�,x��m�?0�18Ȇ��[��"D3�4��
�}N��ɎU��o8�c�pb�C����S0�FifGI_FS�e����⊔�,_C���q�N��^�[:�3^p�`���r8�OJ^:[���&�h�Q��gL-��k�����U�7	�.���E2h��hx�e{{�'�^e(�3A#Q�3������I��7�`:�;��+�>C|F&�u��w��8|K��=�.�����`���OCz��[�~��d�	m*3��^ȷ_�B���=�\Ж#�"�"o�}h�)��4&��m�;�T�����˷�:)�=�_G�������/����M�cW\��3+��w��b
e	�FK#u�M�)�9�k_�9��
P�Y���~~Y5��4��&LQ�+��vxF�4�+ʢ��p��=Bg�e�UL;PwmG0���u��	_�zg% �-P}�>,0��W�����K�=�R����ή*NK��<ڼ�����?��P�=Y��Z��gC�kX��]*I���ù`U�͟ ggg��������!�r'RO��^�
;��hC�7&è��LQD�-L�0.��?��k�$�U:�E}�/��Y/��nͩ�T���y���+�ڦ- �@��Hg����>�z���~�]�>P u:��,~�����ջ_�����gm������~"2�Ѷ�݆=��A��:o��d	����
Ԅx:x��~� H���'BV% ���ߒU�Zy��*M�z���=LII/P��C�������n����8���	aOum���S����g���l���,N
3����R=���M��c:8��,�q���g���������~<v>�p_aq�#�������bu��Z�ܳv���"O�@�u�X����CE�I��Nr���X����2�%Z�������O�\��N�C�꠽��+��Ș��|ְ��F�!��*���fK�W�=>�J&3���m�݉O�T�����8�=��h��~�딻1J �wo9���A3�f��t��'�����w����Q��;�r{�q�'�---@~���̲A3M�P�>wݣ�K�=D"$pj�A{�������^ ��mN���
߳�
0O�?�c�ַ���.��7�,Gf���J���%U��K<�8xk�k���"e��,/�xIx�+h��V@��L�Tf�s5��*�z4toj���J�ފRoވ��ΘNd����:�'�x\� �E�!�)`i@����_��UQF�7�l��� �����~�H�9�F�V]���W�0���k\g�i`;���w�[ZXS-�
u��v�O�c�O��7Ό�����V�K7������뷵��:��#۸Z�����XAT<jݑ~�&�&P܃�-��7ދECg�e������t��7��h�ó�Ī鰫T�I>*ǝiQH >�c���7L���_~ROl�(AsTZ۔�suh|B&�2 ���4k��d��؋��X��xs��*��@���-��>�5Qo˲С/>�2��o 6�Ǡ[�
w.��'O^�`O03�����>�ѭ.5�\�^�}�*��S���6�GRW,��"�}�5�C�`K�d{�Z�t�W����ք(����nƉJY�Eo�,�9~�R@���ɪp���b�ql(o�^a�ߌ��L���u��'�޻��
S��U��]�}� ���9��7m�띕�MrdI�c|l��Z���н���_��FM �|Վha/��r3�XDrUֹ6վ{��Q�eq�� �9LU��#�:4}ы���>w������s�1_?1T�y��W�V�Z�z�h��Жv q���c���ʬ{�Do�����*��zX��Ր�Bj�;=E�UV�a@Kn�4UHh��N�k�.�/���C�LgF`��hD����DC�/��b�#p�J���OZ��?�Lx�1)}�}���U߫���]�u���`���m��C��{3��@;e��v��05�<1��4��o3.&%�Y�!��N|�A=!�=�}��z��w֯�����9�2���wU%@��j��|~�iϿ9j���H�:�/s�`����� �XR�.�[����l�D�� �Y ��SC���9��SAؚP%L�)�hn����C���h�f�է�Y���')�p��^����B���\��W,ڲbnr�$zKJJ^rrQ�4�tל|��K�P����i�O֔�o���Mi�p8��S?��O��?��u�#���R��-4d#��~�-���۰i���,T����gY����$�I��yݓ��;�+p�R�����Xnx�?��
w���iIiNk���sգ�83�yf�g��6^K��2*"�Fbl'�N�����d!��-�7m�_?(��	T�l��:1����}{��y��D]*@Ď�S�m�d$y襒�	#���B�h@h->�y���G:Eg�=���1.es�"�[�������T�Z�԰�w��P�k�_wM��ȣ@�^��j���eM��D��
�+d���JU�0�p������"Ǭ�-$�|�Sl�U�'\P}����FP���Y|�Y�qYx)��͚*ܖ:50}�+)�O�g��0�5A��PZ�}]s�]�>u�i"���4O�@�<�)Y�������t*���l(Iќ���RbՊE���"��"�L"mI�e�����C���Ӻ��:@D����^'i��TIkµ���_-�$ďߖ����v����e�Dr��ݯ�}r�ӰS��?���T�rCjM���J���	��E_���e>�IudrY��{����^�,�Z����o����M�}թ���u]�����6ہxx]m�ۣ/#��t��=�ww��m +����&��+Xq��;�J�gU_ڪîqu��q+���I���G-�6�JԎ$Z�ΞO\ Dm�Td�D���6O/��nHU��e+���[[�D7���x�տ�;uj�-9^<D+�Ke:V�������ĸ���I��o�L���#1������9o7��9���_���!C�R�����.�3�>���_7,V�����M�VAݜ�c0�'���c?v�Wz1J{��m�(%�� �x�u���ؑj���i����mN�Ϧ��V�ҥ��i,BD}�{*C/�h��j$�!��+2�\�P<٥��sL����f��;�o�☿�鈏�_�`�bK���9���w�Od*���eo�}��N�u<���A( m)}[}v�b���Ũ���\��'o�}=e��^�
�w� .S�<���=����x�͆g��8���F�7�:>���;S�5"@k��tJ��������H�뚜4���Jb��>���r�4CD��R����[6�[��'#Gn��'E�>3���L��x��%[*A&c>G&���C�n��t���qg��t����=�i����'5��eKn�Z�H���d{M�p8��������=��T�xw�af�I.˸k�ϫ�߾"���x??(���B�>�'c�2��G1���7,|b#��B���'\֠;��ʻS/��J��2}e�j��(�l�t$�{�� Ó5�H	��~��sǙ\Y���t{G����=�w�՜RXh6ο��,���q;?_��e� 9�)ҕ���	p�Ӭ5����&�&��_�J*���S]x`��le�q�����LHB�K�Y�l��ZU�_���e����Ճ6����>�� ���2��,���Q��ir^�-y]�NW7���`%((��VCY��Ϳ�t��QU<G����&�i��BQHԳ�Jf���:�5E�`;L�tM�/�C�W�$Iox���V)F�����V��l�����d⌓�#�7`F�o	�g¬9QKp��_����a��JT��Awڸ���@,�&u����A������s�mԤ*�V��9�_�wrj�U�[O=�aFzP7��;/	�:���������dX�U�3� }�Fຓ2�.�Y9z���᾵��n"��4�Z'� ��hh�m��}Ι���0p:���mē�2�I�ϾlH�Bh�kj+�ٮ?�2~��"6��َQ���.
�?�4t����q,��r����V.?�9���(�ij�����ACÑ�}c�]���瘧Sj=�j+�R�UA�kc��T�`����@bh�4�X�~�=�t'�u��N��y�-�͋�(y�!�b���M4"Q[CF�u|�������c��vG�h�w�<��c��qIj^k:���KD��w@f�L6�A�������6����-$�퓉�����얆����U�΃]�k7�����Ō�R�"W��<�"��l+�8�C?C^�	i��9�M��f�6�_b������/3q#BVt��hǧ��4�BqN��dӃ��Ov�9�{t�EF�E���}�y.�R%�ʶ�Ҭ���7͊�tו�5E�7~������l�|�ŭ/�<����aP����M�|Ҍ,/g|�o}M�֛%T���c5qʱ�sK�Nӹ�h��ࡎ~n��m�^Ʀ�i��9	�qf_#�x�o��ZZ�0��\_�{X��|3��@���_&�~4��u� *�a��~��!�#��X=��QQ��u왽7��X��ֺO�+����P��������Qs���^�j>{݂��.a0����{}�6�} �ĮC�4ٔM!��rccc�z���I��W)�iYhg�Q\�x|+SUU�P1���ӓ��`8��?$$$<��z+Z����H��JuAX��}x*��|�m'Ȥb�Vʡ����+�٬H/EZ���s��6F`�b�_2�m. r�y�a��L��v4��i��L�e����+W��'l=��o߾5k�+��8�����li���e{��4��2@�Y/g"C��E��7�í�$�Y�J�����ԦUJ������v��\�'�Qs��=P��}�@�g��J�&�)�R�/��������˗/M;��/_�����䟿j��K7X�bŊ�Tf��/U��
��d7������"լ� �k���F��Y���FD��b�ʱTs1x_R��9z���#xQ�֑�qT�1$1b'�9z�<_*yN�κc'�ܕ�����|�dg5��51�BHM�>{��OG�s6����s�	���a�Z�;{�7c�t�e��������8�$�MY&`�|=EqW�����~�����oh05LŜ�������
�,��s~Xx�V�}у��	໑Ɍ�!�Iԓ%w$d�qus���~��=�� %T:��6HiX�'�.o�#�~ͭ�U�qEc��������ں�T�J����j�M{ ~��^����[(��4'�����]���ǍN�/H��(��gȦ�'�;��.��('llk�=�3�W2��~I�!�)eY��[b��>��C��TZ�iE������|�����o*�ne���)�ɦ������A.��P�]}} �s�]�3��|F�l�����|�j��h4�.����k���.�ʹV���B�l�/�qʊ��)]���1�[���ЕaH��妫�4Z�,�_Ƕ�����D�|]�J�rvs�^��Q��)�X�ŋs{�Tj���9��{*��� ��$x���n����l��1~s���A=N�.�xw]��r5����ԨL�w��7��q|�f��)�ԀK,vuCÒ�y�Ǖ;������֤�
�^�z�-�Mq�![�Ls"��*�=��:?���>a�]m�Wr?��� IM1p�A�X �PyWm�ҕ;�f�W^��X}������۶C��ʊW��X^j'�t��q��t�%^QI���.�l�p�p������������J��]^5ң's����S��05q���A}�&�������yte?�CK�$�)��-���<���'�KyxZٴ����v@�oC���QHs���5�!��h����q�H��u�p�e�Mg���2\��;��yxx�r�>��?��s	󾯟n�ݛ
G����������m�X�[d%-����GbD���Qu�v6�\N;� ��a���
+
��t�t×V�p�;0`�^GDb�V�:H��ȣ���]S�����\�p��6�ޱ"�d6Ir?XE/��g�;)��/�����v:���7�"���-�T }�'�$}~���.>�����]<=��Θ��9'�m�%B��b����|?(��~��B,󫱡�����jbv�W�T	��G��5(���Fǥ��;�y�Q���]���Ԯ�{��ج�2� A����J"x��3�u��'ƦD���,�{���uТ�c��cn~�x��Y�i�u􏠧PSiYhT�|Q�?pS�����x��T���?����>c��u@��;�bA���v�,�1G�a$��w� M7G���'���,9�t����	�6s��]��p�c�%3�ԧ�l�7��;m�n�ן�+=q�8S�b�W��U$�W�(`�~S܃}������c�E�`�hd����������pG�t8[i&n�`8��*��U��ɑ�,�;��d�#����K%� ��Q� �%i`���u��gn���'���s��~�����׀e�~���}��D�iNj����)�E��k�͛�:jR.��~>�V�d�Q�$�TtѶU�}�̚��"[̶����9�O8�W����e��{����Hm܊�ʵۥ@r 瘂"��*�F�r������2䇹��a��E'�d�
�f�mQ-G�wƴ;�>2#Ƴ���w\�3��a�bT�3�j3&���7<\�z��\	),��+J�%�����	�RU���s@��3��E|�g�w/W���z�.���)Q��ė%�/��9[ŶA:n[;z��]-蕸8;�p{�}��v�O��W���E- x��-\���!�sl�òD��/.MEz ���ٷo�Ϩ�Ե�s)����#4���a��k���77��� �P�|���q�\���!��A�Pd����Z�٨�?:���bB�<$L�0�C�T�L�.��=t�c����̽���»��膭[̲Ԁb�������a�
���[�m;����
|���k���7���^���W�,ƖE�i۶nM�9�@ >�ROw��rf��Yq���Iv	KmG��n�7�������m�>p	���Y(x���UdA��ߐ���Âi5�E������M7 �<�$��:4�{��~ �G�Z�>>�B�&�ݗ�X��P���4�mͣ`�E�D��h�"f����{o���}�������].&����Y�'��j~�ُ�Q���ywx�J���!7����Nw+�d]�����B&DYEܲY^�kϭ�<UgY�H�+t����9x�.@܆�	�g��o�9y��]#�֜��������K�>����;P�u���"���9d�Z�ӬG:�z���1ZA�B���"�{g;X_so�{�'�~�^��K�_�P}��C��^���2O���EY�Y2p|Vxp_+����\���{s�x�|+;;;N�l�=(O$)�%&�Yn2P���+��T�!��V���bP�-3i�O?���9�!�O��š�T�ࣲ�t�۰m�j���qG(~�Nu���xF����S���P���<g�r��oN�c�m��ץ�(�v�ӌ����M��I9�z�l��4�Fo�TԷe�7�T��Т��x��K�o}}�E�6K
����A�λ)���<����&��m�sm�2(/zy���������G$�R�/�[�0o��4>���$4�^��ө�Rꌭ��U��������3��ܬ��>�l���"I�w%���y_Y8�F���]]�J��RQW�	Y�!��sn郘I���S�B^]ml좹c�U�(W7�g;]�f�UIS�Q���Y�b��Dq7Q��L�{���e�`;�c�^���|�c2�RXe�K<�)���޽{EV?�Al����B�]�ܶغ:�//�\����r�g����v �}pJ��ą�YM�����A>չ�^X_#�)G
J8�L�3m)���Ke�Y�<���TRx��1.>��j��]/^<y(J�������-Z�=��Uk����6B�O�^���kIIH��E�����a�W&0]F��p��!���q^�����)vm�"m��h��e�F=�b2��]�/��c�E��gV��TF)�(>Y�,c��/��S����wL�X:/ύ��|H�"�u[GP@�+�r�6�!�-�ї��Io�ޭ��=%��k�o|3>yiW�E��|Y>������X$d�|v0�h|�#��ǋ%C!i{��P�lK���j�wB� ,}��m�Ԯ��m�w{�� G���m���ٝ{|����n�����k^!z���O�^�`�U]eS�7�$l���Vo�H�`�iS�1EEE��f��������!��ʿ�.��=��b
e��}��z��uSY�,j����tb�TJ�W7^~������*��w�N����8��~�����D�q�qv�@m����=ԁA}#$�mӗ�j7c��S{[(�(����^��E��u�mv�e#���Q��b�Q�,+k�W/!6���Q�Ԛ��1�.�Sh�����F(3x��k�;�QWڭ�M���kM�Z��n>��䍇��a��Z���a������"��7���Y��>��P\Y�v�h�O�����BI��'�����Yl:0��/<����|Z�rS�kݑ@Q=���������~3<����:�K�K�����-�u2�m�.��[*Z����##�u��a��b��@�1�$�gG���3��{��T5��ʹm�����օ0c�
:�A���XH�z��-`���Ww�m�\��R�d�����:G���n �oGh#\M���
�V�,�F���m5����uhm���A�߿Z�OA��}���if_=���c��*��NĲJ���Z�&+��iH���e��e*�;98,]�SہH�8��<E�H]қ��u�]!�ɓ�G�|5�0v]+f��r���~��-��u���u�ZTԝ�ߜ^�ڠD1� yٛ� �5b5��ME��I���nlj� �x��P�����]槒��3��&���aH��E������px�F���t�F��4�PY~�C]�Zr����:m��GU��d��VO�:�\/�$�픚A�G3-�$I��vW$O��5����L�4F�C����É,�	4@��g('n1���%x,D�1w�"�^=�C�.	������q6sW�������nt��s�
�l��dok�"���A�5�,\V��n�w�L�����yEZ���P���1�����ƃ�{xb�v�*NI�SV��������������8&��-M*ij�����ԩ=�B/)'����EA��d�m�|W��Å�Ȓ������}�z@������F��ȷ�Έ�~MuY���#��G�n*IY�r%�Up�cc�8 iF���VĴ�Me�B(**Z����	~����2�#|����,u�
.����i?�F�O���0��u@&����6Ǉ@�P|F���E6���7�{�o?=�3���xT���=�o{1d�l�GF)�w_u&U�P�E*�n�@��/H{sg�_E2��oI�Hh�B }C	�2�ov���3
_�-&[u�R���s.�����ki��7$A�y�'���CaOȾ�˅n[��@��}�m�Z? �1�]=9h��p���O�ff�?��l;.��L�������9�P���L�&�`���ŋ	��Z���U��7];I�k��Y��t��=���r�p��P(�6��=C��,b˦��k8d�=�k�0� �yxxX�Il���Q�A@7K�mI�Jo��=�z��%�Q��Ą�-x5͛�������
t���0�⺁��f�m����?|y�D�Rѱ��;�t�)nz�A8$�6�����h���
�Ào�Y1-T<�Y�e��򾻬���ܫ�K갋9շ����M����ON�T"�ݜ"hA5#/����1��V�bQ�z���<"[q�-�_M���2I�j�S���W �0]7�:}Y�N:�3�0� ��9ற�5�k�]��?�IӃP�^���<�@��b��gZ���ADۂ��ZO ��M��$��h������Z��ۘ���Ρ!������� =��T�uj��&���#4�߬<��7�9���W|���Ŗ]��2��<C���î�ғYL).�X�tم� �2⾕�9Q�,�&��ūV�.�,j�{�2�	k�G����9��:�KD����:��I<�?}6�ś�7o���KdjNL����Q�ݩ�k��\�B&�����kp��t��m��%c�-�V� 5��ccc/��Ի�Dg��0u����8��A�%벗ATH�	E�-�'�l)�.��I�K�y�~�+O��#��8�J8p��A6T�ȳ�V֭�xDA�`A��pg3�.
"N���`N�[ʫVUU%NK<���z�����b>!��z95�ͭ�~��*>9�Zt���]�5��R��H����=����z#��`��
2$,<��,����N���1˻�w��N���Sk��{*\�w�ء��PP eh��ŷo�.d���g���yO8�S�T)Po�O���U- 'c]����ܞ��.uq�ҵ_\8�������g��!�Y�I�p�4�'�ɤ?o����Ҍ!�v��J:�^��<5U_��O/ߎ�塁 �^�܏5Sʍ��&�r]7�;�U	&O4H�9�0*9��<C-w4�z����xP乹��D/�Ή8�5�������B��j�Y2?0!�穦�{-���Ua���r��\o	kO�o��Pf��%�H&)��A����,�⩬�����e��R<���(�<�Et���|�qZ�x9m�r�6$���n��"D.���ݳX��ǟ�?V����O��`����-�U��"�wMk3�����-y�v ��]������ѣ�t�����O�B��q
g��tݐ�2�:�L�b+�����S:�L)W���Q5x)A�FE�1�V�9�?�Va#Y�nA�_!��/�1
<�e���;4t$$xc��e�2֚Ӥ[����hV�_���q|dd䖋����*=E+�n(��Wc�??g�Z *�d�+roMq�3[Q,x������8���)����q
r����9�KJ�ĺ�/=�s��V�kj�0��//�TTR�b)����2�����(\Ԭ��y�]f���c�������"9�W��]dqS5?'��ao�^mS�c~³y�������޺��&;҆ī�I�N���VX�z�UI�	|�T�() Ru��,
N�{ MŮ��9m��z�ut���n�VN,{[qcqU��\�³�d�w���*�-ySE;vhG})�&@5�w?�vʕ��C�Fy�R���^�u���*�v�!O�}�8g�*�#n1������jy՗��ni>�:nQRi��4,:,;��r�d?��z���7�(��k�j�+X�M*��t���� x�}��¢�:28!S��}�ú9 �l!��6��]�@���N��y�dւ�j��N�����a�*�V�b����Uu}�i��GF�j�3=�`�� �E��s�q
w��}�zː� �ibU�����E6q��[  5V���lB\dcS:������+UUQ�+*��a�X ��++�.�ml)O�C��;7�m�K��Y��Aaw_ےy��a���@@���8n�A5�l��֟_�A^��?gfb��aR��t�M1ڙ�	J�G[2>�>�9������;ېr��.����{S���8�d�7rRA6��k׾��f���U �/^��t���Tn!ԭ��Ϧe��_�_t\~h�3d��4���y�l�m����.mA�e��%�)
Ҽ6�?­{�ĕg��b���� �g6��^��s� Xѡ���Ï���Hq���-�Ÿ)NA}����gth��2��]���m�9/W_lqjF?��6�ZK����0F����M�\��k�D�tQ\|�	#�����~k�KL=Ft��n3)�̫&j�_KL� q5��Y[t3l� �՞F�k�����+}3N�)��m0�������I֬���V��76����(,=o8/P�{����(ƙeL*̋b�7V������r�w�5�!j*"��E'�Q�q�v׸���c���_��8��^����r��/�/y����~�cΉ#�_<�bժ�
%�d���[H�����~Z[~�����ܿl)띌Fw�">P.Dr9Q�?���>�-�;�<i��L�����A(a�;�r��`M�Ԏ�ԩ�@�7_��[M��)h�b��N�-䶜V���#�My�
�����Q���|�����bU�ng��9M��}n4�!��E���M(4�)i�[s��W��hѢ��οm-��s啊�"����9�6{�Ϻ�0��}�|z'4�F3��^��^=㘂��Ą��w]�H�x���I�/4|^W-i�gv�x	|�ј��6�����)��l��Y4�
g�R� �9��ǝ!a�������<�) _�����������ܡ���|c��K�J���,[<>K�����U㹭� 'M����I�#f�����z�Ӣ] 8��)�\���h�����m�=N�᱾��i+�Mq��D	u;�Ѿ�\!!!a.կmG!���y��}���Ɩ��ْ;��.��Z��~6��'�:����u�����R�vP���c0����MT��9f��(�
��ʆ-�&Ϲ[�N5�?��<����n{)�"*����eE%BD�\"C�21�iC�d��=T���$�N�,c�-1�h�2��yu�����ߟߟ���u^�y��<�y��I�d��Y�߻a�bt�����M�:�4{^�.��J���9�������Xs�1��� Q�}��V�����0m9|�䱮h��ẶHЂ4���wIv�\���\O�*iL��ӈӾO�]���9�w� 8A]����������G�4��fD��x�i�/��nS��#��2�pK�|��H9i_�G$�U[&k�W;g)Q���t�� җ\;���G���{5��]��S۬��?��~Y���oYX>RI�D�[��x�<F��USx���\ԕ���e�ӰJ/�d�XmC^?*�~G�����s �ЙB�=_��*�JN����n�jL���~�"���p��l~E>Sk��Uҷ�֌d���!u��[j�w�0.�/�+���N��= PMiҮ^ell\���P7��'��i���$x j�\l1�+#Ds�z*1�-��Z�<�y
�M��G� �C����fc�
(#�D=:� $�i���iZzzS?hnį|��?�_��ç��F��e�����d8�F�~Z;��#�7$e���Β�T@�ɛf��zE�$M3�f���a!ϟR�J�6###��~�q#�鑝�N#���?�>OG�/ݿ��E�o;��V���0���U{��Ĩ5%Rr��P�����nn}<'�p���ˡ�fdb"�~��B��G�j�~�&����Ã�J;�0�������5�ۄ�����Iv2R�����Ӫ2��i����,;���
�#�3����j?о��)�yH��M9�����l<h�(�	_��>����o矰�7�E���R�o�D��O�~���0�bo��3��.��ܪ�[L���P*�yu��X /��c��^&���B��_&�GFGW���u�:�|%��6a�XX>�\����|���!FJ��O;:S?)S�$u�@�y&����yc�t�?�� l��u����B������w�jN����N	�|�~J1�s(�;b��9Ǥ��S���c*�R��E��H1�/�����Ϸ�7)��x܃��s�-����r���z��X��S>ף�t��կkM�}����Gt"�5�������O���2���mC[ˁ���\t6��7P��^)�7'���>��= ��ƣq@�����8�H;�a>�ݾ{*�Q8����Ko�k}��z�$]�КĪ�K{ !��-���;�sI�`ėm�>h|�vN����%M/�Z��"�o�=Nn�t7������0iu^��I�������Հ)��P���܌��}Rzv���]�0�.u2�6[=�~�<F���9�֌0$�J�"O�ۯ�o��p��\/
IAB-k�[q��%�B�Ӱ�"+T���p��>�4��7�:;M��[]�ӯ[�_F��cդ���׼MƦgg���*+�,v��o2~�7<�B!ctfRbb!\�n�0�+�U�K��a�n�*cR�l%��5�:WJG�^��B�o?�d��GWD��:���N��jc��	�gX�Pt�&��|��[S�$]�����!�Dk���9|�碲r	�w�T�xow��Iy�a����������>����_r��~�vQ.���|�#O���s��\��
(>�i���)��e]����	��Ke�<���	�:��"��J,�OѨCt<�;p�ضg'�v���y�{�n��.聺�1Vn3�D
n���>����1�^q���_��[ ���8p_`��
����.`���:�6hF���/�-@�0|��o���O��W-���Hڂѫ.g3~��P3�8�A���]�Ky^ywݢ+wK�Iy v��J��Cؗ@�q���ͱd!���Q�����M�WPЦ��*��z�F���l�8kw|���0U��Ð=o�����o9z>��u4����N9�W7��D�Zk�^ZxPf�wF'�DH�e��;�x4F����KӋZ~;�=���N�=d�d˥eu�ʸ��,�p� �@0|-�,�eOo93���^0�A��.Ve�;\&[8qbgH��n�'o�����6Ji���9���v�?��˗RSSs��p;��H��H��d����ͼ��s�y�����Y��	L��&��,qKӁ~Y�!�3N���,�I�
��$�#�>��0�G��N��-�ͣ�U�����RVv�}AV���䴧ha�ӆ������'�~�+}��/�#q����<��.���U�G���ȊS)� �m`�2�Y'˗`0�} \g��P6�����4�$�&��q�h��h�Q���	M��o�5F߾�|������X��վ��N�8I5n:�o��o
�q��*q�ϛ0*��ν4�G7��������mAS�i�}��zr.�]������1�G77Q�QY/!t��;������e$�S(�Ӟ�����d:���N-U�x��[ɶ�1Z7ݍ���~Rơ_敖bB@YE��;9k���?W����:���Y�!F�0���R
��"�'0ᦉ�D��#��ڗyy�4�"�ݷ�Vɉ�I�ɦc1�z�b����ݛF�^��֡��� �R�	���n�C��F쐐(�8����z���ͺkb9���羇䋺���S�!�G������3eɥkQ+W,�t|}�\��j�L�v�\�T�\��y�?ȋ������,z�5���s<��44�LԇXLMJѱ��/@迤���}�ZL. |V����z�����`ʮm�� �C���^T��;�������@	.C,�_'�0�sj�Rp��\��؇b�Cѵ�#�#����f��-���_NLSg=&���C�*l��YtH��Q�8�����df���P���\�YY���~v��V�����W}��=���nnh��}�&�PV	��m����Y�w�N���P4A�w^"�,�kچ}�e�L�7q=G���r����g�h��_�n�0����NCض�+���e_
���^Ot�b��q��\���:#������PP&�Rj�H�8�?pQt��g�p�����K�1gO�3�*����Xt���+<!w!�[�4T>]�$�p��3g�8]�7�%
�#RC$P4�%�?��9������?TؠM���u8ŢS/U/U�Uݔ�����5��ϝ�55կ������`x�Fj�fN�n��+�ؿ���� �n���ﴲ�j.�ptԳ��3
����7p�*'���q;����0]��<(�GA��W��K���%&y4;�W�>��t�S���d&@Z��ؙ{^c8L��j���n)�њ��9�5�)`����ܰ���/�u�t{�2D�)焆$tGJ>q��������V��0p���5TAm����O6����g����s%T]�sa�d�AzW$6.�����������@�5\(^8M�oA���.<r�tJ	݆Beu�Y�g��|��>0s����'����CCe�GՅ���h.�v�NM�����)�Jg�k�p���}]������	��X�$�E��iT���'XgD����-�ɰ���WQQ�{��$b�^�`6b
Lu-�vW�t�DQ���100��*+��#S���.�ą����Rv�Y����T����{�T����Յ]EI�3Â�t-�
���Yl��q��0`S�ԩ��^�vb0�V^=��:*#������S[m+�E3>J�7��qc5�XhR|I��g���,�r����F�s�lv�����l5���B������xH%�g��xN��B��R��]���D��'��i�o�Ҧ5�|���Gqn���' � P�z$Y�_�qqqy�j��_���P�M�/=���sGr��b��<o7��Y�Ԅl�����TF���\#�D~��I���_�"*�ՖbƓ�w��M����C��~�ʀ��]iM��;:�*+�C���d�s�ٽ�?ȶ�U�Y]����?n�s:
��������6쑌��+A����"s����B�p�:�(6�ݬ��nz<�(�Q��U,�9__N��ZO�$�j�A����5P�f!���,��N6g��K{֬��n�UX p凞���2x����"�����c��C�;�f}����(��xV^d��O� �_����<��k-��"X�DN%�����(_��@�O��*0��,�t�DW^��y���I=,�l�-��}y{tt����fJ�B
�T�@������
�!Eg�5N�/���Q�Ҷ�8cۑ$׿��a8�W���1��I/�՞&7*�����W��	*N�k�#�ȵ�"h��k��k��D��N ǃ
�1��[���Տ$MgQ(��
U\�S$�.�����e�����o�D��?Q�m���^Tg�e��b�LT__d�kv��VA*��8�׸�ĝ���y
�ыa��?]�C�"�qM�%x�S�Z!PSRR�8?�憃�Y9�c���{��&�1�7���j�g�W�3m|�[P��ȉ#1R-ǒ��Q픦�&�����~c�Y����LizP�"�^YUtV��]^3�^b�M3�!�����#��+�;��e���
㒨�����9�O���l�bN�GG��/��lL��P����a#���j�վ�FN�m�rֽ)�i@���y�5�Jg�/:���e;y�JM�I�##~���_�L�4�H�#��`{��'���#<\fr�6�����Bu��	�w֑�}c{.]w�jW\���>z{�
�~III=��U}�N(�$j
���\�����jc����
Y��`G�+�6ZTɝ�Wl}�>9�� DJ�����M�*Vք̓l3����Ti��G����N��9��as��̛��Α��
����P��F7��ћ��t�����\z1 {�����1�,j��H���|�����:V�0��r��$���ϟ� ���~�>(�"����9��싷�vm�����2�~Or���$�S�z)I����%.M��e��Ӄ�{G,:�-� �1��ռ]��%�R�G+�a�hN�c6�w�8+��CW�Ķ��e#k��53�J;�[183kcgU3=�Y��ڭ}�g׉m_��:��a|�ڴPp�iq|�^�6�z�OT:899891�X����k8�u�_[/���#+��ι�ɺF�i�m��$�\��jY�=�������3Ƭ���}�RE\������j_���<����ˆ�3=�Ś�Ì�I*I�|�lu\�������ۉG���נ�P�V�M�Pg~;s#��۷ĩ�����E߃J�%+)���]�|���]�d������������{C��1.���-'-�Lu۾i�E�|���J47�失��m)�7(�zO:}��|f�l�K��u�xPp�I>vQp�,�c^0�m�g�,�> P=���C�\�-��m�k-ʦ��tE�W�q�F4vV66MN_=�;�	����`�dƛ*Wx�A��*)J�%��m+eXd!ͣ��n�N�� i���I�"]�����[�d��]iBUhO~��QV�7�1����O��}����'��H�,�-��g�R��$�NO�q��T;�]�j��#{F'�h��6�S�tE�S���@ݧX�+��FĽR���J J�s��0֦����F��u޺n���pKx��xJҏX�F%�l�%�P&�Qx��ۧP��U�{Y��{��4
5j$RH�l��ϋ�D��<���"bp"���4	?�oo��#���_�s��������8������_Cp���7
ʇ�����V/���i���U>L�!�}]�|�-�I�Pb��[���~z�3(�H�٠������h��F��@���r�n|X9�Y�Q��&}������I���$��Y��ol��0�����ni���'�h<I�-Kc�}��[kW�?#`eG$,��9��7r{�=��p�~Ǐ�忾�r���>��j��9��R�^�j	���������4iII����-�iԱH�BZQ�ً��O�t�-d&�+ʌh�����_Hg��w(�ZdS%Z~kΫ���&�bqk� -�T|���b!ؙ�]�[�sff�R�!�l�r��]Z���S*����G{��N��Ǣ�׉-�X�...����T-"����������1�������k�I��Sݖ����pp�,��-H�XF"'�lXô �N����h'�K��Q�ߍ�?~�����	w�7n�MY�`��<	XR��j�!w1F0��r�*�-[���Z�Q��&
G���3�]c��$�>��FvC�����v��f"��zi�����A��L4N�av.#�|�~���Ç�x��~�
kHѽ�4"�k*Ll�%c0�̑J��/_�(�`��CC�٤Ǌ�{2�����~���3sW��$�D+*8�!`�F�Y�+j}���Ƈ	6F=�����{���\���<��"������}^�o�_ً�3�M�Swm����<A����R��ꪪ2� �p�	y�]���1}#Gxѻ����T��OM	m���{_;�ɤ[!(�-u����7֨�����Hzƥ;��|d\�y�}�X�f���Ѧ$��R>�[� !��Y�Q\�	��a���M��Nx�M�H�4g�7����n�ϰ�a��G'xmp.����)��jKIF��uD���ԓI֓���7�� 8m$���J�KI1�����J��LoRB�I����@..?����PK���q**����&�q�b�VJ����k�.5XvG9gX��Ɩ����
��l��E���@�M��h�����v�(�o z�mV3��Xof]LLL����F�!�g����r&�5�*���� �lWfgW��M}�ǻ��FC�4}Ksww��	<���
�>s����q ��6~A�@�L�X��v��cI��O?�:�������9y�ǰ��q=w|�S�Ǧ�6�B� �y�>.8�tM�̥'�A|���D���|�yG7�e�J��&����ϷK�G�1G]�/�(�F�cU�s�b�nL�������6>�X�o���'#�)�H�mi)��Wl(����6z����;-yJ@Q������G-�R��NS�1�-�g��~�ڥ��O��FIf���{V,�����J��/%��zۥG�ۮ���{����Çw�7�F^�~�֍p�9�3�F�D@z�RO��������~��X�C����ѣcۻ
�'F�2��Uk1�d�/�^Eʖ�C��3zF]wr��c��5������Vj*����`[����7��FEe�@>|Q'��,�����Tk\n��ƽb1@֩i���#��q)�{���_����@�
��5�|�HE����ݜRO����,�x�G���`�$�ʘ7F�3�R���^�ü��֪�����$#�-]Wt�A�)+ C5�^�-&ֆLD*����@�+P՛q�n�w����D����~W94d[�ڢjMu��n86Y���^�]�?]�΄��o=�0�}V�����̷WԐ#}�)yV����s�!b�������"y�-�3v�}�M�D}��V意y���YGDOP>�L��4m�6�R����������+�H�5�Pz�t�J1�W;�ܹ3��\[��S�,q=����V��j�١���=$ z�����I�%���W�����<'�_�Q�V�g��C��,!u.�۾���Z�D+�3��9c\���� ����@,����y/-�����i���ǐp{ݿթ� �١��z"��_Vtmi����h*�����? �r�!Ah�t1 ���%��!������C��HFd #Y����(w�|��|�C1P�[��&U��qJ�SnD�QV���&;'�Qж���-u����(�^NT����|�|�M�|���5,�EΥo��T�J&�m���Zܱ
?��6yZ"ɇ3�6YF���E����K߄���4��B�]�R��<�S�EB�5��lͶi;p�smDR[}���*ɑwʜF��.bv�ʕP��'IY�r�K=zTW��,��r�*���i>���!�Dj��H���i�O܉�g�T�&7ɋ����~`���ihh��5��^�ύ;!�����]����B'���6����,�y��>>��e|��Ύ�������� `x����?C/~��fPntS���>7��zD��4��a��Pǖ(Cڂuq��
�̅ޱS��RpP�9�rqf.}k��o5'���u��:&&\r���0�q�['C��Z9��֕1.��m��u�a�@ �?xy5�m��Qe\�Ɏ��N�)l��0h����PxIq��o��5$����!+Ev�]�'�_�M%�www;1�H/��UWlO�Y�ϩ�H1ғ@]l��e9\�<l^9���ع	��_a\�E|��n=���١?q7��`��/Fv��`іmmKyy꡸�ۈ&W��Z�=��Ӧ��P�&�Cgg�E���B��δs�?���0ZEZj���97"H-Ο�5��ok�5:�>���?�5��mX�H,�����
���8��B�ﰺ�y��xIEE�]�i��ȹl%�3��K# �0�e�"�bݰκ���n�Q;���3� �U�$�S�N=7ю�waΜ��Y�� ����v�曤WB����ݞ��YRT����A+�����?C���E+��z��.��T�PO������3o�jf1�@ڜg�,H���<!��L;���?��|b58����~�R�bȈ[`:�-^�O/��s`����|Y���B%��7=���a*7�T��v�'M���Pm����X�E΂ȁ�H|@w�ŪTl�72c���#/�vb~~MY�ͪ�jk?a�(V2H������.h,�8��d��?�ȋ5xN�t�W���^������'��OϺ2���L��A~yW�'đ}�>~��3��z����d�71��Z\���c����-�C������3.[V���J9��q��!�`���uc�(�]Q��WPṷSD3*h��eڜf<���jq��
E�R����ӑ�~�����Ր��
����v��g˝���Q~ ��u}��lKqZ�Al���xE���-C!ok_���_��
A@5��?���s	n��!F�[h�y�W���`P>,B��L/����9V�6 �s�^��ζ�3�|�f��`d�B�==�[\����IR�~�]�"��g�i��k�
6dZ���~�Pwh�8�&\��>ho�ˉ�(�!���{P3�'�d�D7v��h��F�$7(�������rnvf��@~��UM���ʐvT"�'�t����i����a��w�����C��2�k������ @�~��*r��5���U(���ar���%�]����,����&�$�_Z �u��`�gQ�Z��Ģeϙ�wt���e�m䗒�p��_�Ȫ�t�sqv��>����s�]���L )S �V�(}jɅ���2�]%<-����if�S��l^c4�s-A;��46D�F�F5�����3A=%�V��b 0>:!Ё�_2߿;�h~��=�1���.W1g�׮|~���Bގt�Q��[�~�N��7�fG��LorJ����<y��Z�V�H#y��&��p8�9S��F�X�q�-~�4���Y;������;�	5v&�g��*���N�������e��'}Wo�h)��x8|�:��ğ�jqO$�N;_���1�CU:����Q$|�����9�� ��=T�¨�J������6F-��4na�Xr�U����lSP5(��.�!8��A���k�~�G%%Gć�Cn��?��mh��ͭJ�A� �2H�c��ƶ�����^^xY��t�׾Z�?��?�����0@��C�ߚHZ�5l +��Bw2����()��<�#g?vc���犔�k����|?�s��+���'ι�}I%	���u�ۺd�?��!�ʣs7�9�R|Y*�-�ٱ79�.FEë�7������xL^���KQ%�.k
s��+f��vD�[$���q�Ug��΄}�4��j�[�b�G�D���5�����`-����T���/͂�w��[e-�E��yg,�N���w�4�� i}[���j+��w� �2���.r��PN��"�"Q��gs��痾\���8��i�IzK~9�c���W��?�"�9�g���#O�55�=���=����-����Ha �$ :��G�]2���?� c2Kю����L:me��@���$v�^�yuռԟݭ
Il���F�:�f^��As����]��㪐�f9/'�WV��"�w<k��lB5	8�}g��%��i[cg�y���b�#=��B@���Y���8�ؕ�O^޽.��>����)Qp���ha2s��ݾ�����!�/��C���Q�m@��&7��Z0���0�#�&m!�?�H:�)�!�^z2�0�e�����ש4�������7�[?�^o��}�¿�K�'�M�y�q�}ci�OY�v���
���x:(P� ��e�G>�
TL2/�%��Ӿ��E$߿�����[��L��Cf��	�,{s�����o�,ܺ�v�P�
��h�}��@!AY��v+����ȑs,UoT����S����c�`���ՒԴ�����@������閿@JZ���]����ӄi��8����ȫ�݁��Yd<�oRZ�J��_�>��G	�q�\@���n�e2��̿�?+'�*j��j�d���$�C�7ڮ�/���u�K[��<����5u,�/_>�و����i�F>�+#]g	�)(ճ?L�O�Z~5A��HA��k�����؎�t���k"3p�h���ge��\��ƹFY|"l����{�79pF��	��?��,�gh6�ni@M��Xi�l��[gju;(��P��Y��eh��܋ �q�"S����a�1Pb��w{Xy�),X�$��.9�ׇ�R\~"����e$��w��3X�yA�K"NU��y�Y
�x��3YU�a�j�*g��xN5��Ν��~�Hb#��"ը��r�"�L/sW��"���~C���?��i��Ov{�鼇�E�	������P{0;3s[�S��u�z-��n.x��j��A���?�V[���Px�^��"��(O�c��EC���
K�����ș�_�% �V� ���}����xrncދ����������|Y��i���i/΍U4f ��@�����UPfN«.b��!��9EC*�f�\I��Dc\���Wuy�q�%B=G��H+�T��V~4*8s	�ѽ=
`��*NN?��K;H��
�<[1�:���h��?q�[~�	Q�dsC�9�Q�'kZ��f.h�T�L�۫�rx�ĺ��D��h�X�5��r�Z&����ļ�`�ҧ��SV�hTH�iI�o�i��;6���]��<���5ʁ
|���J����
��LOYY�ųgkRT�Gcg�M?֤�RN�$*R��n�K>i�(��[ � ���ת��q��{s.�8&�����W;=�U�L<#��#��S�a*P���n�8H5#�B��~�U�7�f��O6.J��,4x��=z��8֔��������vY-��/��Aa���V5��X7o{�겆KY99;�����{W��]u���^縇�g���vR�'V��={�A�m�Ҙ�4����V}��䟕��FZ HO�iw1��C1�QU�k�`Xt�xz��.ϝ&� ���K����������3c�6� �&�*��� }��J���_۽�4p�/ ���&p�����n�@�M�$3nKH<�ӧ��#��c��"����m<��0x*E���Z��ɋ60׿
�������|����c
��Tw>�	ʴ�nn��Z�I^�p#�������4���s�<)lrSC��W d���%��G�h���I�5I��P ϻ ���|=�����o��U�[z�P���҄����A)12@��zג�ݥ�ڳ.��U�#2w��/|��(Ԩ��k����3�������FA1����+�s��𲡡3�F�������8�Hv�^�[���h���;����w��$FH�����ZC#Z�(��:0ڔS�$�ӽ���k�����:��k�;��hlf��u�[T"�j�W�|=���4ע��5K��E����e5;ׯ`��#R��IK���gdB\����d����4��?�&�~��n��Yj	O�I`.��(}4ZM�m�ȼv�?�4�䭉	��.U���Dty&}����;=��V��ju2�A;<�UGc-wh��, {���/R�����+@�~�ǡ�|46�����*�I� DR�T��p�x=B��P��i3�����:�D���~�w�"�Pjg�ͼ㴇����i]�T��&���i��36Z������b�[Zı���hS�='a���1����۬CL��̑�eOU���������ꯍ��ݘ�J�E��A� t����=`oqc�%�:��0/�WZ�Ѻ�E�x���|��]���$��Ny|��RbZ���G0��hB�Ma	��q�̈́4�C-�Wb��%�n�?��r�ͻe���K: 8��O%7K(@_RAAbW4�6�d:\��P���s�,���S)s�%���of�ؾ��=>3&�����E���rl��;a��Y������E��ӟaS�-PC�m�!.6�4�i~z�@�ha��@����ᴜ�+�c,\�P��(�e��ۧ�������
�� �϶�j��N��Ǡk��'���+��V�^��6�=�e϶�V���^V�G��Y���C
~	˦�#\r���S���tQI��u�*��0���	�3�aA��3g���e�����Qg<M#BV���p�k֔���3jl *�.D��Ed����!k�gl"��<|3_�t��^ڑҔ\w��>g�.���V�n�X������#M���{o�"LG=ۂoI��?�@�̛ر�rX3����t@	(o׺EXb_�Uc���B#���[��;�GO���d̵$�_c�R*���(�<�=��U�}��HO�$��Eh���ڤ�E�N��0�#e���ot��}�~����y�W�I_����t��'�+|)�w�7%I.nd#^~�@:�N�����I���֥�ڕ�_l.����V���	�d;/+���r�����*u���-��?���)��j�"�i���'&��&�����޳y+rX�����D��
������<�<��A��3��-��:ǪUl%�S���¬x���g�1�hB�t�7tD��m������dن�M�kW�!�|�><&�Zoq;̆M�����m=���"�~|�4$�;�n��>uk��jn	x!��?e"ǣ��v���W3Ot[�&�<�npQ9,G�?�aGe��ȣ�kYD��z�a�{�����\���I���H�7!w����fy��U�|�������H�k���঑���ԡ�}��x�55�4w��j�AvTk;���pE�#-2���Uc��D�C'%~�����J"�we��dز��-x�t���{B*��e-��CQbn�IjdDOW17b�R�}W�WU݅���h�oGL}����Np|�EGl:��ձ�G�O[:g̶��œK�}V^��@ |l�[� ���`���U���4ՙ���[��ˡ$��F�%P�u(�9;;g�n<����=���ʄl�̾}�۴��w�ލ�_�W���d�1�E~b|�H�MbUډ�M�O����j})�t~L�`���_�$�FU����h����T3}����Q�0�z���������7���R��D��y��@�_�#�k������]��װM�zL[ ��Sz0�SK S嫙���n�}z��l�~�z��}�`���C5~k��z�HXU�Ƶ����֦O ���9*Z��x���U>��}�������U������()��b*�Ǩ���>�U������Z�)~�5'rX!����@����i�O��/P�������T��<e1�0O�(2���� �"B�t������$YK�?+�;��=�DH�bz�^��@E���<;<1��x&V��o l��NM��[��UW�\92=�EE��7��T� Ϧ�j�7Q9���ׯ_�r�����."��t�g�+p�?�C��\�qhi��Z�l)�-s)�"�x�%��rQ�x3������Q89���I�s=DCs�]O���V�˟'޽�m�UT��D������W�=̧�m]t�D�i�"B�5T����T�C���OD��O�v���K�WU�:�"���PJ4f����tdS�3/���?ga��q �/Z/�d�&�g�� !݇�T��+U�{�Ծ�*��7վ�� N���d�>g���7o�
�]�Lv/S�sq�9@P"���*�[4c(��D�'�j�N�"6j]Cug4hu�����@������nl�ڗ������#^V#,a�Bn�h˺��m�aT6�9���_�fQ��c��u�|���P姳�g$G�N�$cI�ӵR���
Ʃ�w}��-5��C�f^&�O�5K�jO�����S�Eօ]w�n�<g�#�;"�NШ�J1k����.	4/�A�X�:š��,�z� ������F.��Tx��F���]��:�"��rQ� �V)���G�_��Rm�J�����Q}�.D��qu4�O-Cmc��E��xMCɪ?���,�#~�������\Y���ׁ���G��d��7�=L���]�-�I���0A'V�}SP��6�\�z�\�&
g�r����_�9�����t��<���M`���v���s�%��Dʷ'g�̞�V��a�im�n�2̀��_8�X?��y�`l�p�NsIwy�jp+�E x0���t���e�
x�G����K{H-&�#yF^���������K�>2�RN�w�K:N�ŋ4v�~y~���Y�����A�y��+;�Rɷ��}��0@�cF���g�B��^�37j�f�
�ь3m߻kfK�C�VV��3���Ӵa6i� Gz+���_FWN�?%9>k�aB�� �� &��r�#��ќd����D-����V�L���c�a��R_NL�j�EDD�W Ȩ}���s�'�غ{���Ǩ�b;>�f��G�dZr&�$�������m��vҶ��;lj��p�X3iJ�}%){2�
�0�μq�'xm|W^��O�!��6���v�O�gg3B��3H���aaj+�}Fk�n�/�b��j��iA\���= ۾�QLt��m&xW��ѣ���
��h}q�gf�YX����YQ�D>�S ��]I�u�\d�/��*�h�-�r���a�TƟG�-��T��V4�Z~Ja��#���9��cdr0Y��i�тf0��:9i�.y|�M�F��f�[L~`�*0������f��0�[�v�� O� \�Ab���v4���`�Ǿ~Y�Q3s$έ�		gN�!7h����Zow���P���	i����HԽ����'O'>h�Y��4r)h${���c=ۛ�k����CW����>{ b�M��@_���QD�su���kW�s�(Y
��$iDSȄt(���ٙa�v�Nև�<�Yd���������ҀJ�K5î��:��#G$?���R�Y&
m��)�Ǒ�U�gZ{���C���X7������ ޤ?疕h�#PK�q�D_xo$��~h(/��F����54*�	�sĠ�/��uA�JjHЬ��8��$�~�K�)féP���o�d�_x<:��AO�u�iWO�5>�;�V��yy�Ojz�@?[��;�6���@�-	��j[�)�]��	W�O#(���h��M�o ŵvs��`�/���\ 
933<k�BkC�tlk58�E�˪6*8z�[��������T	i�sl�r_C$�j{F]���w�[ڱ�"�����Q���� _;��i\x��JD�ד,>��"���ץh7ۊ�Fr*^%����xI�4;r�x�Yb����v=��W��y�ٱٙ��jPo��ͩ��i䚹��V}[Z*>���A�p/��vM�yeZ����m'~��S�gQz9{O믌q!�EO����`t#���N��Q��N�� �uK������~�=pQ/��K��G�Y*_M�Of��L�|�fL{Q�/��U���r�moE0nx!�A�Ͷ�8CtY�,��Х��%��X��Q\�q�#ׯ��;��6�������ZD��I����b�U�얕�d����(��L;���$$�ep�2��9i�˱[@st��Ң=I'��NE`{��y�g�5k�:�2m֝�˙�e��������H��'�:��ɖ�*I�N�cuaEF\''�q̿x�@�J�9��&�"R�IHj�iCxP�o��A�
��=~�a��\,��%�z�^�0���.�r�M�!IT5���nM�75R	��� �0pb�u�F��������`
u�� �G�tf$d���v�̲����#m�l�-����6�޸�P-$��h��1ɘx�u�[��;���4��?����D˟���D�Ъ�����)����m�y z�"����@�*�2�����ck��wuߺ.�H��>���{�g�L=zt�LY>@�jͷ�|G���F��6y��:��g%Zf�~���Y�[m~���RV�׌!=I��΃�ԯX��?Q��Cj�|)-��1c��|	Py2a
��:��T�CA��	|~o�{5��%����r#:.�����T��L�:��+��=�rIp��I�4���9�_9����NVw���=��@LLoeH�|���g>��/��r<AK�V����c\�1��W��Y�ޘ&�H�&��V�N�m��/�0�w#�	@�\F��ڢ�@?�xL.���>��f���s��H.ܺ��fu����\g��ҵ�,ZH���Y|u�tȔAQ�da����#, ��H­`ϥTmJ?�E��~��d�A��#����7�I��"�$h����B����>��[�J�T\Y��Gs��f��l�3�m��*Y��F���VW��ղ�L�m����߅ΗӍ����E<l��ࡀ�i�Y���}���nKck@�m�5���䆻7ڮ��VFZz{qq��$j�~���ϴ$r��~x#�D��mV�4������$`��MO2FBk�߲!�Yx��Lc�a���Xߘ��v[Gj�%�gH�8<��e�q�?y�7��ƛ�_a��/zrv]���e��[�&����ӟl���M��C��S$����*{�Q3]��sS
���S��x��U=N򞹣3�L(��ݾp�=���l�;�'�T��Lo���}�+������=����wF��� 7�������Ƭ��a�3z��)fɝ}���>�� �'Cg�H�P�$E�~|���s���'.��IǾ`�\*����6�|lI�1Y�N�&�H�^��3(�̧��E�%�I_�����L���nD����W��t�ϓ�����~yY�M�@W?H���������q|�D{�߮�����p*,�ȅ��1���}�m��|tF�P��ɱ�ضA�qn����Y�����@A�\�b�kו�P��jՠc��ԩx�=rGc͈������Z�j�nt��}ɓ���{�����PkyktIGr��iw���!=t#��ro"{��hK�T�M��Z��Z�r���K����!&��k���Y�j�B'
����o�����ㄆ���3Z���C>DK�:y�}}}��[:ˀf^ºǷ�ܩM����ؤ���ˤ�H�K�YՔ6���I�U�:���J49��H4ZAJHb|�6XF���:�F��N9�<�蠟�_�2'�ͦO�9ty�wo��K��l�@t���Q��P�����-V��3�x!�c��� U�S��N�1K���b��[f�R����G���m�Y�����Gጿ2ܚHP?o��J;w:�%I���-�R�N�Ҟ?_e&,<<�p��0�p��0h��X�ܯ��uK}�l9�A��|acm����W������*���J������s�V.�0�.�����ڱ^w]Xy�ڹh��`�2��p�;
���QR�Ղ�~�M�m�:�²��u��/�����Lz>3�LA�J��������Bᝮ�[&>pz� ��{����^��0	�]��$:9��ūM����*�߄����l�hnTB�Gj��W��[Go��KXB�,�_h��|>�4����/���P������bN�݀��(���������3������
W�ߔ�~�Pg�ͨ8;Q{�ť������ɩ?������AF� ��A�x)�o�uLL���<��[�7<���|�#_J�`x��W��.~��q��?�Ƙr_�a���=��6�9Ռ�_݋��>W�`K��5�P��@�%h��:7��X �9�~"�d�-��ƪM��-�s>۩W]ֹu�,<=;�f����S���y:3����9cI|Rpl����V�B�][ ��T�K�h$w�ɮ�+��(�9�#q���NS��ʘ��xu����A�ml#}�z���ɪ:j�M����ipn�i��{��9dm�8�0u�z�������wPv�����?\m>/Ճί*N*���⫝�w!`ѫ��w.���*�CHq��K�ō�AK���̝�Q��KJ@_,Dg�����M"����DH*��?��@x@��6��$��MY�*�rޤ�\��aWW�I������]��x�~�;np�G�^�W�3�O�cC�PFmR�S����'��ҿ~%���
�����/��w9����� k����m�^XEPQ��,�0�d��l!�̰i�UT��f�%�d��"2#�	�%#a���@�O?�����ӧO��}�{�k�{�}3���"߿4�nڛ�ڼ6B��՛=�e�����氶m���*��ϕ�F�Xǜ�Ҟ���5�65������Q���hyi��������������AD�U�ي�3�.�"�n��tGȈo?�����S�N>k�P���lo8j�'l�e����s��W?d{Oᖑäķ<�k>-�C����^��W_���?��n�G��8؝��M1�+��A�w���.������� Y�k�=rl�>w$��1�`�i�T\};ޠ�����c�m�H�$+O� =.)됭���P1	�J�d=�A~�]�j���z��6<wg�W�t���s9n}{��R���z�{���f��iq�9�U�!jd���=pU%��_�zzX��+?�O����n0��
�k����5?M��f2hG:g����QCT��UO5Sy+D�t�Lg�Iu�qX���X��sE���[^���	�b�������/��F��{;��Y�Y�+�pu�2�q�I���z�­����	T���RP%�>W�&Oy�� j�☀XJ������
�^�+���2\cC**4��ʸ71Eme��������ު��w����v>��2+R3K��yo�sh�>�(��>%��J�e۷J��Q2+71ڂ���e������"�wD���i��7�n:�t#q!j�����/ǁ*���/�����Y�����'&=�]=vYJ\kN�¡���"k^��%&�B<��U@ȅ��Ax��;�:��v*��\���~=)5]]��ƶr�PI���Ԃʂ *�ѹ��)��$P^�4�8�V�p�BS�9���A(>{T�4PE������Dg�9.���%�a��A��5r��F�/�Eh��l��։r��W<O�m͵Az�կ?o*�N�<l{��KI0�@%(�]l�uBK0I�tv�t7 ��i���2�>Ƶ%󆡩3#.��ds�1�kL.�R59)����K���	��UO��n�S������I�A"['R)#$u�n���{���2���
g�������y�m}1H#ʄ��\j{����C8dȔ��4�;M�ߙtN�yj(�]1���mn 5��c���*��Ƕh�Z�O���S FQ�%7�I]����#���#a�. g�%~��r�ϓ�CQis�ߢ���M��J��,>s[#e\������h��F$Y76O�l���T#:裕��.���RO��I��Ѿ�-9�Xx��3<*�S�_�i帏���f8�	����ϕ�Ɏ㳾���-�Q	
�B;7�X!�Ikxj�C!�t���S�L��R*�[C��w��'?��v2�Z}G�3��ZKJ�熊�o�G������f�g�288��-1�8�t��]]��C���c���se"u�`H����T�?��Z��_���8j�הi!�j6G��������\�tA]V.��:��̳hVj��ԱP.>����TZ&�*T��?��+((���>f�ľ�b�K�=�N���^��WS�����/B�?02ֻn�
y�!tuA*�<�V�#���G��ݎ(�R'\| �#�4������[�j"��r�)���ڑ�+W�k�	�����z��8����`�l5����Pǂ�mv]]"��un�V�Zv15�7�\A���ua_�r�ښ�2t�5m+:ٳf����~-@��
��OYE�X��%����<��^Ӑ���H���o�^�iB�HG���Z�s���E�5�!2�$�l���HL����&&`��(�1�ݫ?��CU�ta����չ�rB�����v^Ea���$_�ż�Ǒ�+����(�c���3ʱẾ�w�Y�y�{s��<���Mjz8d�Q�	X9{ ϓ�J�v<�.mp���c���|x���~বS�جl\ `�q�I��^$�˕�;Kcw8�E+z��/t�U,X�`k����4��+��>�7�#�f"�2\�qj#�}x�S�2���&���"n�cmo��_��/��$�^�"��WR���}�UY�Xn�c2PQ�'t��J_�.\�+�����c�	��2�Q�$@Z��˴}G���W��7{�7$9�負�`c�ٛ�2���� ���ٗ��S�t�N5�X��|d^���w��@N���?pL�m��u�����8������W�����r���OQ֑mۘ��%�D�;�6FՔ��GξLB]�����_o��#~[��%����kWWSc�N`U�(��~͚͓��#��U��=$N�ޚ��t�ϴ&B�I~e�ʒW!=�ʮ(��
^,���]}3�0�m�~�;��� Q��+��H�ڋO�	�~�SD�aU�樂�WY�P�#�u�r�G�f���F������^�ۺ���9�fЭ�.�ȷ��B��J�СCH��'�3�>�O���^>�o�ɳ�l8����]F���|+��������=3H��|yЩ���^��A�d�
عv߉��6��(�ׄM�nL�� ��(H|�.�_,����.��Y�����}�S�e�oG�e�]%w�nn�}cp�����X*9����n�_����Ss�Hӡ B��Eo&�]�YВm�#�a��?PqY��E�C=�������ns�~(�Yh��@wbW�\Y9�9�:�Y�}�Oo���T�,���(�G���mgg�B�;`��!-���:j�2���+��QGo�ȯ������(��☗�O��ixQ����p�Ko��Ԍ"M�H�ӂ�<1�^���(a�=�[)�G�0^�	Ȃ��ti�>� �u,��LV�kJ� ����ak���{?ݯ�m��7mfdj���S]ʄꄍ-�g��i�0;B�E,���y����t�f�]���l�����/T��?S�W����5��� �E��777W�h�s�tN�g�<���G������4>5f��Ѱ�H�y�t���1L�C�$�=�$b��#�cvHl)�k8�n��U�-���cOͺ�U�.�ƭ%~�8A��;�716ִ�I�Qq�xk{;.�vC�7�LQ����?5����و�S���mXSVv�;�56"�q�I��|�>��J�;�P4��hL/��-��@lH���q[p�����Tf5Z��SA�����],�0u|q~���.�����Zۦ�� �mD�c9*��("XjqN->�w-�����k������W��:����L׷V���=�-�� ?�(�����.z":����F'A�����cee��	�f3!�8�g^1�l��̫2��Ϗ�Hk�W
B��ȥg«J�7r1@��7���󟉋Rpפ���Y��k�xD�.׼�>u*��/���1Ѱ�Y�+]��o�J�G��s�/���uz��3�u���r���!���ǵ�k��K{��r���mP�;�(�]ASo������t�5A�96}�,#y(Y"�V�7�:�0#�����AM��H�x�����<�o�lC{}^��Z�ͲZZZ.H�����:�P��vN�=���H�I��D�
�qx�`�x:;~?���W4�[~` ���}aA=ڱ�]>E���g��������4��~�Rq�t�C�yp�a��?�Oç��V���f>w�g�7u]�Z�~z��ȏ��P<���{���͠)�D�$rŲ�-Sӳ����[�2j�5ǥ�z/zD�'��h/��񔿆���+�M�}[�����!?]��(��F����/^�|�c�?���1��ǃ�� �ܽ�8غ���	)���W��-,���N��hE�\�X���t{j�ۻ��O�/,#�gR�,fr��Σ��4s�1¯ԋ�OS/�*'�ρ~�R	0����Y��@���`~j�O��3�L��@�;���T����S?�@��_����CK|>���B���ǒK���^���Ӧ��N<��ZOK�n\HW�-JJ�R&���v���`�t�>}���OF�n�x�G��m"��\�F7���mY�f�?��M�iҙ��YW����ۗ�������mw)��{��H�2��x���]�&=�5�ѣ��B;7�ƫ�,����uɱ�/�d%pa)��?��	����.�g�����UJ�$
�b��xVZZ:"&�9���qz�%��/_Δ]�M!��}�騜\25�i�lk���������Gz�D*��x��Z)��%T�X��6���>�c].����I�RH�GBh��7��G	c���4�l$�h�w�M=���M֥�7o���	Yo�4w����d__��@r,���d�kd��bWi�Z��(;�X�*�Վa0��ޚ�Z���!h�Bӳ��&ߛ�d���W�0���iR8���v����-v�(N9r1��g/U�.�f�����B��S�M�J�+��{�+��>P�OA
y^��+�M1�V{Wh�Z��۹qh�7�$z)�}qUbd���¾�xNS�x������,��ﱶ����?��M�.�����w�=o����I$�ْ�"/��III��56a�O��г�a�-xrB�.jK�,��)o�0���^#0N��U;�	�jr���{v�-(�ZױrJ$��t�����E��իǟ7�E�,n�u�M�)��i���x�	m#Qr���aͼ��˳�g��s���RL%R�	��k�C�G2�
km}zi&h�9� ��\1?�ڼ�nƪ���'�0M��h�a�'o���x�p�MN����+L]��,����������j��ˢ�5� ��tb���w��m/?�tt�ґ���'Z���B�/Lt�'��a�R��腻���d����/���0�ai  QRr򆹧������VVo�|Q��;��=�>�QKr 4��[��W͊G]L�$87�`/���>�
���[�˧�W��,��Ez��S�&���)�Py2T5�n8D����S,ehnj�ȃ����=O/%�O�o*����[�:�u� ��د��Co� �F���־��I�4����(��^w�#:T����!�yy��^O��s��\�H$��ǭ����ohh�[R��Y�h���8:f�~��k�ȉu3�66�`�ubB�'�/�e��;]x��L��"Ж���W_�
�Rh��W�:�A�\��d#�w[����v�8�D��L�U�RLR������́�U��b�l[s��͛��qU�w�
O���=�H�0-�j(�y�*y�����߯�]�7�Of	���P�Cw�dLV^ŷ[G����ȉ�O���6N��4y�1Q�N�+�r���ɱ�.�'��sCs5N�ݯS�o`--U��&�R��C�Q�����?Fc�g����v�V�Ap�լD�+��a�e��r����Q�����PI�u�E��SO���ݛ���Ѷ�GꙠ�n�=����rI�SFEEe��t��pojk����6��G)/�����,�wN!�i�i�-1��D�p��>����Y��0[�����m��L2�!��c�� �5*::�Ɍ}��?���Ȣդ�j�63��Oڢw޻�*�8KY��h�G�@�����Ez�bM�<��C!_@�7"Mu���5���ݻ;h&uutt*Î�����u�����V�y;5�a�<�H���^j�s����vz�䋂�n	t<��j&bN��a����3���'��F�����>wԍY�}8�L&�I����puk�K���i,N�N��)��Y?�5/m���7gZ4�V��+����Y��Љq*�����Z�K	�-�?��N�[�������Yf��R��ƴ���o��}$ā�[�=�����ѝ009k����Q�=��?	Z�K�S�^����t��6#{_ U��+w�(��XK��h���&�珶����Ex9�QϺ���C=\���Vt#?����C"�!��C�<�8.�s�ojN��&q��K.��F�D87��n��;�YZ�L��%yW����Y�n��h��0O�t[Z�st߰cs```�K�}	���S������
�uww�$^e5�?I-cYZ�B�ײ�"ZP?�zyG��t�]�"}̪���#bZ�|sZ�W�3����Ix�]�<N�qh׀�[����S��FFu���%,���D�\�:1m��Q���6�]{��(���$d��gj&^9���Z�j�A��a��e`�ls��߫;�����	,�,:K�ok�m��x:~�_��8�\�����DoSz�#R�aQ�!���n�3�i��=�vց�w��mV������B��U��A��H�'gw�!��t:���b͌��u�VH�0O�l�au��&�_K��d$$p�Ѕ���z���e�۷oG(��A��O�Z�*�աa69�M�Sxш����A#%���{49��&��p	��`E��*���������7�/A��C�?q�r��sr�)^�5�m��گ��=��W&e���D|��!J��ݮ�ql�>��3�B�0����<����h������ĄG����!H{���I��t(�Hx]�m��"">�	|~���[ʸId��E�GG?|��Qά�lG�B���F�Kan�e���M�g� ;�}��",��$z$���>N��3L�c\�����ܼT���gų}�s��tT��!F�mx�"1??�%�Si��׿u���C/�@��یfL�>�Sh$���8�H���0R�y)�3$W��.�� ����z�����ͺO5�g�T\�8����������.��6��~rn�!]"##�a�݇��;�>EK��:�^=�d	��\��#H�>
�ޥ��w6;��79G��z�'ƕ�"��h�Y�*��쎸��֚3��iB�T�烵�~i~�9)'?��E��F�#�#k~ġY/�Eg�%&�6����ΙgH${��֬=�T���6��0xԙ?z�^�B���3�XSAG�����{Td]wp�&Qp7���k�ж��zM:��^zw��fE98�1�wn�����_p�ȁT�E�`�3XC�� =;�j�N�M�>�1:K3a�m]]]��v��*gn���1Q���xs����@jNnn���k�ڂ�C���"4؂P���7|v��d�Fg\�HU�_��}	��u�U��q�@-�VF�<����tꉸ?�j=�-���s*܌n���56^H��@Fpz��9^=(7/�f`����{׀Q�����e�t0�x�b�m����hg��;�@�V���M4{��n� �j��ex�^ɡ�8>e
z�ς�)��0���Fe��y�[FTh!,~QW�f�[��m�逥���h(��׍5�nV�oVc�?444��.�$�
��ȼ�⚓��z+�/aZ����(+����m�WWW�:�KҠ�ޘ�;�@{v�-T��H�!�*�p�I���xo�l�:;�(aml��H�i�E���S�?��'YE	s܃�zЏw����,p�+z��׬Kö?1k�1 �8T�������?�.�mq��Ilm�y�}S��Ŵ�Dx�L
�f�:o��ă��c��P���!�u�����4	z�����%m��r.���d�MM��Ə�8}���
.��u襡ѫa��+�67�^t��hrOOO��~hk�`NO���u�P�z]|�iH�3�孥��/G�ـL.
�v'��ϱ������,�+�!�@���>VO�m��w�_|b�J9b�
!z$%K�M�C'��F
[�RU�Om���f`m������G����/�E��:��=F���Ԕ����5��7��,m�xil�50�UUU�������ߝ�v����5��h�@���!�t��)u����0!]�mN~DZ��Li�D�%�M� ��pl߶�;���"�;P����@�W$[���� �����λ*�׬�M����w������ݻw�cwl,=�W��;�^�&�l������ �[�"�/���3�¨������u�F��L����!H��L�Բn��n����mAX5������j�t�kNkr\�%s��\����F��\�mMssEM��D29�&g`B��U69����$�H.��j	��W����]�T�9">����w����݉�*���ޅ��n))#�����e+�&5:���uxT���wvu��Du�b�c�SRD�
��>n�&�CLOG���P3����ϋ��)���ʻ����B��3c��h��X����.a	#�FQ܎�T|����K�9���5D60~�YV���h1b;G�ߌ�@-�ȵ���l�R+{6~*'�A���9�X ׶��70�yx|a�+@X���?~��� �e���X��^�#F�zeW�4?��n�K%��}�HAUr��j�_N��3[�/���h��rUj��YR�@4�7ǁ-.)�z0�a7H�J>�݁M�{�C���Ϝ₼�O�,���)�#;98�ZՔ7�����(kf��y�됋�a`$��� g�GFG�'tJ�?�� ����WI琍�ZN��0��>兘{�����a�=��txk�÷uv�̷��Ō\����Q����Vo�œI��̓i�,��:Vw�����B�
EE<�B��
D�|��H�Քݫq�ŏ��;9���ZIA@�_�� '����<�������iI^�(��g�]
b�$.���M�&s��aگ��'%4qn�P���okk����[��S��=70R���#��f�7�M��J���WAF�0Lm��pI��QMTDD6�&Ӳ���5��_�y���Gڢ�MU��5���㛍_�=F~{�&)��� B��MM}�f�%�c;�KJK3��7>>>x����Њ�2L����r��	?�IޕW��*t��� 9�3��s�E������M����N���@�G[z����\$��΋�κ��������͸�-�:�Y���u/����u쏊� =���°�ō��Kb���ܛ�������l�v
�C����.��N��`�ag����TQ�b��f߽y�����k2i������J�C����?����OD��{7}g"*$�[�^U�/bE1��r&a@d|�/�+��ۤ�������V�0�/���r����^����oߞ<p��Ҵn֥P� 2u��^�z�ݚ�R�.�����Ě
*�a����@n�Oo֥ ���p6�<�}|�c�c6����L��E�bk=��듔��xm#[��?��W5>֊�;��R>�� 6�fxE4��E��H���v�.�j��@�����h���e��{�]
�U�4o�����q ���3|���khu)��n��C����<�db(Me��4����H�fyg����&�AOnFo�'�_$M��_�xdy1挳
цY�r��<߹�mj�3��Dkjjr��.R�������Qy�<�?�f��
�����R4��Ljϒ��_�/0�a��3~�w.AO����� E0P��76����n��)�PZ�,�g���1�,{68U�X��q���+]�W�����e��k��2Ll�)�]U�l��G9�R��pY��4[�=���v��?P.U}T�r}VC�-��,�}ҒAG�� 	�f,�����gǔ7��f�����k�~������tp��C��Ǔsd>�@�1�Yݟ�Ÿ�����(=�'�����&,3@P��K��N�p����U�.h\s�� �u��*��k�����%Ju�D�4�I�<q�:���	�60.���BhD�w�D<̹a��JL�^�pH�V{��-K<d���GnA��Ả"��;���G�tQ�������q������s�8�|XCS	ʶ���m�A�^��PE��1ī q���(�H(����xג�j��W�M���S�][ŝ>��۾�iW��\��A�oV��#�!w!T�\��q ����^��ޡ��^1�9��
_��=Q/%�x}����X;��)#Lٕ��K��Nw���?�#�J*���~�|�0�<�9���{��>{#��<|
R��q�Y����|�kzǦ6�_�� )Dc�#������I���_�7�?�(�-G7���?#���MWƱF``av�����F� �����\ɺvLz�=��*#�V*��r��i�	<i#��i��`T}��]=�5M��}4ePhj���~2��(;c3�F0�2ӱ?��A�Bti�dH������tDJԺ�$�"���诜j�a�`���La���,��Cx��r�kI��M%��i����	���B'��l�+`�����8C�����s|y*��IL���G>����0����x�ܹF4ӖZ�3��i��rQ)��b�u�$���Joٕ_vaM&�\P�΋��nׯ_V���BH���k�m-�O�\�a�+)�@J�ă��ۖ-��\3ҵ5�Jb����J-a��H�%��S���Ң+{�?��L���L� ����u�(Ȳ����ؾ̨R�
�1U�TVc�n�ԗ����������{�%�F��T%�cB��&���_|,T�Fu&c~U��ʨ���Kɢ�����mT���$Y=&T\5Hm|���@`�Z�y=��|�����`�C��:k�$�	h糃�ӄ.�f��X�ب�;u2HlE	>(�,,�l�[4���>O{j���tSh���7�eb�ߌ�͍o[#g ���<Py��s9������kL3��w ������c��q�q�)]*����}����I2L��P�P��jѡ�WZ6�Fsb;�)��;~�L|�U��ۦ�9g� ڕ<c�Q�3�q5�4�\�t�S�/ݲ^iyd�Ǒ���޴+��`qYfVs��<|�@Nl-����`�<!H�_�n�)c�J��#�4�K^4����)�v�*����k��M��֚n6�μ����II:�J�+Ј�4B��P��..W����RӤ?���m����Uk�� IڴO�Z�'Y��Q@.����@�0:Y#�����l�S���ݯ<�
2'g{AK�X�|f*��RXRkjy�:��C�d[�o����_�{R�W��Q9ӱ��}�O?K޿}�(ao�I���Q�F��xz�YOW��ڏ��DV�� <l���j�7���>o(pb���݆A��zyAn�dy�=�������������	��~��7��q��������djƃ�SB�4G�.;]��C���9���������׹k�������Z�֧��\����3j-�R�̾���!`?�� ��Ԭ�փ�g���#��KY�%d�^�sм�^&��غK�l��t�VZ��G�ciY;;����[�?I�`\1�򺎇$ëpD�w**����`��!Ю��:Q�����?,%fJ�-Ƿ�k��[�$ja�(i[���p�؝x�g�(�#!z�7�l:�m������Rߘ�?����"���5OmD{a�Q��<r��
�����
��H�FM�SE��z�J$��3����,�܀v<���d��D�4�.�B���b�ĉ��VR��������^�1N��y*:��մ�4Hc��Y)� ��)TX��������SGCS�Ј���3�1p�ҹ)�ݝь�t5H"��-hJOt9]��˷�鄛�<1��NMz��S���o��Ib����ϏXǱ٘��`)�TF��3� ����1�Bʹ#јŞ��N�M3̬a��W��͡}4R��+~��$�m��Rh�$K9�o��8���":jQ����՛�ֆ�q��ic�	m�vu�F�#���$�� �p�t�tt��)��Dʺ����Z�����
���������J#o��z�	��W�Q@��=77�g��O;SX�u��;s���"�/L$�L�sѢ˶J�j��&��0OJ����:��0��[��;�y��{�ʔ���@��p���$	�KJ=���ݾ��[��y�H5�$	'C;	V1� ;&�ҿ;�,�Q]��%c�X��؈��^z1�Ϣ#��j�pn�`)U�̜v.�&}����<���J�W\+ExZms90����i��	`����Aփ��t~�`g��L|�E�4����Bdd����d��%|-���������vrÆ0誎���j���V��B�����O�:�c䈺m:t�}T��x��I��&����SG�rN�y�C�G��2�nI��wT�B!�T��^<���7zi����1:ȩ��򔯑t�p�/�A*�R�I�&&��^�/��v�(���C�n?����>j�ϥC�:� ��5@Rݘ[�a�8�}1Oڢ	�jY�F�X������!������\�K���L������_f��zN�.i-����̼ �Ǚbʙ�h�s�F
k����ˇ��J��}$��L���@"\�U�>1�Q�up�I7�{�u�}��\�M·w3w��ןh%~&���<0Q���c'�Ν#�� 
;#�@\3����ÍT�I�#:���þ�7<$�N�U\���|~$����w��2���}x��ݹ��}�{ɳ}���V�1JA[����jQ�@��C�c8 ZH񘫔�j��l�1n���J�oo��2s�� �|q%N@�͜�	�-!��N-���j-�yd� ��V��- ��k�u�ʶ��+����Q@j��W��O��i�y�R2a���Ul��`��#����6*��siO���������H�<��J�*!���~����v��fS؃� �|��_ĩ%b�vl�ǰEﭸ�Z)~�!�g>�D�J�`��� E�p������ds9�7rb����̘y�s��h�s�0Xu�U�vtA[-�w���:m�k�L�S�0�()+b���؜~ä��	�N���z��r:�n�O��ÛJ���7�g����;�s��ՍD�](*����'K����(
��0�y��U9�b�$Ā�&`�@Q>w�.
`��C�~����i1~�=�"�I3�S!�2<2bRZ��yyFcaF˳��!DeWx�F��<�$�5幑���Ⱥd�4�l��j����Tm��ԢG��W�����;>��h�]HLL�����kum�7�l����$���5G�ZoTd�J���3�U�ǒ�	��ml�6������+(<�ė��������~�1�L噃�V��6����Es/�`r�����jk	u�U�O�*��r֮7|V�/z%zx�;&��!D�����,O����rh�!['��#$�#9��KpĶ|*��E8N%�}�N�p���3GZѱl/�?@�C�r��+�A]z;��kN�B����o���B�zE�
廅5o�sms�揪ᳬZ�/�r[W;^����-o��`�ZuW}�~5/>��jFM�Q�p��S��1����R�h���'_��Mٱ�[��VQt�c	��kǦP�,8�Ef~�C{�UN��F�C,�y��g$q{=H�d��n6��f�b	��u�����E�61�V�ވr�ZL�ёG�+MT������~�A����C4v�	ʰ�c��{�t��6]-�aa�8)9Y�P_c�DN"������.{JKK�}�R3�p�����倀ιi0&�66�ء�c-��#P�$'L�Z��3y������^(�w|uL5=.�tH�%�Qf�t�0�Ęy������z+w#U��q���k�Z�\���b_ޏ���@�Y�鏠�#j��`i�׍�������TBe��{�m�<�<L_�m
돲=R+��KLݻjU��
+"k���?�����t�'0�ٚ��̕Rw���hק���~9��y�ߩ�(x�jOŌ�R�Fs0)ŝ�ͩ���f��/PA��.�4��;P3��`���v����8m"����&�����]1ݶ��Z
	U��n�u	88���M��ѳ�$��H��	HT�~s�lIv�oUAGG���KR��S� �r=��S��d���Vl�H�� 7��1�Y�lkp���	��5}�J�)�ó3��^�.�ğ/��V9��FY���B�a0��@�ݳ\¸�!��׹��6������Og�4�X�P���E^����ի
F{a�D?%ȗ�d��{��}��$Z��!�
ؐ3�n�]����;�C���4ix��ٍw\�� �k� �>�Zi����1 �e��-�8���@����+r٧9�Bzu\]h���Ō�����q��̶�o��H6��\�_��;%��	�m��O��Q�E����V����n��Q잛+�?4��`>B�6�*�X��_��&�"w�W@IYYY5e��26_��� ��..�_C�<�`����Y5w����co�G�m�G��M���-�J̐1�3N/]3���
�;�%3�+��o�07m"j�76K�#�a�;�	/Vӧ/I�0��������]�lm��}�6�0G��.��wBU�dP������}�X|)Ϸ��0+J��3R>>>�j��1�H&�+�������-�9U��7P����Gw�)����{�x`4ǻi�.m����	���O�=�]�چ��8`��c�T{y�2�����Lue��!	���O��.6����DE97�Š�e^7:2R_Q9��ԽVSa���ĉ�S���@�<�~�Æ�� M[04F��hk�b��h&�Yρa���K�M�4�H���҅^�C��V��er�~n�-G�O�����m--{f�u��2��
�ύ���_]u�9T/ZUo=�n��J��!���r��������#�T"G�p���+J�^�GQ�O�H6LMD�.�U%��j�:�����zVK��WS�Y<E���q�,l�ހ��j����+4@ߗ?��Η��i�H=��7�m˅�B��Fּ�$VT9�Ԉ��E=��W ڃ�O��iz6���Y:R�Z�ڃ��[���i�,�^�h��sp �(U����_����قu�J2=��w�_��eI[v�K4!�-�^6<�Z�'��\�������%K"�{��Ka���cu�?.�u���Ů��n{NSe��z6ُ�i/K,)aT��&�F�M	`@�YZ�A�|�̟�K��p��K-<YJ������P��9R�P.��\��5f,�[c�|�T$g�D�
�u,��3<Y>�]�Z}�1vm����@(��]m�V|���^��5���Z�/֗+��A]g�Lf
��&�ԍMM'�W+r��cY�X�A���&&&1�ڻ81L�R�2��(����i-��sѤG��ho6Ȯ�7dW��}�˪PVJ�v�-����r.�� �ҰB�R�$��L��B;7�1[�
N�U�u��폵��n˗�d�*��vڕ]��fX�A �	���X9�|�eI�D�Hv�˲Y��ve���U�'؝��Q��T��&0%%zk3zѸ��,:ޕ��A��΢g���WM�ʀ�N(D7Q��Ҩ����9$Lg�Oz�=�-�Y�}���i��&M����b	"U�[��/b[��D��19P�@->�LÑh�Q������m�~eߙ����=����[N�=�h���S��V��������;�ߘ?(H|�II���ˮ=G�cF�k���,W~�J�:4� �h��B�9��g0��k,ޝo�M+�F�^���Rw����ˆU1�.���DJ�K��[�v�zWkw`��K�F��%�W��� R��O�������������<�<B�/�RJjSS�\��w�:��^M�?��Ρx��L�ֵ���)�$�� �17?��h�͛W��bg�o���VR�r
��mo�_U�l;�b\�VWn�q��ܪ��\Y_�kbR\1��#���A��/���juL��[��m_ծ�)��~L�H/�&'ejj*�l����K� (%ED7�}6u��k?���c>&�}�
tvl��g���O�%+��`�?��F ���wgHy��S��.��8�qQ�R	��C��W�����QS��8�^� ��^7;���A���u��=��%o�����4�g�@Q�Q`r	�������+Y3�Aw�`=���3(���:��W�rC��=�CQ�r�g� uuu��Ґ���@�R$��L��cݴ�Bd|#��W����h�<n$��k�մ>���ӍCSY"D�i���Rո��#-��?�jI�7�f"v�4�l���0[[Gs~O�-��۰�-X�B��epp��:�k�ѭ��ʙh� ��!��@bvGU0��s�4��d�D�Y���eW��wo���r #=1�]n��������6�
�NR����>���IH7�A���kG�!8'6�8;��M�=�_�n�y�T���h(����7������sf���U��_|Յ��n� ���k^#�u�x�[��	� l��8�4�3GhtC�� �d���m��$«%K>�[�TH�����*Ԉ��w���Q;��ZI�uE]�}W[�%Nv����e�n����}��Z�o��FB���&�ǔ��z)��ࣼhR$?���"^e�k%<c����s)�]��WFu�����d��p,eޏS�#X�P���D�FP8�ي�z��czـ���٦�\;��֤��\"�����^Rd�*�E&�G�;��-\�H;���C����A&Zu�	�3�r��'���H���/��>nMt�ީc3�8"�� T3�|N����>���+-��̧�s�Ks����}r���H|��O��|u}�����D ���q�\"��u��P��\��J���F�uxI�+)�T{j�	M���eߘ a�ħv&_k�U�����R���.ک2�H�y�
����
F��¢��!<O����`<�;|t���o,�U��bk���@�($�=(y�_����ID2sȝ2������2�kkNq��w���x�u|ka|V��ߴ�.
�O�
V��`��Fgkl��޽�<�?�J�d3i�C��yt$凱��u���T09H���4�N+���:/���?"����p�����>�V\���@�������ؿ��B����Ht,w&��C��Ӱ�"D�Oh�\�6d#/�N3�4�+�'���$1Cj��OYӝC �N�R�}�N��g�R3K �V��Y�:u�u}^�4�8�K�XB�)�b/�U���3vn�:�'��<�$�����!v�Z�KNW�-_u���hgQ"����.�F���1ÀP ��x�>�rߍ���x��ۙ�8]�7��n%�.�#f�N��u�F�ѱ��oO"z瑞.�k��>h��K��מ���b�˯�(�Co��[﹪H_�S��G�3&�H��8:�����.��{�:P^F���ba�6l@�8>>�ao:��joXʢ;�ω������ԋ�����z�i�,c��:��G"k�� ����U�b}mot�d�7���(�c�&"!���<�z��qĈ��/��索�A��޵)�.�~~fn�999RE�?�P��fU�.���>���9|�:v��r�4�YSss�\�4���hc�*tnd��9{��D
tQ����/�P���os�ꃵQ����ڸ�}ҋ���_�g�-l� ̂�K����{Q����o��T�+�[���,�\��\��w/��"+�#P68����~s��x��,u�����4�^Dc*s-�b.��'ˣ*��c���@�u~�*�]���c��J&�6Z��܏�����L��w�l&����u�tg�D�K�����bݓ����i ��3��m>�uI��pI��]��#ll�Ңϱ}��<�=<-�g�^y������%�������!!S�f(Bj�FFꋆ���Yk�����zl���LL\�$�U�u�N����\W��n������$Y�׮����C��������6z���'�����i���dsP��,% #1�p)����C�4���h��J����Đߦ
$֣�ߕ���#��p$�s/ڕ�޿��c���?J@ߨ��A��D�k><H��nm"����F�C���K��Awn����qE�T���n��)?�aq�Q)���ח����5@��cJ-���������V�͖��^N)�������U��J��eH���#�.��Hm�w0���
�H�-��'�F6FP����=�ϓ��𢏌�x�h���;�����|ϧ;I�q��,���P����=�үn�@����]��>k�X� ��>	)	l��,۸��$N�.��Ѥ�^�O���Z��x,���p|���B����Q�	m����B����2{�������'<|��pH�+��S�L���i�7��ơ�׬KՀ����8??��N*O╬��ʺ���Zѐ��f�=�܍k`��Mdv|��j�E
����H��!BmQ@@oW�BSCE^9o$���vM����.M�BbQ��a, �����6@UË���Au���A%tL_}�Ԃǜ�Bzk��.��w�q��~�ZY=��j`������}���.�x5�k�񨦴�jF��E�X�	�Qޠ#�g�G@Ф0����I��N)���������/�͡���+	����QK��3}�:�:��
c���Sb�� ��'+U��TE�.�
�3[�_K�ЦFa��φ�����oJ��J�������.\.����ɚ'c̗x�0_�[�V#+]+5���o��/�+s��@ЕD��e��	����x���k@�8�#A��&��Ě~�<��G�QQɔ,]�c�]��W{��ٕ�L���d�0���1m��ů�&mˮ��� �_���_S��J�+P��t����Ԃ��ߚ��3�WJ�[?3����Վ))������<�T�6<�y&j*��O��-��'UX,�T_��;�2��p��m�H�dnaa�K�0�5"1Q3���p|���c9c�9_M��#������������ ��j������Ă MAA�ZA�D\Ddi�i�%H�  �E\qi���t�^P�RX�9ς1y��{�����X�s��{�{fΜ��X���E��k�'^�`�')$���c���a]��xG��@��'W������ƿ���-&|Mf_������v�I��G�����D�M� ��E��Q��������|͟��9�R�"�����]��e�q�Ͻ,O�~3Ū����(<���4tu�}MP������R�|��X�1�����.S�����x���Țz�]���� >\=pBc��R�tt�%Q?�;���~m
�T�eH�w��&0%����h��ۉ�F�ԣd��p��{�et(����׌"Ȉ�Qj�����Y��樫�nt�{Њj�DШ0��WMt�~f(�@&����JMq��A"w�T(岹��<(��閺��@k�7q�gi�;99=����E�;e�Z �c�<�N�k��.�ymmт�#߶/��
��!�����I�����֕��MNN�q���>�~���.�s��&*j��u+�@rO����`B֎4�����%P9~�`9_&|�O ��5?�! �dcm}U������]�l�����!�&G��	_C��_�Ūcw�� P$�s�7�e�Ne:r@yUz�v�~T}�a�g77# 2�sc�yl��ᅅ~kkk���5�Xخ$��m\z�mNk��$%-����Ȩ(=��1.����Y�� nF�{4���a,�� ��I����[���� ��^�xI����u�_Z�MΫҰ���Qş޽��q��^��|�3[�ηX�|���Xm�����K�	Rd�Z�������	���-���~�J��#�&mâ���E�Ip[�:2�E�������M3��-ȱ_������.��m���6?�KIII贝��l�nrh���Ocl*.iOY������#�,rDj����D�Fݹ<�~�A�|���GCOSN��Q��gzO�����?�$G����C�'����:0~>����`�%FR�u]�!�%#@\�J����.x겫��c	��{R%
f6>�\IZ¯l��^*7�B�d:�V�@ôDx8�ב5�>ǒ��{�K�ѹ���&������;���6n���-��x����T���M��Ol�;��T�N��r�(i���C�ш�2Q��B�$F8�F׼ij��9���R�j�nQ˲％��H�hTX��|�]4&�ekG1r��nmaq��dv��%��]
�m��l�;�eR	�y&���+aUm2gV�h���"Q���z����~�nO�I��t�"R����Q2ލd���q�ٞwu�Xqq�(�S����b�ڮN.f��a:�yrH�f�x�2�_'D1iQ�B�&?.,,�:cd�,yc���N��\{ �8!��n����<�zR��]�\��qLp����G���MkTNj'�j���ެa��(L���h�Zr�>�p�P�����&ܮ�m@�Е�{�z��RM����ϒ�3�?��.�P�;�Tw�.��}\�&�H/V3���0-�-@L���d��dg$$$x�����������qF�V�V�.<:19%e��6U�.f�����c�����R��OG����0��vn�ֲ�M������Ot|�]~�@�Zb�]Bj���O����^�Nĩ���zIu�J�{���զ=H _y`��=gt3m���Bxe�j�'���������a�S���(#�kX�,19
7�G�b$$$�<p���7��b�z�1�n�P�+Tqȅ疢���`J�����h�m�C�Ŕk�@����tR6�>�^>�1��8�;�`G��a-N�B,��eV��,@"i�̤fb #�SəlNWכI-��ϟ5�.�w9�7lڴIQ1�W&�/:�ܓB,]���g9l=�����W^k�,Y�1;��9��nTAAA� �����hp�X�srWtY�����h����/ s�qt�i"�D0J�E��^��I-��g���dO����N###ަ�N��}�K]�TCA۲���j���og��ReAt��hHܻ���¼|�n��@��&YW;���@����ܫM��@� ��[TE3*�d!��
���������{)�M0ݰ���Σɒ�H�Æ�(H=1.999M,3&:�`aa�5LV��J~�L`��]'�g�Ʒ�zCV���Y%t'�f�+�um3�����-�<����G�uD_n�Cg�7�\RfFia�V~���1���֛ockI(��2R0[��%�X�g{����e,�o�?RrI%6ۮv�k�ֶ��;���q�������iW���ķ�:��y,���x��rUH��,�Vxϭ������o]�f�^u0�7�A7OQ�R�x7��;D9^�3ח�y�D>�j f~:f���Q���O��R*��h3!��qW%�����͉��S�e�(��j(�@�W�p5�6�?zc�3�pЈ��v"^^:F���(���#�*ε�(O����d/�m�D_���H�a���n=D��J��.����<wJh
��mV�c����u�Xr'c����A}ck����o��hߓ�S�pӬ���mU1W���<(`���#�Q��4 ~�n�o,��B<��yQifD��0��(Y���>��e�wj���"��-�����yt[+++���N8dG����v�����.�h�ʨ4x#ο5��Uv%%���^���I_Gr�Q�}����)��,��I璼�-j�����9F111�v��L'尾x�����H̫C˚��T�
�����7��
�*M�q��bI����S0N���U0�4������;Qυ�u󅴞k�^Ҿ�"ɻƓEwAGz>0^V;�i���z����4��{c�v��z`a�f�.��h(^Qg�3��Z�L
�����(��;��7m�~b����Y����b��������&��<��c:��S�� �Y�]��>������t�˸^^
�!4Bg~�n>A�|i�/�z�}�H��ިpǎI<�����`�Q��{DcHHH`)�W1�zz�S+T�fdd�ۯ��@�:�Y��͔Zk{oU�1֥!��L��K�ԡ��_�Q��[놌C��"l3����Uй�R��t(3Co+ơ]+�_����21Zm�R����p���;~�׹�ޚ�����6̍~��+����O!c�-	))���j&w��9γ�b��e.��u:V@D��1Gm�"J��e8'0Z�ͯÏBz��F�>�%�AL������.΁?SC��,��s�^s�h���#��{6�2�P�,���3�vjQ�E]>���PMd.��e�MP����i���N#<>�;ڬ*`w���u��燵C|R\�!�u�E"�_<���EKx � ńX	��B�"U�)?t�<$���i����4�UTRr�I���e w��1W4�vv6���q��>����:��-N��	š��Ɋ�K�����M�j��GX
��/Td\���:�-� 4�סR�'�*m�6��;�����IeS��6��n��|(�=r"�f��T :ɒ?��7��܂k�L2[f�:����]]'"""�[֜52z��.ݾUCu{���U�N��Y/@h�@h��u2N�pɻ�U�A�75�)�4���K�%5E���<�ejj�pu:���~��1�u����W��(�z6ӶI��U�D���T��?�LP�"*���A�nn2��A?1��I���6�r�9��uz%���ϗu�<� $U�M�.�jЍ�y>Ti�1��P������I���.�3��(&�,�&�Z 5����i�A7X�.�B�/a�����IT2�=��w����!׉��槦v�7 �ۿ�ؙ+|��'��`'(��z0p�o�-Zk� ��+y�)�v�Y*�`_�u�!S1JLw�Y��k����yO�x��1󳽨|���v>��u���P8�ri��(� �Z�:���%��F1J>�SQQ!Q�LSyՁ�σ�X>z����e����j��6�� EÜ̹ �JW!� ^{�S�V�<4����1 =����NBDB3W/$\�}��"�O��I�����_6�׶O��F|Qe�E�T����$�e�w���H�V(�g��^�$&[?ZD���6�#��Q���Qg%����o����(s���(&`u�M�Z�v���������BXF	Pg�؈)�:�w"N�N�2Ag��y�<�;yy�~_�em��5}*��Kx�К�A���Ϭ�"�_����M�@��:�ju`�A�)jA%��Pp)x�M�ncR!�v�E�ݚ�p��Cx�p-�q�B�#����� х+|fQ�J`�222/<�e���1�(����@��|��]z�Mb��
e�P_�bf:[p�P�r-�a"5��X��%��Tx���E�@�(�ۜ����5�\�u���]g-i������~ff{};��.���Z��	/D;���? �B�nmd熩*߽^��������^�8Q4���+�;���)Gد���o��q��n�ޔ��#]f���67��1,lK��bo�v���edf�,"�����~�/��Mjݪ�J�C��˷H������4+8��+�wm�jW���z��y�5n�֫��u��ϻHNN��%[X����g�N;��56Gmy	K����'&L4�f��w����,`@sC�s�O����ܞ��޾�9�����zE�Y"/�����dbFܬT�[,�}�B�'�e��aE(Q��75eH�5�6�K�q s>�������� �W���%�s6kx��"b��Z[G2��FVρ=�T\\��ܬ�X���TG 9�eyv�+!���[�}�_��;L�vsu��c�%�-�W>�§4���+���{閳�p�Guuu���%#�p�6�t��淟��!:���u�^�(�����kB�Ov;H���~�k#�7!��Q�^���l�甪��^g�Kn%�:�E{܎"�����k[�v���?���sHLLq�=�k�t(XyXO��ۭw�.��ASB��W��{��<�PCa����oF���-zi��_~����#�O�I$���;/w�*�ц���"�/��ݗqa�L I�}UB฽a�u��/w/�T<�5��>�do�.��R�W"����d=`��@��M=�X�y1�s�x�e���[/n�g޻���sG����/��2Dj3�^72b^���������&�[���/��r�������+_"�_��@��mm��W/�##k����R��)��/ ��[X�+L6�ӳ���d4:{�����մ��| �Q���'of�ŉGai(Tcl3J�z�����Jug�y����^):�[SV~��Q��Y��iwR�CRn��v��j�ú$.X��C�
1�egg����%U��t�śp��)�M1d|ʗ0�^GxS�'�6?�N��If��$���p0NoB�匒��KH��ݿ���~?o�Ɋ>�E`��r��5���#����$Wi�/����
�WOT���b'Ebۣ���"��ٙ33q�ק1���)��O�b���/ڑt����h�_ѓ������'5�F��wQX�e���8��zxgt���J֬��=�Wc�<�o[� �^SS��2ttv��I�K֯��4i߉���,A��R���
%-[��Q���{���Em'%7/n�C�h֋]�D�;|%�X��˫}���Z)(]��
Nx���g�<3qO�*�vZU�6��*fڬ��@�2��Z9�Z���R|"!4w��?�S�	(���XNzk��@�
�tE�ȒK%$:�1.��w�jT�w�[R�",2%��N�m��]�GT�@�F�n餖�Q�5�����hb�ò����ƮW�Y>��]��,s6�3�ai�'RW���x0l�K��- �8C�ń�'�ꉆ.��SRR"`UZO��
�����9�c	�,_9�D+���kP_���M���hF9X���L��� �/�y_u����-�MG
ރ��~c.�z��O�	�7�R"���R�"��}��H+q4���,��
|#�;Yks\g��>P����z�5�#)#W��� {q3��(�
���RL������\�2�2eU?A�Ѐ-�v9�_��x���U������֮]%+%���ׇMD13���>�Z@/�v7���I�,P�&���z�V�N@hRQ�j ��C!��IT�3�r�SA�%$$�
l�]���Ⱥ�����g��6������4KJJ���$Fį���<�LWy�K�{��Z+�U��g�ASb5S���C��5��]\���_$���Ƣ���oW8cg��I;�ځ���q�F"���^��F%�̘%Ւ�@���Fb����la����#h���8�Ի�ǥ��tw��i��V��ۅj.46:��HkίVUSc�\��>ϝe�g�;��V������C�S!�W�36�-/W}��k���ں�𣝍͚��e,1r� U�}��ܭ_�Z3>��/���!�7���f�OJ�@��XKB���ۦ.^Ak�n��*Ea9(��0��@^YzI\��ד�5՝�Ÿ����.�l40-n��D��΄:V�+Zy���J��<���=���%Ѽ��{3>��۲���T�x?��º�͖E�5[�4>���A��(!@�Xߣ͞��ƺ�tȺ+_v��^}�����)M�~s�����������N��A��q&[���q��Q�����z	a��6�#"&��]�3��RR�o�Պ.x��򔕕AP�^��?�oj��a�Nc,�������[D"ꆁ�˕����m||�
���ޝ�kPmVʓ������0uܴGq�θ���u�Xdf���m��!w�af��ե���յ��;�i���؋�rW���J(��~���/ g� �o�F�4�p�%ԕ�Sv�@�ڿ��n �xP@"!�����0��������R�C@�#��~���un�jP���b��B;ŏ;ac� t>��}f�ûjN�����%-J+�4��MiX�5��/^���z��H��5��H�y��9�~���9 ���m������!���2�ňS��w���z�����U@���70)�����;5!�5b�����/ܣ���d�c� ��=�>{���L����ؔf(������ö���۰���j1���0���+��v]t�E7���^tQ�9G���v����`f��&%3�b�'��(���I;gz��%'���;�lG�;2�R%�neiy���A�*;fw�X�i��C���*b*L��s("����w���*o����p4�ˈkD''�n޼yd~�VR]�� �3s�G�d���f�;��w��s~�j�lr�m��R����幣3�!��6|��4�d}�=�!j¦|f=Z��Q���܊�Jzi{��,�0XҤ�=�,��*���&A��@P	8�Sm�樺*��,�!YYv�RY��[�A$$'���ﶼ 9U%��w���j��>�0���̙3�(�w,�<[`W��$������I)��n��F�M<	2�xÑF��yx�}q���/}I~���H���S-Q�c�dz�}��c�xTQ��fq�E�ҚW�O�yxx@�Ƚ��R�$�?u��4���nԌ�Oj}k�J����ؠ�z�{W�#������%S��n�ef璳�D:�OJ����ȞN�h�\3^�u�\�p·UIj�R5��5��8�0U�'~����ŷ���X۽�_Ks�a�y����e���+��6���b������ 	����L:\~;5����q�:��� lh]3�s�%�����\��sL�b�W��-�G�lه+���V���W�aMT�U�eee�~��n�vO @����t�bAl
�;%--va�����`%�Z)f��!efB3�x|��������\�`�xLC��k�F=pލ��yK��}0�M��w�&6_�k�.J3V7�y@O@�.�]����dM��UO3|�[�mL���E�<�11���IaD	��ĉ	gy�)M/���\R����j�֒Vl���rr`(CorIu�� H���^Ywڣ�~��C���Ffн[����1�,z��f>��\�H�kmy�'�}*-��km� �œ��,�ܮ�a����ځy;�#��ݪ���C�#B���<b_*=���P���]~���đ�y4��ť���oc���_�|����D���2�&O+��XND�|�p!�O�x�B���!%�Y,�R|����m۾�[�z/�����Dܩ���!�\H{��5 bw�Fww���y�:��F� @8�F���\�^@�����VO\?5��WTTt{����nPM[ZZ�Ú�3��a����-L�L���F�٥ϟrL�G��iՠ0Ndt4�.+����ƥ(?D���L�����X�'�9�h��>�F��f|�c�K[��pn�U9[�����_{{�(��x�f�	#�]��p�q�(O���(����-�Ġ&,
F8���v&贠�a��I�>U���:]QQA�&?�ۮ����T�%��_r��ذcr-b���Ձ�����m��O��	]0600���f���NpeЃ՗u�n݊���x����)�v+�Zl�������ݏ���V��/�5���M6|���l�/��"ɸ�ש��Qc�����g��D�+�Ū/�񞅀?�@�k���E��*u����˻��J�/[�Soѭ�-B"Xu+����%������ ��2Q�� ӵ"�}nB?5���⒏uS�`����"���D�O�>c� �D��R�%Q��z�0�_u�J�yi`$�a~�m������f�;M�FyP�h�����R�i����<vw��Z���i���r�G�F����.��&�H̿�6�AiS��CQ��:��A��6�}Z�v�"�|�B#!SAA��1��|��~=��#��0�dC@�s��5f�gⲟ�Z����{�#�_췻Vcna1��QS��P�`�ao(@��gς�֋��EG���i@E�P��zjٟ[k���>�x��e�<|�[��B�P�x���ZQθߴ�!��@x��B�R��|s�L��\�t`����:w� R�u��|�O<~v ���w^��Q+�y�^K,�?X��.H�X?���߹}���ᎊ��Iz��_-lH9� ��vb́{%��^\�&<�A��-�lW`k���9���U�ς�EyjtO��ǈ7��� ��h_�iB�kLj���1�������6@���'A���Q������z���3�{_Je�DF�s#�jvR> (�M�"}��)� ���:������R(��*��X��;�)T<a��Dǆ��"�ب&�:zݬ������!��*�	O�{��䊧uO�8&�7U����ڢ)Ǽ�v4|�p��n9�r����ߙ���tI52=�t�#����缙)ͦٛ�-��X�����t�QC���w~��N?� o��sxX(�b_P�_W���2����;�m��� ��|*Sq�ż����7���U(�kg\T�
�o��m+�ۘ�����,�_�F3���<T��Va�Q��6�����0��]zv�cE����t}~�
0�U~��׽�tW�>�=�d��J����U��q�������3�`�O���b�?r"(��|�ԉ�����L�S�G3b[�`�h�d�KFԽ~}�2���eT��A�U�}�����Hœd�h�D���1�I&��!ۺ{�cn��[�t<�7�&��N�s���Ȯ�3�k�CtO��"�@H�6>�)0���4`��(�ł[�]#4��oڄ�b�D�����<s9E
 ��W<�%�T�����<�K*�,��1P��&1�Ɣx��8X>Sm����h �|%�{f�(��,p��w-�XB��'H�,d���QR�7��&c�W�s:�rnf@Gķ�Q�^���_����5��k��
���[wP*�o�GM�%P5���C���M�<�"M�پy�D�5��`P�{��EO$#fz"���L�p���z�������B�}N��x�;��i�<l��v>����1GE��[}�x�֎хm� %���?��׺��C��RLtS�Ⱥ��;w�خ��y�X�+{�ej*���۴�s���ձK0Rh	}�X����һ���w�D�$�6��I1��xg�ndh�*����0�*�y�τ���~�_�{�	���g�'��O���G��H_ﱩhO�KY3���'ǀ��@ �H���}JPޖ�b9�*hH	x�1|Ow_<�@�B�����x(B�������޽�u��Z����I�c�����A��������+��5���m���#��沨��;�f�<Z��g���x�_X�-u'[t�R/�z��y���l�Ak��χ�Q���(�{��	����@�֞���c!��s7U�k0��qʳ�8�Iu �1Yg[�޽�0=�?��n��/�[2Wc��;�f�֕���F�K�v��d���Ok���Xv�M�P��\<����)��@G����d��iŵ|
�L䙬P���NG44�3�=���Ԥ|�3��3�:m��o�~�UBB�es{'�����Ŗ�Nc]@�$ �M����4F%��=�m�M���DA���&_��پ���7��d3�fh�x��]��>��n��]ml��M�"T�����ެ�F�//�(�b��u���L��� ~���J���+�#�r���[JH�����/�i��&x_>P�R�;DK�Z���hhr{���<�%��B�(>��3]#����HMFk��%�����}Un.�1Z=�O��w�lS��4�B7'�O]��d(����-��.���s$�[�@����7�B����1�@	Oi�h$�c��f(å�R��k��>"xr;�dʜ�ԕP�%���R��%n�8�2��H� ���a��];4D�v����HEEe�{
b����j'�V榒"�(-�M�dϿR���kh 2ǯp�jQ�G�z5�������'������$������=��D2O�G'��߿��s�(C)��g3m%A{ݦ>�N��zؐJ��聉��v�B) C">�� ����u�B<���]��,f���:��ŝt���$�X��ϭ�)3&
a�b0T
��쥑�B�bB(�@L�i<3�	��T���@+/�mfR��I?�h,���{���*��-�z�mO��h̛U�d��%/��6r����8�>֋{��q~����5�O�����^�hȕ0�����d.?KXQ��N�H����� ��5��_�ڐ@� ~
����$,�@Ծ��p���-�`t�e��̫��>F�	Q��B[<<�ݩ�*�ljz=���e|�/��K��#��[A���;��K�w0����d/��_�@%�_L6�����:���� #1����T��l>�C��6��^L,�Xt�c����n.��k?���
�!Ћ�\���U�۫��W��|�
��|Ƿ�vW�ܚ�l|�L�hH�Z`�P�SWs��U�6��)3�d�;"5�v�hyy9���Q@�*T���#� q�����V�O�f�����훆�n�@��������"��<I��e�ԔaхꙁS%�����q��gC���!��BހR��R���].Z��'����NS�˽��S����X���51��@��U�de=�����EFFb�2�)���������.�AڸriK�
J\�.�А��K�{�L=l&�%� �tn=zLU �s�YT�k�怐��*�/ �[V�I�P�#�?-��S�2�Q�f8			�^_ҫ��鱣q�M�8�m��aˍT�G�Fs  Bи8;;�&B�22�i��Tz��������� X�hwvpp�.��>ӷjhn���-�#�DṶb{w�<,�f���ph�ݍ�N��1W0�-�f.�ӹ�����v/���x��I~���g<�~n�9�#�CW����4��UK������UqkxE�U�u��ԭLM��\m� �
��+�iX��d��`�>H��K�`��?D4Uƈ��1���`���|�-f6�����e���!�'!�Nm�Em�|���~���3��@𼽗���칾�M�DN��U��2g(\r�L
x[f;	@���?��= 7*�s)i�::��knHYZQY�/�jL�L�M�7 xTTT�nv�=F���P��3c\��F].�ı�<"1}�͐�C�%q�U�sK�P�A]�?k��ܝ�X����?��#;���bm�w6&뫸��{�h��

/>~O46q��P�ݕ�f���-��T�;����3�D��T�*�rN�};��&�V��$˾˄��Y�p����DW�z�[WRRZ�=��t;��L|KK�������Y1����|>�ń�U���i`�Z?�Bu#t!�v�L���WI(���-/<��O55s�5���� ��XG@���p�ډ]���h2?\���˭
91޻�\ ��k߃Z��B�P>�98�HQ֋ET�>�r�W��y8N?	�(�ĖI�g�����W�gK���cBS�Z�z���,���l�^k��9B��u܌�7�>�={�=�u1/r���3k�Ua"��(�|��� ��''��yϚU�I>Ae�J�@y#<^?Vs����;B�=��&�NpX�I����nXoffv�kL��%0�(���6a[v>�a 9���yCf��E"�)��`7�f]�$�]�٦ŭ�֠Ya_��o�%'51��؊J� � #����nY&&&ݯ./�s�n=�h�t���<:<��a�r�_�v%�s###�<|C�^4d�u��6�Zzz�V��{ѴCx=TX-B�n�-�l5�T��u0a&XQ���yLNf�:�U��VA�WEd�HNps
7��Sm�P�[ʢU��gH
^�&�T[n��BLCm�n{�sZ���X�����RJ�@�Q^#�����B�쭢dD���_����x~��޾��N�U�f�'�X"k��B��Ԓ�?zNZ=��=��'&�� "��+ٍ�yѲǵ
Y��"^�0��������Swq&$Yd� ��)@���'�'!]H�����i�B!w�ݣT �僄Y�Np�������q�΀�X�J>B'��n��<4hO��˻M����Y3�Ft�gY��6f�HJ�����aZL�?b�7������C�&�: |�K����/���.��v�=��bD����
J���ǨIoz9�+�<سn=�Ye��r���lvlvZ�t�e�5�Z�O�����L�V�����]5�<а���p�&����	��R�X�޽{�sc]�Gkk��z����=]]����(���/P��D����?�d����db��J1� Xb8ɠ[Yщ����i�U��GZ|;�����?a�'��E�/�j�*��)s�������έ^>8d��X�m�����V����5�[wb��kk��YYY!�Dy���pe?�QQW9Mc;?�H��A�`����`������a�TS����C�P�ц���b��P9�,L ���S�=;�)�DwRy��ʻ'v��0wl���#PӽU1@)��"ؑ�7�#���K�s��K�.zz��d�>\L����ˍ
�V����tP��_u=�m�77�	����/��;g,[d|����и=(�w�����i�DN��)l8,���NM�;�<K,�nG84�V�Mn����-Je���A5�)�Q�׿��LNN�/|���no�g�2z9��}� DcYj}7:t�F ˿��q:;��� �<�n4�~=��|0� ���6�n�V��봰6��k�9k���4���\2Z�=|��Y:F>/�r�2J����T� o��%k	� G��MXweT���lƘ�@�V�C����C'o�!�u+�Kp@!�O�Q���2����m���]>�OXX�u�$������=8Ce���Р>+Q#F}��[l�C3�c�wo%~b+��O����L�"�v�<����:��/uA{�E����$���y_x��ꨗ����?Z���7;�bqk{�奥W����+�AN��U����j���[>\>��ȓf�K�}���Iw�����!=㶮�'-��s~��H�2�qv�Q&;f�9���A�*:��_��?�1��ۻ�+�>���3��A[�JbMi����8����Zb�Ű [�vOV>�jA26p���o�q� 9�Kk��핳�_�ĳ�g��uSܗ&�R7J�5�2�_���A���*�E�.?d��9�m��5�1rAΨ*�����ቭc�������;'v�ϓT����B3��"�S#��i�P����@n�����q
oNC��a�zdݕuk��ⴸ����z�V-�����}Z����!��.M��W���P8��dV⭩Ke��YCé��������ު	T���{�` ��`�d�k(V�|�"�2�c��o$��=E��o�=�X����U֮#����7�U�Z�}�Ү��$�~�M�T�f�������0����dts){�f�)a-���� W��"�����\W�����4�u�zu�;MMA�}��2������v��t��\�>#L�N�1�!Ԙp3��.���c_�*���P�aMbU���WTU%a�>��H���'�r��E�8���:bb�2�߱�1XM\��)@k�q�X����/��q��JC�8`��'R�󟣫]���I��>~��d�Л!�{�k��[;�����ˠt��(��H��x�K���	�\�<~�Gx4�A �\]>�ߥx`� �wT��@��Re�%���6.9��O��vx�����O��ʋ"�i��}��l�V�]/��$����]?���A >��޾��o`0��<���+���͍��w�$'�$�m�Be�_Y���/��,<�^��i�GY~FX���G��_;��-<З�k�~)�'���T��@Y-�2�Pk��)�Jt�	z��X��\�����wa��*��d�Y]�x�{������OK<m.] ��/#`u� x��ټ��7u�ఓ4��c����"o){�5X��a�v����yx��>�����4�b�_�{^Tt�����Jv�Ganx�CzF$��Q�6*3�X[�:Z1j���@��p���w>Ʈ@ȠE���f�z��s�	R�G�'�Ĳt�U�X�R�{&�ߛ��l����S�ј �_����!t;���y=t�p��j����x q ���ڵ���.��p�I�?;5���*�8&V,]��1X9|���q �c��p���R5C�#\Q;��L���Fn�qOv��i�<x��vAI`����G��� P�6�����N�i�A:�آ>1�v���h�Ž�e���^&''�9\8���~��QNǲ�{K��^w�ݼ���ތ\���>������m4�*F���4þ�I}ߢ��*%t��\����]�{��QJ!��G�5�d���o�'���n��)����>�z��R�����o}��K��5km�[^4��]Q�8w'���<r�����-�<���5�*�����*񓉿`{�x���}�v�������8�w�#C�`�g�����8�HUαM��s3)od�L�\z��ʓ����pF�T?��kn�v���"""�\�l���i��'Ŏ6����m77wZ4���j��=�\+����Tu�D:�Mks�.����giF�y�t�@�u���y%�S���M�	���_H�Mݙ��W�v��Pi*?M�ƞ�D�au�5Y'P��w��Br���X	������q�"�^/�u�~�9]N�BU����o�W�Pu@�C-�������5o˟XE��v=ټ�������^ǻ�qǢ�ϑukN����V���1ڢ��6�>�y��h����YKb�h��������R�+�Ŷ��j�#|�Rvm]��<f�0���}�*�����yA=��a#�2�7����������뿱���!җ��M����Cs^���z����T�]������,՜+l��C�y��D��!���300�@wܿ퇉���9,��L���m������'1BMH�l���]v�a�uB��Ύ�O�>f�����Ox���Ii���))zIu���pZ�, u�TH�Tz�j;�%%� ��^�Z�����?I�˝uLw���2՛��3	w�� ��w��y)�fo��Q�^�x�3��~�a���i��6['�#3�$��d�����̙^�<y-���4C�]��+��H�#J�N���)�9xpo&�]�=�N�Lo������
MMۧv���=��+����+r���K�$6��v��1V�a]ۈJ/L��j�6�G�;p5���C�c�c����&��%-iN�&GF~$�9��@`�s����orH))&��B��3�9�Ƴ���_*�~A�a�����8���m�N���X���7r��hIV�|�9�����u�U��m��M��ʡ�y�1U>�9�k�(P�/v��v��6���I�"Β��,U{�帏����0��K2h%��ma�{͎��M�x1 wz�d�6�*��Luh���)���yg�����L�*\���{� �efK���!��w�2E��X: 0��
-���'�����kHs�jD�WO��<)� �a�M�E��G7`��R�ߏ?�|�K?)dĹQ^OLU�&zU^��a�����=�a������/ճ���`��xq���b<?����TJn���Z	;��hp���C7R���G���8�M�zބ��w�~LM-�$P�������\���b��{@r(a�|����K��yŜ��#�U/C��Ƈ �$�O��	�lZ� )�ݖMt�v,e�03ҫK(�TOWO�GA�^��L���!ef��2���P0ˉ�@h=mnBL$�l��DC'f&�8��W�Oo�{s�W�����Z|g��3Z�A@�ec��]䕥2lоV�������8�Bm_ѐf�G�$�����Dc�����9WB������F�Xt[��ޓ8Ҋ�ɬ�{����L\�(a[mB#��;@�?~��=x�3�9�D��ȰJ�ղn��SA%�SM:]-�j��5��P���6X�n�U���Yv3W�,�3�k�sg���s�_�R��T�)���(�F�1�fB7�O֌YWT�r%���e�y���y���r�R�C���'���mG�>c8�[N��4�<�$����i�[�@e�Y?	�A�֮�q-��zM}.�RC+����k	Dcn��$Q#�����f��Բ��dMؿ9�(�v�K�̾*O3'5ѝ�K�'���NW���f��У.�YrYB����ܻ��{`.�+j�{�u��Mt�XX�r���t鑤͓�|��G��1���4�&�ߋ4JNpncd��j�p��@E��m��S�mo����ڦ���9{y�T���� � �'P�HF�f��=�a�'s�0cA�3��x��f���CRBܴAZ�AJ�Y󃰐Uԋ�)��÷��05�$�Ct�&x?&7�/��J�4F��rUc`2����ڭ�X���|���I��2�������,��vZ����׭3[�4⻂JL�&���h)��\?~��aۤ��iُ!�IX����L#R��H�F'�'���g����E���o~B��Zq�3��m~����C�����> ��������Ig�Hs̅7�Yt}Pa�-����1|���Le��������d�efp��C�����h��_��$Y��������V&Q�:��k�@�FN.i���C�$�޽���u��b�7�w��+��y���{��_�]D�Dcb¹-��^�M����0�h��y�$#2K_��13c��gX{A�Z����[հH,+�����7&����IL/��������H�W��J��1#Q>y������z�bE�����juW���4R2z
0z���R��ϿrH|Q��Ƣc���V�D7�XQ�]>�@����-�Z�a~s��1�[��7V[K
�#ď\5�����
!�{�L>T<h[Ĵn4��	����<|��Z���-��P�m>��C�'v�p�NJby(B�����!�B��L��b����p�`0�L"NQ�������t�^O���)��*�c��h.�V|�e������D[X��s6`O�.T � lۣ
U�ŭny�Oo�i�7D��v�:�옷(�������v��s�s,���c�6��ل ���x͝���$���[]���i&�Yn80�QD�Ɍ��	�~"�j2���HꙕC�����(�$�7?�X
@�1�b�[tr�n]	bq����l�t��BU��/�(Þ�c')¼�]����	�p�/t/_�L_�sn��T;L�^G�>Ļ��8R&&�gQ􅥺���6ޔC��ڞ�hd!��G6�F���(�h`��]4��@4_�YJ��ѿ��E��!��k���%~ q�Aa.F=�2R��6s����G�����ڷ՝S��L�!��Q
��'���9��r`�my�&��v��z��e�{��&R�.����
�7����&�޹Ô��=z���
46����@O�
��.Ԩ��l����"D�0�U<��w߷Y�����$�m	�a\q��QM����L��)x�O�`	��B!���ؓɤ�i�<�1�a�c˒��߅����t��;e/P	��.�c=�*H)�"��
jf���:�f�A�d)$&��L�m
��G�z�/{��۠�fy���=�6O���p��qH1:%�6|wV�77uQnL����"3Ӯ��NuAN�{W�x5�k��0�v�|O��꜊�PV
�su·�`�s�\�3�~�k��95�M�9�H��?,���wwY��%�'�@m_��b1=4���!����h��Xo��8#�~��� ^�
��`�jeG�0��h�/�) �FTD
d48�Y����dZn@|�m�_����A4�΄[�����5oNj�u=b��� 6�e� 蕰<W��73�3cU�	�0m�&Q#�(Pl��[s�����0c�J�n����v}<S�%vY�+�����󇣘3\�G���D8s�����D{��_+6-��=#zg  ��PN(�lԧjL}nX!�$�[^4Pw�d��²���3�ݾȡ�by����@Q�'[^@��A�,gXx������-Df��kk�P�/ac��k����Q�-�YW�l��->S�O
Rp�$�s���R��֏�"�*�A_�h��͌�&]G��57�8B�ω��v�z?�����@E��2z�P����Q����YZ�8$��n��ͫ��^BwYh��U9�y~0��K���	�,5?l��|�?�M���:�rTE$�6��Sv؊G��<g6llC+�K���W����de�Un,����@%~U��0���������/�Q�m�������:�O�?�b�b�O��rL�ｔX;f�|l�������@3��C�a����G堟��zhl/pfd6�LL@��V�\�d-Y����_fl�ņ��Q�yltX�Rֱv��le�$@>7���n��E�L]�Kגd���>8���^���؆^MN�(X����kW����B��5�B)Z�u[����4ڴ̴IHBj��2�$�1ej����&-ӪFj�֩���=gr�Ͻ�{�9�����]�������sLJ��"��4�|F�����gjh'�x5E��K0/��8A�`���,��!]��;�|q�+�7��<L�-�>�A�b�h��IZ:-ۭG+���u��0�D)��C�Q�&��+Zא�W}�okk����w�IAHi��B=�Y�X�����A�xMwq%I�2���o�$�*�$��A=ݪ	j�:#�l]T�'WQ�m����.x|<���L��������W�Cci�w��Kx�QbE��;�o��pJ1b+^I��{T�^���,���	��:�<A�yF��"��P��<$�eB�"X���=ɡ��ml<���'P�����Lh��il$Y�Tf�P
��C������{��Q�-q|��6�^��xR�c�]�&�W�lW��ũ![�����%8M���aE2N�Qf����ݺr$��OY׍��,V�(�h3��Ҕ��_@kTu��T�"��PW��T/j ��o�ow��֏z�T+�bZRK�C��#�gtY)���m������{����q�jެ&D��1
7i�Rى����9=�.�K�ܑg}�|��rf";l"��pz�P_��
=�����TÎ��WG)�K<���gp����ռ��H-k��ϺȚ�n�`FN�SY��ůۈj��8���>$��p�����׺��39H������5ԯ�/ V HRX2�t@���S�j�o:�~����P�-�҄�~��F�_5-~Gz�uF� �h5�2����눴/���Bj�6$�"��ދ�VP� *��-�r<����y�~P��<˝�d_��	)ӡ%^��[�7��Dˢ����͌DÄ�U6H��w<Rp �YD�h��
I Z���u=��I�
KZ�I�ۀ�Hĵ�wȀY�Q����h��R
���Kcd�HIIi�� `R�^Q��啄L���n�0�%5g��d���R>3z�`��8�Z&��+����"HD����gQ�n�n�!��e	�7�x��y�F��ӈ�s�:�܍q�ׅO�d�1>� ���<�!gK�͔C��#�u���0�!}�U�v��L�����>?Y��r��rVU��'d�4�ƌpc�­�C�]hY�o������#k���U�T�g����.q#��X��g~�s���2I�vm�!/��f�v�V�[H7D��n�k|~C��4~�jw~���ˆ�󝕽�2h	�ɀE	���GѢ���}�s��0�/u�F��L,\�J1X^7����Ul���C\��m�QUi�����tVR�͓�q�b����Lh�2��yl+R���ejBG�)0\Z�����Hҡ:Dg�״tݤ(�вaTVK�JН����A�O����<��0����0�����ܢA� o�L�,�����u���s+G͔;ۢ
��?�Pʋ������#Oٚ�$;C.���6L�zt{i�����y��˵(*|Ӕ��B�w ��+M���
�$UeG_���t�ؚ<�U�	쑠��*��� J=|Od��[�I��N_
_v\}Uf�`Lﮗ�2�ed��\X,Vo���փHi�ؕQxB\1 TA�#���;ri~��RZ�wv�c��NP��{��+���:�N�M��fn�Q1��0��MhMK
��O�Jn((�8k_�up��~��^���������f\�J��G@�re�L.	��17�2����hB���lP{�?8V ��bK��3��짼�Qt�(�V����dUݏ"�<2%P�'��%�73-n�C�W'�$�����0W��;�մ�tAXY`�R�>�
Xw��\�D>�+�:)ʊP��<�2+ `���ڐ]�#�����(9�
����q3��/�@EI��z��)eeh�	�a�ܢ	�Vâ�B��ىG6�K��(n*�0/�/*̣,"k��C�ޗ�����u[���ӔTӤ��>7�6�}i0%E�zSH�3� �f��Rs�]�_mG6���>N��**D92�4#rme��}lH�GV}���Ɂ� ��Q�V��s�$��~em0tHE�Yyx�9YLg�0k��z-������`��u�V�\l����p��s?���Ɣm��v<)�~}�Ŵ��st�@mKΝ����"�\�ʎ>S�4p�2م�����|�bA VuA�7��~��.��B_�B�w�T�����_2?�h�NY�ƪ)���[���_c��;?� n]�2pnm����V��LQA���3&3��f�͚��͹o����o���Y���ە�X��n�XQ�XP*�·xAx���e謮N �'�G��s����O�T.�Q�2V����++��ؑEu�	f���C� Ȕ��	��'d@n^2�* �U%fI&��M�Y��y鏏f���x�ѣm)=@ ��Y\�M�����g���?CA9R� �*Q�sA(��I��{�N��77����q����I���ć�D?H����$��)�h�D����Q%~!���C�Q�J������H�+�{h�� ��t�5ٔϫ�`Ƀ-S��ONN����*��B]<xkGD�jef}_��P��t��Qz�m(
D2v�>H��Ǹ�8�	6�7���3�$��(5m[����O��Z�����(����,�ݰ)*�����g^���е����>>�N1;@[/&�[C9\m�j���e�����S)f8Ah���)�w ��(�
Pz�}�ywC�k�Wu�	�������8!�0�������6��,e�b��\��.�|����g%���q*��B�R	��d�>��@VYoR�%V^��3�*��A�694�qA�MҼ�%���Z͍.�vq!�ڟl�P��e��J;	��\pLo
6��6���u�P�����I��@�w�Ϯ��/˛�=�SD����Pq�z��G��{����ܷ-h���s!5"�����9�a��?�rz�c�@8ňn�����7j�ɵ�ؔ �[��E��.t�wf���Ҹt��j�����f�I���1�0�{ ��:Kɨ�bS'�p2��o*uV�D����&j�����t�{��v���m�Ƈ09.Al�ٽ����&��":n���\�n����J}N���GMF^��@��!ڟ�w" bG�;�H���|E�{��k�D0?Rc�����^C�͡K�%��:��yg''&��)7c�4��#�J���R�Y�~���g���oŖ|��� b(د����Ǭ����*r����p͚���;O�2��,y �R���(���?�b�9J�2�e�#�!Hk�2��~��^�V:�����{�;�>?K+Π������Ȁa����	�*JO����_����h=���g9�mU�����a�7O�Y��+E	"I]"����ڡ���
n�k2�����V$K����6`o�״7�^�X��k�"��Ҏ��S�9nn�q*u��ɱUXl�)��Ԅ }����u��>���vc�
[�繞?+	i���iu<�^�t�ڄ��l=�գ͏��G)�r�ҿ�tz_U�l��~�Gř
:��5̧p�$���� �\��НR�}��@��j�l�Nj=�V�iR�i�3?j���B��Ղ�6~��F�ی� �m��q���0�3h=�qĎ>���w���L���Ec��ؙNl�i��ψ5IL�ep��	h�U�|�0+Xw��
;�1�C���$�����Ԫ�`�A^d=*���5�e��~�T���b˒�~�)g�7M��ݔ�p{g��X%�R}�DMg��c�j��^t�x���m��J�.�Z��=��/��J$N�<�k��"e��V��^8ß��&��e�V]-��EcX9u{}��7ى�ѷd���aJbD�ʏ���_A�����	Ʊ!K=��u�or�n20�7�Z�(	�����1@JR�&0�������\A�����P�vT�X�B?�<u�q��}�U7�x|D��g�����)t;dr!5d�&�<U���^z��)�"n�Y��)�5�9��l�+����k��P=$�����)!/�U�`���-��'Wnk)��|��p��+L�8��:\�0hw)�$�φ��9�=�� ��T_�����Q�<�%��r���T�����9D����p�\�{֕iL�t�V�&��rT4��[li܂�<гڷߖ<j�N�+�����q����N�4�ݞZF#���$ vTe�B��~Vx�d�$t��H�-�Ub�
�Q����M��t!�����'̘���f%�4�s:���M���7Ц���^��4G��؎X���Jk��$�ۃ���m�:�s[��쓂�ؤUp4��No{y|�R��,O�P�\��`�S*�&[�%㏻f'�咜��^4�=A���A,9*��*f	���M[˹ҡ���3�.0J�H*�ҙJ{O��.�6��6�^�d�������k3�img��˺����y��?�,vBx
����BV�˽E�A}ׇ��+�O�#=t
~$��tIt���l�+����ꦻhX�_;�����Sߐ߂Z�1Ur��x0@߾$���8��υdU�%��a�D��F�K0���vvT���ԝ�g4HDr��s�y6��G��uUUT9�y��KD�\�S&wmg�� �E�4'�bJ��}��'#�P������<�5����3"?�9�x�Y����xv'�N*���Я�?F��m���T妌��\�:� ؅�)N�%��� ����xň��\�āj�q��u�B�Y �jT���:�9ъ�e�~��V�T��Ր�"�p���ŖVn���I�F���I������9℺m�U���k+i=�� Ќ_��諬Q���Y]�����9��L�,`>�d�y_�e���|T�Hd �x�z4g��@F~b ��"��OvĖ����Q��s���L �e���8��F?q���{'4Y3�r �?�#~�/�`�N~��(��Ӌ`@Π_�)��#ܬ�
Y�o������R�E
��Ub]p��$�Ѧ@iB��\��P�sb e���m�0!��5{!�-S?��81���pU|~��H��UW�-S/�?�4��u���\]����k������5�x⯸pz7�������>����O]g��Z���V�{����GP	��z(��u�Q#��ٔ��4�/�S;-p�3٥'w���u��	P�:�{.U���f�&��=��	ƈF���]�%]�l1~3�'�]����6�c�����>�޳��@ˍ�q�x��b�;��E�Ae�25ի�=
�ՙυ�A�0�p�%z�`�����5ď1�P���z�'�ۈ����i=�.��㫫��nU}*���e����BMP�������4��:��c@��=Y��A6&��e�H1\��p�w;����٥!+�#GЅ�]O(�8w��@($�8��,��@��xָ�X���2)3�:q*I&������h3�W���Gpr#��4n�=����A럂�+��ۜ�9���lquI���,n���M!w��8�>�;��/��sSx	�uKD�h�WV���hT��E!�\$ӥ|�^ऺ��RՃ|����,�d���ɾ^<��{����4'5��)����J)=Z�P�]8�O�����{�İ�x�w���m%�<���Ҭu��Q���TYF'��;�*>0rs�fM,M�������i�����>�ǹ+	�������@=�lh30h�A믛��\ŖӋw��r�����D6ȡHL6`�e��p�1��Lߥ$ӽp����3���@����U��>��1�8����g =�>Z�u�D^]HVJ�"GsL����C�	IF�e��e����XP t�k�4?J���K�8)]˰���#�T6����ޯ�wm۸W��NQ�v�,���?���ܳ�9����)%�n�OA��{�8���eI�'�ڧ�I`e�@S��O>�e�)͎�%i��@���^�>�p�
����9��~ھ��:�z^X4��3�#u��o�C>����� !U.����7�^oRݢ�M払kH~t���+�d5��! 5:<1����z�!�U�U�:l�yM�������`[�!l}�^�DE��,YZ���J�󃛹����0'���ك�O~sx-J��C&@d�a�O�G��`�p&�R}��Q���Z[��7����ꝫ��[��ִ�w��y����w�]��Eb��B��#� v!�,S�����¤r� 9��%{e`�hˋ����K��:�)BfK��-�M���t��9+94?�17eبu��-�uq�gn9��7��ng噴�}��v
;��[��=r��Rrު>ǌ%��E4V���n��u�t�=F�A��R/�ܝ
s��
,	�i���#f�9[��ھ_��z�e��5Gu����6�#m��L=�����H�
Ğ��F�����[g�Jg�i7�T��p�p�VkK�&��j��ߴ���#ძXgO<q��*a�&	�52���jæ�����˔����4x�H������p��K�z��=Б�<�<�7�������>#�X��%W��5L\��:��UK������ȗ+2��r�`�"��"���U�~��p�ls?�5�Ͻ�{�����ɓ� ����q�3p�}z��H��Ƣ%�k�ƇW���_0F�؋��LCټn��<�K��\�����
ŁwEFH�F�2�J�P�c���xv�7f�X,�f���eMKbT����;�����+F��D��#Y�%��t�m=����7k�ȥS���y�)5̧�>�Th��}�ޟ���P����O�7����� �m�ОJj���q�y�ql�ǭXҺ��K�N�����V�Uu���*F o�#j!��4>�{'Wb�V/|U���I�y5�+_ݨ�E_� �B�b�}w�ˤg_��>�藏)�����ΫV��J�>��\����V�	|��Y(��ִ��񴞕=H�����r��ִ����6�&Y:#o�X��5�z���s�n&PM|�E��p�R�yb?g�2A��4$��1\$�AW��\�:���{7G�wU�(V��=*�D���\����@T��IX-����	B��2^q	Cf�A8R�8��"qj�����|�2�!AAi�	�S�N�E����O��0�s�k��!L���4��B����LOW9�]��<�j��)�^핍<5Z`B_��H(=�2�î:˧ǎ���JF�m���u�қ=	��};���Px��d�]��X�q "H1��%'+C�5�{2o���fHY:
��S���u��X�����a�Z�)�/	,t����݂?����/q�J�T��X^��듑7CQ:t���#��y�S�
�M6�b�l|1�w�9Ã�ާ��tI�A�U�ꈂ�F�3e�3z_N �W�`V�·��'��3n�{�}v�&���C44 ��#��P�vW�
d���˽x�����5�z��Ͻ��,@���7�X:����J�*u"p�S�t��!�Mk����Xx����%S����X���d���`I̓��ȉŖ��t?����o�J�:<��2.`=�V�����|�ҊsHd�p�� �kv��=��q�冊r�Q
�V���Q�/y
�o�O�	��k���Z��H����C]>u�s'�0�J,���l���,v�
�u�J���Q�=^ڴ(�O]�M��:����+�0y~��2����Y�$��6G���aH4Me����z�V{����3�u?���܌8q�����J�"������⦐�G�׾�G��5�..���eǷ��6�w_ǒn�v;�����u[��`��'d�m\-��sE,h�E�Y�rB��'��=_���@$R�l�mpnt��Ulil�؈���ν�H�/���	��̴o�=16�&������df�ңµ��ҋV�#坨�n�UK���x�����+RXn�j��a���q�Q�0-*�����.�f����h0�K*[�
��ŷ:&z>%w�7�-:G�J=Ƈi\��.~���"
A��8�vJc�]u�uc�RAn�c�V��K3��9��B���ߐ��{���ϴg��<��u��Tk�\چ��q���VǕ^e�5�/�Q�����K�e���2���^��s{��"M�p�,sO͚I}C/�2	%=�o�t3xn|D�u�/�ۯ�>X�|���g4m#b\sL'�\C�IeG_Z���NYm�Y;��������J����e�X����� D��w�e�g N���V�X���^��ye�;g���Pw~}��j�R���R�(��-n�H�"����J���π������G��CD���2@�|p�1��Y��׋i5'�tfH��r��֡:ē���x=w5�	2���^a��q����
\o�
ը(�4����ȅ����
��u*�"�o��!�\��򛁫r�࿅?�T�uF�W&�ͪ�7IL����n����`/d��9p��L�KS����$F(�U���@�6�`�1�iJ�Th0+�z�n��3@~����K�=�ߊOԬ'/g�& ��B"f��|Hݿ�7aZO[.f"���h[y��lB�x	)�ꔠË���E:�X };�X�����s�Tlu\�>����b���<2��L�[��9��$�,s��=!�� �HR);q����ؑMe时ܭl��0qy���j��������wHVAC�;�*��3��UF_�3�����>�����s��$�j6�T�죑�"�$�A��Q������2>.R�٤�{пI�[#��B�Y����V0/�v���nCۉ�AB����� /%;�}[*�BkA`�e�+�NPS_�j�RcA���r���WNK@<�'I�!Зo�N_SSͺ�tu���&���@�Ȍ�vdnJc��^����_��?�[d�,�y]>�ħO6M�2Ȉ��Wʛ�F�X�_f.�@$�o��x�}<��0���󲀤.uI�"��/�p{|n��2�%$�����S*'��$G�'��s����%��aNfk�-�4�=.P�'�j�F��!7��{ŪĞ`�2�7e����~r�a��!5g��=U�Lm$"<}<�=2̼�=��d�$Њ-���9b;�{D'���γL��I4MҊO�ۜi�V�A��&ܱ�C���-��U�5�%�
�vH��W��
$�����F@���7}0#����`� `޵*�C"*F�:���.[$We���w�#œо/uu��<��B����t���	������=�~��@��%9F\��<Ͽ�����Iap��E��8M��,s�w9u���_ܠ��$�A˰Z׀ŐI�L݅e�9���ݳ���N4E�+<�{,��k�jͤ���'iޖ��!��'*D��y	a"���H̯q�0X��"�|�+��q��Yǌ���	���G�<�$d����mk�����?�Ѹ���a5{8�\�)if���k�_Nѵh�:PF6��w^�<�(��Gk!���Ʋ�8��܆������b~�x䢚L�D���Q�r�P|j��:q��kBu ��з��s���b�Ě۟��&���)�MB�Uvㄝ���/�S�a�����@`�j`e�T�M9� C�Jp̼�Y��PS$\�A&�j|b����Z[��+Ig�O��`���B��s���|.N�
�h��z����S�h��Ye�i1��?�/�N��Q�^j�b��딖�ִ���GY�^���3�*��1a�Fp��: �C�bA����-0��Q9iuZΝܐ��2ޑ���<�=���q�jS����V"��	����=���F1�^�+��W'��ݥx��|����Q��@7X�W�v���Z&DV\�J��kr��5ή�e�4�n������n���]j2�����}�I츔����G�3��	<�=ئ>�(�zT7/�jfs��u��ߦu(������<u���bľ
C����h� ]iR|>��Z�b E��%9�M�,l	}VH�>?pRk��`}7�g���`��T�ˏ#���2c�j�r�
[���{�Z��b��>rFM��4��)�V�t���,��Q'��}�� �'X8����2d����}87C$��1��h�L���f"=�Ey)\L��QlyL����s̓��f�]��Y��c��o}���
��l����r��l�-�|���agN�%�J���Y��֒�w�WL"�ʄ���C�-#R1\s�����������ak�Z����xĊ]�X��pe��2O���B;�\L��	��7��v]ǶR�A�Nh�qB�S�g9���D�*�w$<PO�+q}������x��S�c�N^7Y!L?�Ɗ�kn�q}��se��N_l�>��$�P[=�]?$��b���##z07�,�#��d�]�ڜ�W��j2�}�k���;ac󐧴\ ���5��R�����PË�*�OM��#��i'��:��}����X�ܛj@����W�)��%ղ
?U?	_�*/D��}��ed�&n��Y��4mEۚ�˗WbI�I&N�ԇ�$Ӕ�L���B:7���ZBab>��������%�4�*e/������q'��[V��?G��,�y���}�*)���v�l���MC�t�ܶ{M"m��H˰�mc'����O�ұG4���ٖ���f��A��@�+A�p��#���C�$K&�}j[��|�4	g�O���z�,O�s��N�Qz�=u/\�b����=�w��P��4��g�g7���Qz�j�8n�	ͻ�3��$zȅ̺U|f�j�X�~X���'3���e�}>"��u�#4�Y�f��㋴�/_��r3�e�w?��aa���1SY,w|-V�[R^S-�lPP������j݊GVI���S�R��j�͉e13v�r�:;��4�71�,�`fCO1��C[��2I���������mBoa�m���R��Bu��f1/��C�+!P�����aA)����!������k���G.�
_���~����0���!�k�|܀+n�|�,��r*���]u���W����z?����C�0��ۙ)l�X�c��P[KK+�ZlB�9i��yIG�������'v�2�n�2����D��y�9c��Ea��S�3�[d���5��Tמ�ձmd]�OϬr���̨^���V]'�Z�t���%&�EEE�w��=-%e��u��L.^\2�����n��W�o?7�}�Q�����L!v��7 n���S]��Ȕm�I��}��~�}�F��b����5��JO�J���i�Yd�`<мY�36���]aWߡ,?̀R��}{��y��7;r�K#m���}ylfX3;�(nɯ�� ��ҹ
[��I��~�c�������MSRR�;ܽ[����N����7�_3��]�IE�j���
r��@׫)���qx��B,Ľw��w�RO)F�ыJ�1��͛�ҡ,1WA��t����C������T����~�	��p��2g���-4��ؕ7Q��~W�=��|�Z뗳 \l���,E�sد��<��f�R�:;!Z̧�'VJ��Ě$Vfmո
�j&��`��5��1|�T����d�S��,��~��|o����m�qh�����Q�θsh����ǅ��/wk7�w�*��`"K��SE����3*Ȫv �ʧ��Ыx��p��㨻b��5�Fj*�=��-(��e>��ic�(��SfQ���0�m�q��7�&�L���M��\~w�V͓����~>�g���`2^����냅s��7�rX�1�P�h�9����+?��^  ��7��L�N�5^�e}�@��P[�}7ke�G�{/���~p���^#�W{��U�����-��a����(�iZLy�7�a�o�Pg�i�xr���5,���=�ͭ��J��v�(�ybL����E�?-�I���Օe�a�b?	�l��у��3��`FUK��9Tّ-��Fe�[~f-�5gtCVT��,���h����)�3iQ������L��=9EZ���	h��XO�1(/<j�n��/n�r�-�r��8f2��bL�'���}�'K�vm��E�ڵ��Ìyc��t1��;i,�~�� E��d:�2�����`+�H�m�X�7�n��a�T���p�yr�z?��Xr-p�]��$w�aB���U�9�a�ǖ�� �duw��x���<<CU0��e�3��O?�Q���$`�⅚r	RoI�F�#�D�v9YVd*D}��❕��T�Q�������_�7�6��^�8u�`ۻ.N�I���l�aΫ�}��3]�|b�3�F<BuVm_�����(R�ܳ�	`KA��U��@�XL4M0v�h�/����jUԏ�&e���6�������/�~���"VR7��H��dt����uƪU*���rm8�9P��}�m̛x�Y	r�9�O�R�,��7b�7����:���ۗ��|���dm�F��>���{�P.㸥�+�`v�3z6)*�>v�ݭ�=K,3����:���傉NY��s|TK�G���y+JR~�%M�6ZC�뗴�1z�5�0s�7�r%��7��>b��Ev�b	𷫩3�D��7�mhZ��$��&E�%�B� ��,Fx���ђ3�M$�p,�PN3]�h�b(c��V��L����։�s1�Χȵ���}�^�*JNE9KϝF��.lM�|�2g��`���;p�@y�B����@��G,w΂!���V�ny��(������CC��T��	#O�8&UN��:s��Z��'�;l�R�1�Yv3�2,i����Ab����PB}La��$����̆��Ia
��v�Al�߼6��)�u�3�%�_";�\�$��\F��G�V���,��>rєo�$�iҽ����j#܃�� S�1�/;Ny�d;f�e�f&�N0n�	�������/�V��ߧ��͈�����T������������].G﮷Q���0��f�w��i�v�r�B:��oC̶��i9}nS��;o#�0k�$Y�L��%H"�׈D�Ȣ������#��b�=���<���h���'I����3�d��ޠ$�&r0�L��M��u�g�����9?~��Jp��(7b!e��N���EK����T����)�V���Z�&�](^��S߳����>���@9�f�:�D,[�a<�Ŭ�B/�ٶ�L�J��s�=���ց�R��5�3�7�Dh�-ǲ}��է_���O�Z>Q�AQ����lzī���s���̨*���u�'���5gF��7��$��Vl0bs`����Z�bK�JtԜb�(�x1�[7t���<`ȟ�!��c�KMƼ�����sg�%�9o����C���iy}|ӫ�Ҩ��Bk��lIq1�jr��N�I���%�������ғ�eu	�ԐKΝ�靤���g�H��7�9#�̮2	F�S�hX,`�CȞ,�g��U
g��=EqhX���c���r����|�Kq��Xjuuu�� �(x�� �54ߪ���{Y8�{���d���j���;9�D_p{U�
�o�4d�x���ؼW��g��@�`�dC�P�PcqK�ρ�w�ಊ�����t�v�/���R��xl�$�xmQy�'���C�r
=�=�*�	Y�Q����f�� Π�w�N[�Pc�^��$�S��MWՆշ����7��o�::
7�r0�6	���ˊV!��(/ 5n�<����R��.���D�ކ��jY݃�������\P�I&!Zq/F�}�����҈s�,����g��e�~g{��v�ўu����sy�qm06\�Nl��.�@�~�^F5ߏ����I��H`%d�{��qnh8�`��=J�v�Q���o��gx'MQ^�k#�������g���S"/Ci�K�i�|Ts���D���f��%r�Ѕq��򝮦�,LhW��֨G/-�ֲ5����J؁#�!^��o ALy�W���l�����ó��Hf5�?�BU� ���60�[�����i%�N�l4�%����U���xh"��ǎ�|\����I�T��.��1�?H+Σ�cVvUG߹�9�@����=��z��0�����<9ZKDn�9�S7��>�ju>�Z;?pӦMe��Y�<��0��P�0�(������Ͱ��W<�Jvϩ
���oFo,��jD���`����r���2F�[gVHPP�KCU����z?�m�f�=5M�z{�z`AĻN�u����v��{d�n���&Ű���+lAv�S:��y%��(檻�D��@���B��BC�`'x���:� @����v� �^UX8�+�-�#��ذA]f�O�}��O��+��NO[HB,Snx�y]����v��E����c��z��!o\̼�Wv/�=�Bne<���HDzNq�����N�\�E������.�����S����7�[�])[)b���s܏�j~�Q/��Y9��3��9�~������XnKNr��>I�����<K����l���t�b���$-�I����
_���YJ�RǅF	���AdD����Q����m��W Y+� !:������~Ո���Ndɱ�]j�̬ғ��M��{l���-�?���L���jT���iV�QyW�����o��9�~�魉��!j�҈pOU�{c0)�-���<�ɓ'����Z9z���́���r,��\��ķ�zF�-az�Gd#����}�.�rd�9�S�N���W�;����/��x0z�YH�SBv~����	���@��*^� P��\���u�>�����#�:���j��vg��1����J�.�T*0>n�EI�����	�ռ���?�2�J\;w��6nc�{V�������p��1�v��1+f��$�"��&(�t��g��u�)d�1�i��`��SI��0?�Jl0��>/��Ea� ���x�?�m�(��L�|�K�)���{V=�t\�U��W'a;�P:Hݹ�O��������&F㮢Y�;�;�� 8D�e{����Z��j*��Uzpo��*%�}޴I` Ǘ�����=)t�y�BU��O��9�p���B�~��/�=�=�Oڟ�������[O�L��l0����q�wj���1�~	���:����lx��������;�����ŗ�s��d�O��_�1(JIB��b�O���c����M���V��n�l��Ґ�I!��4͊��Ag#�u�׻�)G]I3Mb�r��Ǽ���]��)��-�����龙�E�OY	t���?�k~����
��[����^��%�Ǭ�\jr%ֶ�؄m��'sB�П�{��18����'��*6��w���]��:D�	I�3rW�X��m��s����d����V�P����斺s^i��aC���ȹ��/w{T�t+�Q9)��¸��~�쿩��8�8q��uS$�yO^�9�D��)�׻n�C!�&��l�m��o}l*=��Q��p���)9��Dz'w5�x�ɘ�Fv��,�0M�zZmx��o���ۢ�x5A���o�Q����?�Y$Q҄��͓���\n�e�߲�w�e������DF� �C���WSL�y����~�o��o碰޷l�l����������]����A&��%�*���S�K���fQ��.���ŦMȕ�R�;��>�p����w+F3����k�B�"iD ׏�d��U�w���W�y���E�~ӝu+�X'�#;�R��/�OR,S��\�T[��Y �S�~�?!��I�RX>��a��D���D����@UR��+��a����k��粅}ļm_�yh<R2�Y�%�N���_�;�n�l�߸��Ŋ�w<+�u�b���W�>��ۏ�c�^��kyNY�9��ԿÚP�\mX��`��?���^&zԮ�'���]�Ʒi��_�&���r	���Z�� �ɈW��٪���߭���&_o�rd�z$<	���1+3�Nc�v�{��9)	�)���ǃ�g([hs��Z�k��x�ӏkm_���7���m��|��v{5�UP����:4��yy]"�pEx;�X�Py��rC���bNi�h��<&�<�D�?�.��;|%��_��{8r��/ZY[ �t�{��Y�7�jk�[NL��W��eDC�>E��YƟ(
�Y����z��?��ť�v}�ȿ���*X������3��hm%]��/�%`�P��$��|1&D��(������"j�V�)y�m/t���^��:�����7��g	j�֙e�4�Ջ2E�������{��H�1��\K׶�^1����+a�� �f �����|��5�~Śߑ������#1.����[�� x R���]���ъ
��w����_q�\��aٛD0��ړ�3f��@_�b�җ�  �:�W<����աg<fq�|F�7a�勲� I�pX���*6��T�?Dn�AȌ���
��g�/�}KPF�$p�o|�9�EX�U �l�L�&���o&��be̍v��
�r��!}�C�tެ��Y�n�i���w_�����2�c�htRu�D�\��o��/�"]�	_�Ԗ{��GA\��Ca��� ��m�'ߙ*������`3�)DWl�lR�0�}z��b�����e�1 �Mn�?m�gF\!��_`�or����5L�����_�7��zFq�ػ-�E�:rQ�|1R7Y�T2�}����a>�������������~�z<v/Ť��+Uk�C��2��?Д\d>���v��i�$�"}]�n���S7k)����%��c�ʡ�Aw�o`�*.aF�Тܒ�X|��O��޷�,(��-p#?AϚ�*������!�_�^?�x�#n a�5m��<x�Zk�	kň����I&�&&&w�v�I&�f��)�&��}ͅo>~�?wڤci��h&[�6���HL,�����9^�A�ŝ6��ًo�Ǜh��ęg�.�_�����	U��J�v|92���3�ׯ_��q���N�Yصk��携�젧9�ǝ��_��	J�`6ٟDb
b� 	MdK�YZ�ZH�~LAY�!7��A`�b
��wuw;6/;wF������\+�P*|��Mu��իW?zt�j))���� W=b�Zz��H�������BY�Q����~�z�W;��u�T^���3?>UY�n���#�j��9&���ĵ�x���,j=�}̼	�7p� <BF.ZF���+@D� nW��#G4�ϟ�!?D����(<&�`�j�vjń�!���^������ݴu��Cd���|����KUpo�%g.W��n8f,9�a�{��W���ٟ�?�7�Z����CF� Ba�q����a�j���c$�k���I&'�Y�}L��,��O��8X�����SU��T/���s0w��p8E���ÙX�f�+��ơ(i=��fFuͅ�r�vvz��l9''�qv��UQ�"��Cd��0�_Qq��>��S��w����,�NF�z�m-f�|��e؆5�KHNF���}M�w��������������+�8�gddd^N{�z�LA?���ǢSN`�:���+������zz��S�ڝ���ݻ�~ih��w����I^~�]���a�Vo��DÄ7����Y)x�y5�>��NQ�b���?���ԥ��RE�q��m韃��=E2E�gյ?U��!�R���Y9:"C�����n�޺.C~����J��'zzz�L�_o�:�W���u����P��[o.��AS�K�'�;fD�݋�o��o������M���%��7��r�M��v���rؾ�1W-��v���}x�tYyy�M**내V��*|���W��?��-<����s�����g()��� ��S�f�!��$%������,�]!`+�ֱ����#UW�仞?ZZ{��ZC�h|��]s*9��oCC3��h�3����#_��� ���%�� 1%d�)����ǖm'^C���O脻��̥�+�H��;qv��H@Ӥw�dH�Z�
q	��p����E�G:UUA}3)��͛W'�|ӑ�-k��uކ�̥8x����;��j*���Z5�����0��R\R����>�c��ݬ7���6o^�Ve�sx����������L��E�I�C���ȃb�a13���Qp{a�O�_�[�)/�Ri}{�7�Α����7
[7k��&�F���iО2O\s��h���1�{�\���4�$�s��*����rZ-�����T/z�4$�b/��8U§�ԛ�a������C_Kܟ\���k$��q�R1�B��̮�b�L{�C�a���ޕ)<�od�`|��r�o�:�Z�[[��Ɲ�\H���w�)Vj}sm�&e�[�+������&ih��xx�`vY��nF�陳6u��: $Puʱ��[�{�/Qs7�g�k����Kg�����U@	��i�f�����F������>�&�y��	��� ׻�^W��h���Y#���ط�0�?4t�`��g���̮�)��N���7�����>�L?���n�A�N}��b{��g#�:�����9ͯ��V�GD��n�c&+U^^������#��<��1�W]��^��/�� /L���K2��ӂ,~'�� �J�l�@~��W����1ⶋ�9�Mv <������$�e8I�罸ZM�'/��6��TeuKK���L߅�ՓQ���Z����n��pk�����>��{��f��<$�U�d��kS��W����.c����O��2�m�+a��ۯG������1�G�3=y�a��C��={�Ν��Ŕ���w�`<����W���\x��	3V�V7X��V���[��}�#���>SB]f�S�?����EA���p����	��M���a�AFL��D��U�-o����
�7x��1kB{[0�����U�of C9�w���?��;@7���ܞ+��������Ϸ� V՚Ɩ��ucI�<[	�0 HB�����EQ)$��>�Dqyp�-1Y�g��ћ���#��[mS� T��z�S�]sYB���H�M]�����c��án��qWuE�R�JYs)k�
)BTD�Dd_�eƌ\-�W*���(�2H%Q��B��fb,��9d�u����s�~��u�}>s��>���z���C�J��i�?[��QϬ��^J���,.a=�MӚ�lz� �ނ=nhI���~Q2eE�+8�~ګ~�B����R�˰��=�!VIB��Tq�M�d�D2�Ǭg8[����9yKp2?J �h�Q�����r2ژ��:��n�v���+5\����j+(����m�!єa�ߝn ڐ���Uw�ݾ�Z%�1t�'����랢[�����c��ڋ<{�>�QɐE�<6�jX��d+;;��?�
(3m�K�x����\~��M���PVM����W�5�doyvxk�����R�Ԉ3��[:�1.��%y�5.��oW�	E�Ay���7���W��}~�`~�;7k����!\��!	jQW�|�#G���D2��ܣ� R���Z@�h�|	������:�t���y�s��y�X��%WRJ�p��9�9��+H�K�ȺߐuϝS��"	�'� �����<|��p�Ǉ�R���Q�H.�߇��<u0X��C��&@I�
5=Hm��jH��Q[���/�AF���|e��>�V�9Y���:1�3'�Ո��0���¬�AR�++���-PJm��<���F>d،��B��_���Ă_��-#��t��*.�!�L ڞ�0����;���2i��%��m���-*��r	���?�i�RQ
�H\�pLlS�ϑn�q��ź��1rEL�H@��j��������ɽ�2;i?��8{��:nq�~v��=�����{��a��q`��&q�����4��O�������bf�vxJ�R��]OŶ��,��4B>r�:ɤ�KO�$���q��̞���z�� �IT��7o�J"���4ӫ��2Jg���0@?w�T����J�*��.%�L &fc+=� x����Hi+�4�o�L������N��sX@�1���<Z�����2��S����B�ɻY�F�8��s[>��W�[�~5�{j�w��$>���I�ܰo|�ج�rF��[��[�P�Dq��������*��e��/�XS��D/N��B]��t���+�D\{�9Y�W�t2�t��Ą��1}+W	�k����mఏ�V���.�n���N�h�XgonffY:���69��FMwoj�-ܳ��O��Jۯ
Mo u=�<P�p��Gy���i&�B+w�*���U6_8�1n��U���8@���O�[o d����䪵e�ּ^`Bn�=G�s��Ӽ�eQgY��6a���aV@���sxj@��w.�+�G���������9b_��dO���������ڵ�>}�5=<7K ׳�U�ZH����� �D+��FDx\��G�X���S���9-H�gʊW/��#�#˦&�-r.oo��W��.ʹ��5H�
�7�����S#����>?�S[�v��G�v�r����&��&���	+Fa��=R� r4v�J�jjY �'Y��q�&�UB]��л�H/'D6����9�-6i�~I���n��L��\z��Ț���鑊ѡfi����.�1��,��j	X�be�;nWEHj%���_7���K=-�=�ȡ%۶:l�]������[G��sf�J���BCP�F��^�Mi��+[���Ç������!�~��3&�<J����	lY!az����:�u��GJ(�᷐Sկ<V
z�A����>���EhKA
p&�E�L��`���j��

�v���(�:t
�ŝ����+�
1���:�D�م�V&!h�џ LO��v�X^Ҳ�p$ 3���Syw�7���n�)�LZK谂���b �+..�V�'Towǃ�p$��yQV�X�*p�VK�R�.��pZ4
��IW��2}�U�k���ԀOw7�G�rF�'Z^pBR��O�y�
�T�#�ϝ��Q-ZO;��|8'��S!���<҇h���{[�"aI�^LB�]r^$��e���.G$�g4��ҁU#���!��ȂY�õ<�h�J�QCԔ��	�X����u���y��=*��G\;���h��j~����gϟ 8�D���ocb���[�1�W�čMM��)�xR��]��6�U?�@P͇Bl.0с]_�%�~��&��Z=E�3O:��Ԯ��cG�X�2Oػu���lq��xOXN�cJ��� ���f��J>l���ڐU��9�:{n�]�\�d�I���������WdP��Փv�=(��X�Xh��ћ:ɂ��gf�^Ļ���]DVAU�9@� (��<�>{&���o�$$$�m�vT�p\t��o�:񇹳P�����N3�>lHXTT4[q�'��"���%��@��M�w�0�T��S;�B�U!6 `j�p<�"�V����JN����r
�u!������9b��O�e[C��������p��֬Y3
>@2tu�����e�����0>��˔.G�^����c����Om�<�o���A!S�b����/6�:HVx�:=]���slo��7y(r?�,6j96Y� 	�d��~�	���#��=���Q�۟�GsJ�i�h;��>�[K~��V	��iW�.\��B��mn[\7=�:���{-ÔV����85�yGuu���8�J�N�"2J�4;��CN���@�«�t��3��V\㜅�ߤ���'�u�>N!ԁ�=o9
\��h��z�Y#1C�YI�ɨ�t�5��r(��e1&4���쨌����	o�!�d����䗆�DP"�h4�B��o�Qh{�GT�=1Hu��] r(�I33�ލ�������|���ݗ����ñG��ө����f���S���;�0m���}����7;C�t~�-|ں�rnĖ210M�mr��Sy�k����ݮ�ɨ��Դy�}Y�[Z��ft����\�*}�_w���K���q�}��'�WT-�4��a<�Z�]�q��<���%�J\�}3�؟=��]̧�s
T9���'�
�s�;ʄRÆ���Nz6� w��$E�N<�;���(*�f�*V��yAGK�c�l��*j�uΒ�ι��5��u���%
(�]V:[�x>��hkk�8'\SXQ_�v�=N5�������.�z#�*�fN�%ⴷ����C�r��v���������eio��?^Gmz�}�92ύqK���^~u�ho��hgbj�?���izf��_�}���P���d��9=�CY9����M �j���mV�;.�(�`��|��g�5T�ˏ�l�{ǼQS�"J�����ㅆ�ZrR�#iw����Us�cG{��]*~|@�`��PJ���:���F�E9�C�&�uޅ(��VQ#tۗt�V9�Z�)�\��C���̷��4�͔	���gCC%�L��c����E����`Mg��@�ț//��O����"�7P��b#��N�ww�JKi<����@n��̞B�A�ٻ4��W.��n��"���a�͐_��9���C��C�W[�K"�|���R�� -U 3{�)����1#����ֶ�^��{n�B��:�9Iu��|�ѵ*������_�]48�-|��AXuﻍ�l��ɾ'\�+��#`���ùdr�����ul��_{Fu}�蠬�0:����X�����dv{3���d!��63��|��ݳ��t���_�	�@X
G�8�5����� b2��/��?� ���YYaD�zѮq�̾Ч#��m�S���+_��[h�+\)2�[y��Cһo[�=$��{	����?����T��܄9���]�b|<{�_C�����)W}tm�Q�w�����rZ\%ַo߬,,�T��x�;]���)�*{�Fɭ�UHJU���-|t���Ŵ2���h�I$���Ŷ^��<�@V�'������~	P����ĽÏ Ђ�YB�|SQa9���y��H_ݘq�]�˭�s�@;U�O����l0�;3��[�2�,�z��^�MA�����
���������<9̨�y��k�I����N�g�@� ʽ������t͜����YM�P��<$���'�-��r�2����������Aw&?ޠYHO:��Y.��$�2;���l��s!Hq�5�g~��y޹�҈ TM��glw�Bz[:;X���	��w2�w����G��� ��	#��d�z���VxQ�8��S��{ �l>D�4����ɘ�@����J(����j!��������X˹pR�8�ڡ����{����\H8d�Lk��������Q���{�Gm|�6�j����j�'s�?�H-�˱>'�tn/=4X &G�f�D�@�bPs���nd��)�z�R<�9�)�OF�4�l�x]��J�ֻ�M����C[.G�۝ܴiS�5�8�����$�w�`�V���F����d(TϠĽ���K)�S�#����z�v�V��UA����ΓB2�L���ǒ>�����olT�wTx4ϗ���ւ9��jz4b��ɯ��)u�\�.�C�v1�A/Xh�A���L����11h�g�ubn��QK#��dv����"�۱K�H1�����"�G�1�KA`Ŭ���)�2@A4�5��5��Ќ��@ϓ��"�#\�����?9H$��9��TL���T�G��Q�:^@�D�V�d6�����7�gG#"'k��":73d3:K�EY�3wee��K��0��z�b�Q�]����}��W�7q�S�2]tT0��o�o������A9>���%?~C���#c�f��.��O����o|/neF'Cqs�}nR�#�?y�^���U��5Vg�
hl�w+;��t2R��D�?Z�g���&�2H��j����~�ռ:'C~������ٳɓ�,�Y�����?bi9����쫫w�D��e?�����Ȋ��k����x{�с�O4O�}�����&�\n;:b��aV����c#/|��&<�J�iW�
��E��nX��w���Y�{�:�Ǣ��d��3���������K��?xE�+n�z˄���p]JJ�=<<�}���I��@t]�}�(�	ƧN]��J���i��h� �-����9Jۅ,��T�D��w-��z�!*y�.����⦠�Y�A���75x�|zGf�}U�*�$
�f�jf��r������b����ܮ;�Rrr��$"�x��
�ڸ��c	f΃3jķC�b��n��4�:�o�Ϋ�!�<z3�Ջ��Y�W�y|BdD�w\���FC+%MC��9����j�|H�c� �.�]���k���|�2�Eέ�p��c�<���OvBH�O�2�޳g=�F�\����ؽ2����D(�
/�<����J��c��LՕ��&0J���d /��vR�����p��^%�YJm�K9�7Q6~"��b硺�P��]�kq�y��� &�:��1���>�s���D���\mE��k�I�ׯ�̣aqz`K���Rg^�nȕ�pq��XkZ�P�3���u������������?G������Tw��7�������uu�Y��;NM �_o	Oo^�+c�ș���w�^%&8���I�`F�r�t�����?$"�M�1��䜌j��Mٶǟ��v?�QN�V���.��`�!9�� �F���0���p*�!��Xb0
�z��k���|3���r�4���%��&X��������b޶��|i�y����V����O��-��a���l��Ȇ�ߞ����k���r�i/�nc=����O��n칁���!�%�.|\b�؇ �BԲ�'RO�a#��6 �Yk띃R
րc����^��
��}w��2��+�SUU�zy�J&!�y�ڣ�"�
��23kGpY��a�d��Sύ�����c���|R��]��"����QVz�l�V]�¢!���J��FLl����9Q=�y<yּ�� �2a~�yZ`����ϋ��KV"�}��$�I������_�ĕZ���b�9w���Za�7�H^	�R{E�tp{�`_���*�����UG ?�?Ux���Z����S&4��=���n�dW���r1�ަ�D���Ŷ|��IK�ù+-�*���<���ٯ�	�]f�ԡ,���jq��/���n\����!�tw�q]�	��^?S�r�qŵj��'ͩ�<;u|�D)C��۽���==V��p�p�� ���v��>_֘����8���Խ�k����Qn���R3ۜ�FЙ~�\\M&6Դ�RJ��	v�ڠ��3��n ��Y����23��N�nT��Q,�{�r��u�^75�
�$���Sy�l����g���3��ź�����6��m�W�����W޻W�n�I;w����H 0�a�Zi��ګ>eJ���+�1��C��qv�6�u��R®�eS]������_�-�RR����ZB��{�>p[�p��Դ�Z뤑O�F���ovw����7w�O������F����ּ��QR��r�*�<+��bF����?.�Bއ�\�2�E6�Z�W�� {�̰ צM_U���Yp��(�>���x�;���}��8����y4�ת���fF
KI��z:��Vޝ�&\�-�;�� �k �Y��uF�����h
� V*�޲=^W�!�;ʶ��n��gP�KȜ���b��6�6qӼ�<�N=���x߷o���{n�_%-_�\xƻ���ZU(U��'3bg��Naam0�77��Z��	%�@������\~T����tpF����h��L�>q%`ډJX�ރ� O���9��&r�S��̕��/�&K�nnSp��T2�-���E���C��	�oj�_ݡKE�S�4��$J��o���uFa϶�;��+������7��,đ������aaa��*�uaPr+�� ��D/][��)Ҹ��.`��;�P�����i�F�̃�*Ο��X������Z�	�	޸�=� �]/!�fb�W�Ac�t7_$���-�)���tחv�:u��wX L�a���[՘�����ҵ;D�Z�P먗)?��[!Lv��B���}o޼I�OI����"]�!���,]���3k����5;�ZՈ�;R.�ps�l�H��.��� {�ݼ�eݦ�-<�uWH
Ϭ���[R�D)@L@����[��v���G�IQ��[h��(�����5	zX�EK5���s[��N@y�ETRQw,��|��x��3G���!� ��WP������1w��c7��w>�M������bM�$�NI�d7�m�8 �s>��f�z�f���l��,�x�s� �,�+�G�j��1�欨����{Sjq	��G�����ul����*Iǎ+��ٳd,&M�Rn������a6J���%���bn&�8V��˃��n�������&>������T�|�ҟMש��EM���C������p��)��~�����W�N�h�uq��#/�CN9��J-|Z����������jC��L�\��.�;U��fA�}ܪe�<�wz0@=&�m��_i�M�/<���7�c�Wx��2��r��7&6���
E7qqaKRO���^ęW��b׶V���m/��3��ZP�=(Le��� %>>��*�� {����]Ԯ楶�HFM�dnW�����Oy$��C2=M����>(�pǟ������0�a���N��9�����fW������J�����aJ��,5īg�O������@�8\�Cv ��_�b()?L�|����Z�g'��ĭ�Fu�U���xԸ���P�h,����x�;n���m͗�����g�/h���nQU�����>u���4c��1dV^d?�(��Ay�o�`Zj`�E�_��~
g�[A�QG��#jH��T�����B����� ���o����yl6��U���fN�Yy�h?�N0�ڒӷ],�q�(��[FJ�����"��(���� �L��L�Tc'F��WIdn��:W�uq�q�Ë��5����w \N0HE�\�n��0�1�۫�~�J��Q&n�t�,^m{S{5��Ü���{�;��kjl��<�V�1����Q�wkv�ð��ō� J�l�2Xw���@�^=C��J�I�����a�Z����$��
R�c���#�FT=\�[�}{�����-ʪV�q�?I�@G]5���xj?������߾}�7)l笛��|3�w9�d�v��Y�~����S�MR
i�s1S	��uӍ�ڑJ\�}�QX�Hr^Vt&!oª���x-
ΦM�p�G�{��~zLh�`l"`=��lT�0��[#mb#'X�!�R:X����0����I^�����l����qxL�e4��!����>u]f��*�|}�����l4�Â��f*��%��QG��my�qe1&-E�������4��X����S�۶G�D�Bc|ܽ����<�	�tn�_��i�-��.��%�F�"����(�(P�H��-`6��z�>�-X_k������6�5����mUR�}Ѿ��5���2�1�R�k����l_zwb��*S�l��n98E�:��[q�G�r���d�N�K�4?9]|	�+ڳ���#vv,.�
tX�2�]�_fK�`Z䱎b�mYU ��������q�t�Z5@
��YY	�yh��7~KV��7L!N���}}��̫���5��c�gx�/
:y�#����/w��t�L___ﹷk���y�8�j�D��4��eْ��?S�t��IL4�b�Q=�����V�޷D"�\��N~�4���^��v�8���K�峗4u� �m��4dѪ+�����w�G{C�i�KYhP=(���7	4?���:88�Վ�[��0D�}w�g�ͣsFAª�^k9w�K���Bb�n�����ag�b��|.��Lw��f��"����z$�,�H�"�e3L9�IjG�}g'i�|���%�rPJ���|%�"��֠sq�s� c�R���j�􆑈w�s(u%�FECϫ����x�ll�H>U�u�������X��6�ڵ�ť���&Ψ7���{�5���J�O �ߔ�3N�<��&7Qw-�cu�c�!�$66��A3J!`�������;�_LӃ�I��X�n��$n@�;X�C%�_	A�>�Jm�9z�M|.��bpHȝ
�i��KnL�?"��n�c\%{,�<�FL�������LK5�e�f��
��sއ�6�AKrӑ�=fݺ�=���qwD�Hn��nl��g�Z���*�␼%�v�wf�~.�T�G�$����ۍ��+ށp��<���*�1�I�EKY{$�׽Q;�ck�����L��@,x�b�NI��[� ����5;��R�O�I\%%�ϪE���;�6�ߘ��dC�S����Q�S����!	:\��+��4p�<8�3jYT\
Gɹc$��JA5�'�O9y��\���4����֮��W޿_�N7�:C�HH2���vP�eߍG#<�]:�I4����/Y{O��U|�YWE�c�!�:W%-	,��v4{_�m�HSG'lI����Z�~ʫo�Q)-XY;���,H��5��On�uy����6
��N\9§�6.:��{�ܰ=�z
��ql)��vG�U�o�ɦ<��1ו�ڸ7��]�
r�߱5����g��~�(���㚬U��^P��~��>��+ <������������T��[FF"w�>I}(]�_:|Ƣ`�D>�,9�&�7Q? �4Ϻ�f���V�$\%LbpW
E���Z��@ܬm��9�*�͛7_g���ҵ����sߔvԕ"l |�V�fi����W�j��������.|D��s5���,a�_�"�n�rh��PL};g�7���st�����[���Ԉ��'cVkd�o�4 �;|f���M�i������ ��"��<ǝ<АR�S���֗�xh�n�	�>���l"v֣�6�����[d����D��.5��̘�޹�����$��HUy��Q������3�q݃9O8��kr�)���b��U��gʰ� ��Lm�_wh=EQ���:��Oƾ"��-�r�x����Q
�J~�9�މ��w��REbvS��/���^7�Ng���1=s��H�e퉧BY�]�z..��J Շ<V��#��_�U�����	�:J��Zp%pO��D��΢f�#Ik���D��Q�(m��㦭`��ٙ�]_��i�h��@
�U.G)hXJA�IGqt��f�I��>t 8ؐ�%\�2�1'��g���j�A��S�|'|�P[6Q�h�Z��V/]s+؆�X)���BMH�t�b�Q��L�Q���t\�gE�z\L���r�9�[N��L�?4
?�c"~:�UC�i������ooԅ�#�]�w4�_�O�O�;��b��T=5-�:5�$Y"W��r�f���j�(��'}v�B��t���찟T�fG#*�Uf���Ӳ���L||BDǱF�B���P�$&�~Dn���$����P������	����7���|�F��h��c�F�D��c��NAl>]�Q7�%�D�ϯ?˘�ף�pk�|��i��]�嘒M�&�uE�Eužg�Y/��A���ě��bbb�r���}hJC5hV"���b��sP��L���*n��w�Ϗ�^H�d�<)8�S�.��/Ɉ�Ӏv���Y��,�Uz�챌ª �y���P����_�?TA��d�dqWe��1�^Gg�������¯�w����~'�qtbg��1;g�oGh���\?66�BB�A�<q�'T�m�C)�s3)%"��<F\�Zm��)�����c>WC�O|
<����]�����,����t-�;���|_txKl�~�v�?{	L�i���ƾ��_~�Vf���� B�[���?�����y(�@˱F'[�J�}I���x�А:�n�ho�n7�VB��������TtNWw�Ӓ��>[!9�YG+�O��D�2N7d13�Q-ز��ԟ���s&�&E9��|�й������W�ª��L�Ѻ���:T�&���V�z����:g�$���5n�+�n~����^Qי�F�ꘓJc�5��OEP���֯���!�+_������HJ`�+�B�r�써h�%��8�襜�o���~����Q�=.:���LN����F�)?��T�P�h\�sa�# �$Y�n3jKc�GV�͈��n|f�v��i��T�T<���!����Ց�%�dbk�;��C���b�˰����0>��L1��ЖFc�j�vߑ �W6*�f�=�o�8�Z�u���*:,�ڻ���Xbl��R�{}���,Z�(�?((����l����qb�_K
�,��A5��ss(lE��,�B~XV�Nq�����!�Nޯ�ޚ�1��UOff�����L;��3S�Ae���)�ha	�4�n4�BTՋ�ꌣml���"7R!j�_��S���M���<M;m���:�ݤ#��v��AO=�辨��u%۫��Yy%�#A���y��k����nX����M�3K�F
�t��K���%ܺ_YZ��WK�:�b`��� ��y��c���P�J�LB5?M��Y-ۅ\j�!�?~�u�'��8�2��Q�]�t�W��s���BSJI�[��77�>L%{���57h�z�zR����7:C�m�/������}wͶHb>�1[wk�o�B|�wW����v���k�Ν:rM�J\mD�7{%�����0������a�)��R?z����M\_otH��N>!"�Ο����MW�d{���>G-��FG��"�q*
�^^rf����gI�o:XГ�[_Df��UmkPҨ�;qTG�c(�:�k���K������S�X���
�݋�!~�e �2ԝ��s�Ƒ�M�SG&Z���Z��%�g)�DƩp IΥ�@8�i{P���^��f#L=�:�R����W�Vw���pt�r�퇋bߴ&���8�s.9$y�N�ڵk__K�]����D���!ž7��F-^�;��z��E�X,) ����8��S阘9_��}2s��۾� T.M;kl������Q����7�h���KZ=.?�q�ϭ-C�:݃�{�4�!�d�g'.�I��Z׏�\���MzA�o����޵%�+K�A^��'Զ6�6<�8��u*��5�Q���OXqf�sDa:�1e��`����WF(�\����è=�������f>�4#3�y�:J��7O(Q?�x�2u�+�W��*�qUJN��~������Y���H�[R^��V�[��k�����@K�$q ���9K*0��:!���摒�r̎e�c�jqۓ��-�ܞ��r2��֮����N�e:�گ}�(��ǜ���Ҡ��M{Hh�ɾ8�l��WD:��.�j�Zb�H���(P�4cX:u�3����녜{����M9�����k�E	��ϟ^�����3!�a��({h��A0����ؑ�a/��k�b$<<|����(pzvx۠3kk��g^�2����?��tO�Մ�}P�\�r%|�M��SeR�Be�(���6߹���6Rާ�yVd,��p!�Cr�e�SS��G�^{�J>E�Ѯ0���N�ϲ<�a�Ϭ���
�T)�_[0^ w���*��=�*��:�x�#B�VG�V��g;Kp�<�;� Gm���h��k>�;Y=b���й�ZG���%��6�����?+T��<y1��'Ȥ��*��RH!,�����K�B�*:��u���6q�_��۩��|4�e[o\w������|J�Q�O�c�\l*�.	���B(<���An0-��Y2�@�~�Ź�vΎ���F��?���-+Bcj��������M�V����TQ����ME��(����7�~��]՛�w˹�cT�K'� ��ի��2�V�O [�˄�+��ߜ�o;pM����WF;����A$����ڃ/�|�P���\L��L�	yN�m<��S�'�e#P�����V�Ѥ.^W�9���㧰6��V��Jg�� ��ʧ�M#�7�����������mɱ��G�u����������+.3f����G���j!�g��v�����\�n�'��~c�n����y���!:� �&(%%�^T�����$�b}�٢F�Z665�t� ��w4�D�����H>�ٳg�o���������K:�yl.�������zF}����O��":�~J�җcU�雖/_�'a	�]@���?��C9�J)��}0���9Ǜ�O��{�TXZ�f�k
{�m?�V��lv�� ��w���{��P����5m��K=!���y������Y��3�:����R��󨓴~Fd��an��{Ҝ5�N���$�7>���������X#�����]KEݚJ b�=�r�SnvH�vӜo��Ȣn�SÇd���Ә�Zß�&ݮ�g�db�2��� ϳ��:�@��R��y�&ř�(�9#�zO�2ݜ����ݜ�(ތXG�}�rS��a+��*�����Cz[�=f��V�	�Jڳ�~�YA¥]��VV���w��5���J�Z��xg�Q|�i��T���H���턽�aR�T�����7OeDV><E�6�}���S(�`�2τS�@�mE�ij�3��a�|�:$ں#�)`���q.�n
�ڻ�c#�4d=��7BC�5��xWϚeBt�2�vj�T��ʽ��s�.6G�U)�3�Q ��b"v��Ň�G�:='�Ջ����%�	��M�Q�s��B�OW�~�Z橣��� u+I;
���X��V��>%o�;��ڒv��L���.6�P(D�ӧ{;�'�������GG�X�W��>��;9z��� �7���gǌ�v\9��K�LL����+H�i��o�QJ�kYv�;��iO�w�'��A� oI�ۗ3n��e����:7Z(:D�Ŭ��W޳g}��c �Ҍpt��@���3ڐ���s|�,�:ِ��/7�����W
�}��E	?�,�C�bBw/H�� ˺�J�G�^!�z/�Txz�F<����#]`ް���0�Y�d��$iiiGB)RqH�nx�^�Jr��<��gΞ�@͊����
ɟ�/���w,9;��ҧk�l��;w�urr��ۈ�3��dq���g������uUp6Y�|ty�R�����gf�<5?(��ky6�����uhֿ��^QQa	�s��0����H���9�"�b����%ps���Cg�}G�@!����0<���lgϟ�7L/�)+/?؆����L�uD�
r�p���>���^()l���F��d
��<�7�~�X��y��|��yk����\HO!�u򎍍���u:VLL���J�J$n=5�}��Av-�ꮸ9����и�nF����5��������.쨾����TAv�T�4���W�o�w��.5�j��s���~%i݂$�� �΂Q��p���0$�PSG�^g�!��$���pmoEZK���.�g�m��m�6fm�Bz��7>�~��Q���@�% ��_�=����[N�����2^�V�v��SUU��<���A�)Z7�B�V�@�̶|Y��#��T)�6é	��� �)Aļ��^����(�ηm[0�N�_B��̘Vz��o������Ԃ�W�k%~�GL��@��H��a����������`DRRR�YFEy�?�	.ɗ�փ�������jN�(��˗R��on��-�YV�A���ו{N�zI���yѬ���ԡ˂:\��u������B�qTҟ�.����Q1�Qp��H4U1�`brGZPm긁YܔơCg���T���� �I��_6oJc�)!�kV'�6^�E��#��6�+��&�_�(� _B�\Zn�� �(�`���}j�K�G���U��*b����:��>8���sq��M���@���uJ��t���c,~�С�y����*2��-��{���w�NK�BI����l���p��BQ�xO&a����%#����;�v7w��%u�%�YZ�ݸ��&��M+�Z^^~�Q��R�t��[�Q�n~�P�~�p9���P�=�1�"�sxP�ߢ��m�j1̮���̶\YΝ�z-�:&1��XL� �{�\\9���S�~y[�(5pi熩8��&���44��� fjV16���A�,��?��a��<<!_�|I�h���b0�A�����kj�w�}ā���}�l'�b�`��Ԝ�qn�vC]� �9@�9c�-�gp�߹y��%�zzڧ� ���VЙ_��읰+��ۏ�m?6���B�@)��(Y�بӏZ����%^XA�_H�v���۽��V'�W�Ӆ���&��^Fٹ
eeeG��T)�RZFٴj��ү��B/� ��UN&q��A:�-��B]�1>�t�/,]Z�c���i�
][���+�Q�,,g�n�Sn��d���t^���W���#�2i�7R3G��=R����/`�EaeS��di+R��Ϛb9�w��4p^6��P���r�C�h݋��J��2���&ͧ)~Xͅ�@�<2=vb^����`��v:9pbn���&-0�LS�n�߿� E�Bw�];i�R��}�d��cSN���s�^}%Fl�6��4�Loȧ���8
�d�w~?l{a�L<��y�ȭ )i�r��~}�4�A��+{>En�$�8Hy��uZ�⯒9%@3��.5�Ш��f�+��B�'��E�Y��T��+���ʒ���}��;hSΨv����r�ԫ��; 2��9��:��F�M�]K$9ڦ�͗Q���+�^��+�
� ��A��4i,mk�����;_!����2���0d���Т��`C>W4xߪ����}'M��C��p<����Q]�5�c�`yB�[��q쿖gDWn^]�w��(?��n����0B��<���!�cU5z��d��ˠ�j�U���y
�י����y\o�pD&��,�U�F�ϦG4�>�Zp��Џ?n޲�}ѝ���W1F����B�������r���$�j3�@+ێ���\4����y,m����ķ.���{TYL.˼
0�¢G�_np-����������w�jYAB�F_��� �_AK���!�CV�����;��v��2�A����p��mXOs�U�N�ظ0��Y�D�D�߅/�)�9�P2�����Ɔ^�z5McQ�{��]B�� �XX���C���y�`(HWv9�'6/:����#�1����"���ѡB�[n?��K������p�e����t6��|����Lm�t�A��v��ST:�4B�翔������/9ܞ����b�RÜ,���ѿ���t9��᷻G,�n��'�.K?��jҹ�8.�xu��~�yA���vs.��+My<�B.�7�N�z���v���Ͳ��Kt�C;�i����sj���U�Qbtg�t:���j��)��Vq�KD�]�]:OD�nĴy����5=eb�?zb�◜�c�G�T士�=���k%֞ke<_���$���"���.�������.��2�~1ap�e���'Ht]Ѭҿ�O1����P�)f���EzZ�T�����T��������8�U�
Lmd/V?E�K�@b�����	f\�0���r�JX��ѯ!�:�j���0��.�q�2�~F�=0#&����0÷	�X.����U�3�3,2�q�u�=��x���K� ��W�nlg���3
3*1.2��3�ѳ'S���f���k�Z(r�"1�ta ���|UV�v)��%��s�>�*�,���\��bA�(��ۆf\v�\/,��e�}/��9c�b���_5��j!��Sn�C�V���2z-i�=�/���z�g��u�/+�}K�r���V��8��7]����g�/<cgx���]�'��`�f^7����b否�0s���˚ˊg�69#�����b�/���Z{��Jѿ��R1S貢�]-\&�m]K*�`<m���`��,aM�r/�O�?/x��ӿ|����-�l}h1Z.�ni�S���W��n�7�d�p�%}B9	K�cg���3Vxvօـa\?�D}�癋2�0kf�aMa�x�]V̔�k��6w�Ҿ���K���.֡t�en�Z���I�h��&�� $?���<�ѵm��|�6ʠ�R���-m~/���IK�.���3�g}ց���ZE�����=�o[,]ћ��܋|������_�����K�m�T,s]����L�C����t��r5]�G�;���q<�q�;`�^p�l�������f�J-�Qۇ.������Ӆ_�yI���K��[��k��,� y,w�J2�)�R��M*�/��`�.;�K|1��sY�,���=2�l�Z�'�Le�`B*L(��>a��sS��3t}�A���g;��΃���m�����4(��tY\ALcc�g�703��d�}�Ś�,,,����� ������PUT��?�����P�\��1�|����O�09�����.����g5V��d�i�Z�OB��-����-����-����-����W,ɲ��Y�����z�O��w��{�1��~�
�ʖo�?f#���[�o�����Z��S���� ��������-����-����?�#&�+�F��+����´�X��Z&��/x.5�?��V!��q'�c+��Ά�o�11[,Y���
�n*�h,T	��{$|��U���ޱ��z��|�.ےDl��?���rN&��ҘJ��l��D.��6+��	j�В$/��sd�%��7��23��;�"�c
���ma1+�w���q,/Y)�2��\ϸ����1nc�
F�\�_���"��-��E䕀'�Le�����L��-�ҋG߉��e�ϑ����������Ϗ=����XǓl�_��D؊������"��-��h�{�/�x�[���̲BEWWל{��at�97�Ѱ��H�ɯA�����~~O͐xt�c���<g�g�nnv'��B�ց��::�R������^_��ᝣl��{6�+�̵���T,�pW,��'��u��*��c9�(��0Lev/Y[�lV�"�saz�~hc�� k�4�5L��jd���0��d-
c��=6�6�+���y;��n͊��_O͞�������{{^����,ӫ�5�x��;�u�Yg��;���K����-+'�J�R�!!!'�1|�@o��[JpX�rrȩ��������MJy�݄��Y�ߍ����!��������q�0>_�w%n=�Xq	�Y�p�\l(��]3�D��JN�n�5/�OOK{dZ�1�7���#?ÃJvdTZ�Bں�A1�Y�7�v��K�FW��}���������Ƨm>�D��k�{`�ɮ���"n�Z�QeFZ����]j����ڰI���8g����I=pܽ�ݝ<�lp�h$�l�/՝�zIN����*����F*�>�aɼZM��V����y�!T��,WN���oq��da{�����5.�俬�ɞ�a.��"�O�(��(x�x��M��ZP�������>����Y�_�o���-j�C���2�����ﳖ$�Ą�c�]�,mqg]]�x�0'��_���%arx_�]>��Ŝ�Q�7V�jht���h����Um�3NC�� 	�LU��_��^�i������X�e��LL�����0�h���Di�,���.|���3���ljb����N���𣲈IH$=�Kj4�j3.�Ū����a�g�0���t�L9�kI���N]!��j[è�9W�#��1������Z]�/o۫�g�3�����,YZ5�̞�8sé��~f�1ƺ��Ə���<����B��v`zr���uC>�v�%����FJ��vf`X��]�1�[����{��^
�1��ˌ+.�\���e�aO��"ɐ%J�±�L��
�>A����]���;��/�EEE��J �VHBT)"VzQA@���  M��@("  MB�TM�$A����>�+���;�ޛ�3�{����g��Z�U��>��c�,lf�ど�{�q8WN�F����פ��Q���5�!qK:<��Q��>df��S{����n}�s|Q,<hN���\|ζ��5�ϊ�6y�H��n��C�̌��I����!�D��O�ڼNs���u��|qN1}T� Z8~�ڀ�ps�d_�E�}ƭ�9�L�(MAt?�m������OK���R��̮;�#�x���X5f\�9�b�v���u�r��h/�Hu"�v�`���۟�eqK;_��Ґ�	�+~�U�
5��z����Uz�-;eh�	***3�l2q'fW�"Z��\W�{�e �d�&Ց�C�544��h�;��dK�^����a������#���l������X�?���Q{�4ొ۷l�-��&�j\��D�hFn�WNf��؋W�I%Kv a��Y5e�++ǚ����^n�������ʀ�p$��r��ax�H*�����6�$����𙛛;..~m����c�����&��1�b �b��aaa�Q���щ�0'�e�#����
��V�=���S��ƅ.�8��H��2Z��PiJ�fQ`x��YjJ��!�����.��uh�Z��f:�wB_��)�c����,�.-̨��8�wnrӯ� Wjcc�\'��'I�	`R�J�:L�o����G�c;���ׯ��6ˉC��;���Ϟ9��|���lh�)�0��Z�;up�ɭ[��yV��ENM�0��{v�ݽ}[��=.-�c�	��Tmee%�N�����Ǭ�v�[q�4��l�ʝ��i�6��R�]�Y�[лG�"��J��fY��I
y2����!�ڵ��P�c�Q�h ��*�M"�n��&�� %���q�����M4����Q'��jMl�$7n���?ݒ�s3Y?:��:S!|&��\&����\]�Ki"���G�>~Tl�2�����엶]9FtĬ���F2�및�,�A���c�qPK���� |��%�fP����Sf���zNHC�M,Ź;1娇g,j��@h؏&�ӻ,��\�[��S�A�� ,S�>p-�6'��DI>w*�i�6� z��b�Z+�=?�NEQ@8 '<G@~�l�!}͹K�$��J�����]�(�����pK�6¾���\g����/1���Du8�#`X�]b �,�
lF;����6�Nc��ܯ�>�_*�A&A���p4���{@3���<C�kNP��>�mH�Ѣ�/�K�ǆפP�rm��6�XYY~���??�r~�UF;�f��3�ʦ��	�-<C�e�U2�kenJ������)����)�<
<�sD�a���fԮ ���������c� ,�ꕑ��q���ss��0]��� �/�45JV�g@J�Yc�v��ӫ�R8�3��ƻ���pE�~!ʠ���~(�{2�Z�*̥�NV����1l���M��)��]�r࢝Z��R��N&���q_sw��S��7o.Q:6�6�Ji7X)퐡����'�切�4�S�)�@OHH�B$j�GF�v��/@n��"��ju�.��%���@8ӥc�D���;��U��<�z��8"����L-,ِ�y6��g`of*[��|�� ė����Z������GK�����d�}ޤ�"ڊ`c���J���GK��^�n����aO���Q��ٚ� ~��nC�P���:��q���U��=h����&'l .7��&���L��K,��a0A#A�v�Omg�'A�qUʛ�)'k�F�� ��{���E��p�)E�"CK��&�P����*lԤ�~�2���@�Sz��Q�k�;�U�@K�j�8VG΃��r��s���E0r�v`��7O���\��ꚲ�di7�?Pʁ��`���O�*\6�*����e2�x�c&
��Y� ����*����L�1�iH@�S:_��:Ps�$+8j�����J��穧��8�l����M�Y>�2Y�p�ٹp���#��-:�@E����wg��~E����#a��m/n����O/�x��9Y�ʳb_le�Ϥ,�u���;\�x��ozU�[���������7���}+��̘����@��TuW�;\EUu���kRz�|��kN�q���F�|t�;�?Z��Y'
�/r1=3�mc�4<�S5U-މ�-Y��\�lP�N/i��#,,|�J�۷k7�f?5$��%�.���/N�O���F[@5$�����#��]��������::i�\�����:��` ��Z���/E�L�H}=�(�����.+H����)��9��~^�y���R�J�爍oi�U��;Oꤼc~V/�z������-6��z��i6��[�̞���:$O�J�ԣ#����0 �+D�ΡP��!)�uDb�X�Ɂ�س���M�ɫ�Z�����9kamt�%�n�_w\we-��g��W�k�x^nƍ��/g���Z�oU��^���Z��]�С~Z���}l��^��̅+ʭ*� J�QTvRP	~���m�~8�=[FQ(�T�S�f����R��ii�7�&�;�ٮ�\w��=���p�	�q΅�����6�gm��/7��eAh}��0���g*�F��eh�D9�AC[�.f�q����X�^�����g��<Zj.`Fげ��.�8��:G�a,f>�������%t���(e$��^��_:/o��T󯫻\��qK9].((��()l��Ɗ;F+g���,��	fH�'!���oR�����	Q���`8�+�v�3�C���l�[�({�����R��m�C�HZ�ڮW/żN:�-���� ��Ҋ�cO�x�GGF�޽� ..��/tUQQ1"GI��_�nw	')��n��CE��w4<��Ś���d��6DM�����4M��qo?�Ab}����"nd��#�n�sFR���QR��i�-r�-�ho�]���3�V\���SA3�9f\�n��ɏ���LMB��v�]�v�.�k��9}�n:�]5r3���N��^���I���������c�^�f
@u�4�l��G��_��Ĝ�%����]jg�G��'���\����YŒ#��:�'�9��B�vx���T���be�9R��ho���B+C;?ڛ
�ĳ�z����[ho^�NZe��+�]?��<�ia�Ww�-�u�&��o.�Fd 恜>�˙�b���p��̼�1��a\�������6������\`X!@����?���ڽ������mQߞ�b����<G�;=P��7k��,���h���"?�����~���CL0wYr6Y �6��w#�`��D?�!���m��oۢ�u��7q���������jjn���ၽ:��F�.]�����m�;[j��CM�{]�z�QZ�Z>G�5���#x�a�mz
�t�,�,�F]�gF·�I�݃��(���&V�&.� �-�������j�mx������g�ڈ��SSS9�T���4�;���[^�	���Hr	,]	�6A3�/�5���۲礧�6}�r�`M%*�lOy��>���F�[X�8��-��1��"UUU����)v,_���|g��t����"����eM������JB �	j��k2��FK��a2 ���)3+ĸ�8��	_�R̊ۄ����l+�1pp�:{`ic��ֶ3�l�:8��޺��@p"=Pu(P�@6��},�H̷M7Ebs�~�Yy+���* �?�~�������A�JZ�����@�Z�y{r@@ P�V�0�{�?+t����-Е+W����
41Lvn����# Ъ�m�e��60���w���i###mi��a8h	���p��b�:�]�5aC�R��E��Î�� lF���@�.7S�^�n��������$��U��w�`�4���8bz��Z�y�1W�R;���g�-�9�� H���IT'W������S�uc����q�!�������"�3�pX�<
l��9��d���\)M��
�&-5y�5��ɏ����R��>�!�T���X�X�?�w;Z↾��#��P���<�;�����k�.�V�G��2x���7�����H^��F{��J0�܇T�\�s,�̎Kq��3�6�~�FFR�5H��@�LWW+�����\����[{�\м9Ͻ9�s�*@�}wPՉ�J:K���"9X�:5=��f�L&D��v��e:��)Q�O�:ů�>�	��%�K���/�_¿�	���L8_|@��Y�����K#\��Yz[�<ǽ,��?�����O�=b��s�{{�^����C������=�8�pr�{�շYR�e�^�8�SMF��i��6�l��{eA5��<iA�T�e���>x�s�Hy��㿃��z~s-Yi	�Yvx��&�j���!��m�O׹�I'C�����hF�ű���7�l��8m׻(Iǟ�%�M��c�u����s��3��^�+�j���w��v.O��|^Y(��X�t��,U�	�(ɹ����^?����ɁzlGj�+in���~)6��[����H@��v�	J�Z�ꌢ�/�"��%*�n1}Lϋ߮$j>	@m�\BV�%-a��V"�,�����qn6�8�!��G�fZ�h�%��}F�8���/To��By�!Ӌ	OJ�+�7�<�8�N/D�m�#���;]:��+�Ul��*���Yp�Q��;��SW�1�q�-Z��(RaǪ-\'ܖg�d��w�N�m���Lō���L6���p�Ί�Pu��Jq�\�p�E��w��D�-M@���j�u[Y�7����d�Q �Yj�i�~.,����]s�l9�~��dȠ����oP�4�f�'�f����������\�B���n�4 X����uW]����>��[ˇ߸)
���U��\��V��)>Jp��IoN���s�n��߄%>�X"9!(��MKU�Z��sB�N{��d��Z�B2���I�)�nuu�8��B�Kv�${�	I�e���(�7�wO�5��b"�%'Q]�h��w�����Y٘"ϑ9:�����ֽ�K�\.��c�Itpc�J��般𳆲ҥ�?��(Κ#K���pF������ |��3*�>CG�O.��9���"Y���E(j�f�3�~t��������(}�=Q�4��t4����!�8���g�;|ź[����8{��t�E�sf�����}�����P
g�Gm�������<�ʂ��X�	-�Di���[kRh���udK�Dѣ�p��
���Q�സ���At�\@I��7nb\e�\kM6-������f�mԤB��Hw#:B��Ɉ�&+����+sN�C<�h&6R�$�ၾ����orD�LX�u���1t$�	g}��t�k*Qfi�f$�����4�_^���Gut����}�x��s�'�w^��j�t���\��̓Ϋ�%+�΃t�v8�^�Z��[j�r�����~#/'��,
J���N��!�����/t$EI���q;�<��[����H>�����/Y�<+�U>>��~i���+�TL��X�����d�9��Ɔ����$n��G���L8�dHr�M�;�l��b.����P��7Gad6�TJ�?���Q�����c._(�PB��3Ƣ�ua�a���kD�1(��'��z�����l�]\�4�5���;���#�#//_��T`��aNd�Hʙ#n�e��c����OʦϾ�r��	���]�,{��� �J���')�
���s� ӻ��_7�n|*DV*۳?����]�k��+�&�! rM���$��@�W���Rh�O�݉?��
x5z�қ��(�`Ei����?&���T�P�D!�rđ����N�{��4���ch��<Ԁ����*U�珡� ���&Et�"�D0+��#Az�ط��%pA���)�?��]*�#����Y�}t�t��協B����A���o�AR�Q:M`�鞣\��y9�.W�ߖK$/�_����Qw��yxD���c��s���Ӕl�e�,R��	Q��- i���&���6�Ku]�7���4y�$_J�dw�B2�H{`(���G֓ ��K)tȪh��8���H����8#��� lXȅ�%�6�7���o#�WG@W��m�gu�mAJ��XVG��QQ��:�(���l����Y�G[HP���y���,8{OJ��H�6�2S�ML�K���^ʵ�OAk�I��갤��m0�
}�E2ӐM��SK��E!�H^�(��f�}�j�P|Q?��{y��]*��j���&�4�!x�/�E�w�%�"�
��.���U��h��l���P�-2<���$�oNUK�_T-1���Ѳ"��%V�/%r.�d�<@���ƽ�	�IX"5I+����5r���x�6BVU�	��\�I�&	P&�:v���H�yJBV�n��Ra�:~U�f\�o���k����!�=$��-�}A���/<��R -�Ց @C9B|�:��^��z�����*�_;0��mp�*U��Uu��q&�ʺ���KG���N��j��R�lR@ ���A4�4(2��� :��¯ݧY 	Q�]*�)��?
#�XJ}>�z��Y@�	�]Pu�o �=��ʯ �eZ��dQ<w�y�n`����A�k���	�hy��d��Ҩ[�����J��y�h�As)��L�$aClHT��~ع�'^j���*�]9�@謤�q�z�:�<T�S���3��~�IG�%�Y�6��{8l�U&��lC���:�fJ���)W�ZGg,���U�>�[��~K���yZ[	y����xD�/'�$����9��p�b3�_o�6<���u����Y"�B��
�~��Bc��
�"Z�!4����3~r���ʐ�����c����^Ū�tV�9׬?"�at��� ӧ�jgٷ#3\�s�J�nX�,��f�K���(���4��p*
�j�ي 9NMB3�ٛ�=��ܮ ��SU��{W�2����%�9䁒t8%�'N��[�_?Ȟ�%bx��/J�P1z��< Uxm�Z�����X���_LdE�Ʃ�n~V};/�nO��{ �5���B���r	'�,%��k���8Tr���pe�i�󼒓�5*l�K�<�3kG!ϙ��,��N���9gn[�*�\����u?8�+��H��L쓔S��sj�#��i��Pf�y�d����uh��҆[��D���Uc{=G.�y������Lv4�^p���_���-�Od��.�T����6��s��a��{ف������vڑ*��^�e�ʠ�Θ�up���hR��b��U=Duc�o�񈭼6���[��ߤ�R�o���t���W���+���b;7P#�,�j�ky���A�/j-i�_n�5������`���ʎ���	w~�,����[;&�O�ͭ�h	��7������F�m���\��dgΑϥ#ƞ�$[n����]�'�ʐ��%b&���|�"1[�1�ve��o��n�dL�V���������<���n�"�/���Λ��ya��q��r�)�R:Bl'Pz��=���w�]�2U%��g)�{tZ�͓:l���nO\���a�Ϸ���{A�r�#�� ���V1�`�UЌ&J��A
�˕+&�mv-,I��[��nܾ��;�Sa����(9���dU�G8���pl�E���$�����{����Y_.f4" %r��O�� �C����}�;��F���s6�C�Y�'���Tl�p+�I�����1�����g3u��"z��Ny���i�%��|�.�Ew���h	�L�M�|6������~�׌&�|C!���?�W>��C曟��U��5[�S�x�5gS� �FDȦ��BE�S�&0�%��=D�ﾞf����C�I�"��;J���;�DTU�X������3�=��:�����=GdU6�w�x�N����9wV�o�y�4i*5���b���Q}�E��܌��
]�t�@���UĿ�o�- d��4O��g�#U�>��|�v1۩I�V`���������*��>ݢ�.#Z���/���@�꿚�]��� ��Nnf��>�d�q
~ ��_�J��s<b"���z�J�7	��P�Oأ��:uχ�y(h3���n�og��p�=�����Ǌ	�4�-��)�jfʟ)��+�
��7�lô���c�_}�^��g2�7��d{�گ^���j�3�����g��(�_9�%�-q|�JPM*���8�戝%k����~�%�4 �$0� },��h��Y�şOK�;�H��N���m��eXs1E�*��>`29P7[)^�~z�b�p"W�&�	�i�`�7� cw �l{vL<,D���w��'�'�o�����@hېjc�@��F�ʥv���M���ǘ�Eop��lc�,9EKܠ�a��?�5OM�J��Tj��{�vU`IX�{�i�L+ã@<�+
6�.�8	Vd\�i��ԥ��h˺�o#2�2�K(l����	���,ˠf��,g��^�����R�����T.Z��G�����p�sߧw�ݡ�|t��
C.57L�Q�߇�9���#��D�_[�n��	1o�e\�/s˸�� ��23��	l��F�b�Ri���k�e>���j����6?��C�>�����_¿�	��%�K���/�_���	�7Q���Ф
��x���Y��Ǔr�ْc1�n+�SlkD�����e���7٫s���I�����jM�_�}D#�?:KNiJ��x��qv��h�����țO������a���,���_2���m:" ���%�Z1M�;�"�͇���F�D3�Y_��3ȦӁ���gi��Mu�`��E�U��hh*��ԁ���bܦ�H�/pb0|�T��dջמ\ng��Ùsݽ��������Pl�(V��v���u��}�6y��0ف�a�ӯ�r�>���R��$���^���XN �28 N~�8�C�/��T�k��Q *�(�5�Z��BHc���P��u@������͖��^�`�V �%�� H3�=�۷���[u�����A+����-v���|����/�ȭIx���0C�+�x���uz�������:�c@�Va�Hs}��74��!�>q �J&�V�V�+��o\���>�"�Q���7��"��5Qb���
��]�k�S-�$�����d��Z�k��;����1`�e������.�W��c�Z�ti �Y�5��"@,�m�����Za����jʕ�}T�! 7��P�%544��&�B	���:i\$ o_�k`��g���s��uՐ�V4z��ݙ5�F�uK���u���� 8�ϭ�m� k�����˿`��x��������5$P(ּM�}`�u�4V�~@ɿgMF^/ M	���}�ݏ�E��r�\g��,\����\f�0`"�.� dJ��7��c#TL�UR������%;
��=�{���D�2 ��)v<F�q �lYwp�E0���j]�g�3Q�X���g�>N>[�*@��G�$�{��ׯ7$$%���;�U[���l���7@�ZO�z? 8eBh��u��\Z@.n�5���D4�5�C�Wa�O�ɒ`�HE#���T$+ p� �+��q��p,Z�5ܫ6Nu10%4k\M	]ӛJl=�. ��C{�=���CO?Y��X� ���]��P��`x��G�D ��-�i�ϭ�� $ǁ�w�7P�gL���"O�C.�,4;�Q]�|��a^g���*�w�z3qîgJB���0F�Qk�J�}��N�H���o��?���د!=(t騴J�a���-�%�K��lE"��}N��a|��qMg��P|\���Z��ޑМ��[;"nd�3���M�����O�������s�Q��B��
��Q<���Rɿ�2���/ÿ��1��?B�^�ߘgH@/ؒ����[k{;V�<� U����z?��H��v�LNMM�,#2�h�U^��7b��ƙʐ����_�0,������ʲtrBb�@�-��xxj�� ���@�n^I	OKK˪C�=����� ��~�3)�,T��_\��?I߿�3���
v�JJJ���佪�-##���d��R'��!7*:����������Ia�M�R�(�K�)=H�����f��5�~�&��K>�]hl��֒D�˂�4=��3EhA|��`û�������;�s3$����,*<'����D��2����3��h�TUU��XsMEE./�T���b�����-�,��O�>YZY�T��8���եŢ{6�|�<[#���ttt��x�����~��4�-�<�����0���/��ug#�PO&_��_I�I.0r��r������X��veFt�ѣ�g��#���ܘ/��%��\U�xv��	��u�s��7vw^~�q��89�&�%�l���o;e�U5�97�=?D�HNLI[XyK�.�ƽ{p��zW-,�B����#V���Θn+\����ēG��ƿZ.�-7�B��}k��6u��;Yc�
����I���gE�ܠ1p9��ƙʇr�3�wA�����Lk�Fcn��Y��=��;8hu[7h��A���Ǯ�x�<�PEA[z��ֆ�^rCl̽�$��,<�jh D �N�Q�u%%��ѱCYn�	/����
dC"_\?������F�������?��^H7%+�Xp:$e���{NS�c�	����̾�+�]����^3�p�����1'� �HL���
������;,zxtFIA�Gq+~r�"�p+�;W&	&��*4;�E����ݬ-����Zj��-n'l�}|p3�n��[�z�|:�Te���iv�	���0�Ӝ0�<)m"��#���gj�IT�*���ɉ����s�sN|��h�ąh
j��D&�"�+H�F|��&_�����sDr��g<�]v���IH(�{��"}w���qN��A���"�W\N⊷�0�nj�((xq�G`��������{ˎ��d�w-��x���m+]	ߓ��́�A\�$� '"h�a��LQg7�/���%i���!���j��xe����[��}��+έ,�um4�>)�d��m`�p�le�����J��d����L?'U#�D������\�D�V�{{�o/���*�:ݹ�t�cՇ���I�!$�?r�W�T��G*#�d]�ud}&.��#��ׇUf�!;�_%J�IAD��;L�W�C$0)�@���])q��&�+�BP��aC3����]�$�?m�+OGr�V�|(��y���_X��mq�KO>��5[� 7��[
��o�zJ{�׋�������J�a�U����nC���4�Oq���*6���.��Ы�H���~��I�I��*U�3�N��2����BE%�ӑA���~a�/�h�<�y+�����!pz��ܯ�/oٴ���g��qI�)q���3o��꼹�и����V�9�̅7�D�%�I�<1W �8L���f�nD�-��Uyɩwp�͏�\H;��������O�M�����_\bk{c�*f��՞7eU�]���7y����c�Q�u��x�
�w��q��ȍ]"%��VjJ�s���v+�Z��F��A�a �(��t���B�.23O�OU4==�g*���	(� 1@�Fn�ݘ��M���t��w��Ê���C��^��K��g��k�Vxz���5]fBZ�dB����ځ��f�����;�{>X)�^s�|}���m����?q?�ī]��㨅vHk�O��K��~����z�����,��Xlf�?É�)�]g����'a����3��֬޶���3�s8����R����Bσ�*_L(�AQ_E63�6�=}��
�R�ZjB�+�MRvGøQ;��+������M���qwk����v=ͭ��C{e�/%U�Tul��7g�i{K�m��6�a�����ܾO͉�.a���6W�[V�����{#`z���&

C�T�//%��a1��	#�Ǐ�#kTwF?��ִ+o;��~�w�_Sw��G�6�*�V��)��o�MvD��M���֎�D�L��>��ʻ��s��?.���w4fRմEm��I���i��������L��M��۔ǿ_+�n9$b��,¡Ӛ�\�DB��d��H[��r}bO��Xe8��Z��kl�Y�s~���ȩp(-���o�������<״s�B�Rxi��N/pȭO�;8[~H1Ǳ��j��T�i_i����~Z1�'���CH�ś��?@!1������%���_����5LY�=Ly�ț����[ށ��Z� @��
y�{Ə���F�Y%��w�:��z\�«���l�y�?��j��sw�9D�f	�l�c�8�/�R�++8DT�.�X�\��T�\N����Dɗ/UIi74X��l�/49)��t]�*���M�z�ۓ⎗�ؒ��>t������~O*"|��e���od��u`�؆<����G�q�oN�?���#��knS���`^<km__��).iף����E��<E����3!pc62��͏�q����JG�8��X��avN�ZEv�L�|:������@�1�{��B��`��F�]��u��_�r�����و�\z�ԝP��e*~�e�f�������⤠l��>W�ۙBkS�񽐔BIH���\�)Qc9���,�w��"�[g�� }5Oi��R3.�**����H��P}�|�L#v'�쯺��8��N�r9[�X}��۷���V�I��TK���A�P�T�I��&ܭ�f\7��첩�0{T4��HBJ���}�Ӥ�����Ge��~�b��~kʭX�j��� ����x�9�m!Ŕ�J N�N�d1N8* 2R>�v�#Mw�a穂���+� ���w.,88���D���je���w�.X-i�<�e17}�;����/��pnyQ�k�ȧ���8�ږQ�M
��Pp��%w�ƆO�]%�գU��b՞@�pq(��ߣ>�Q�]�6���n�L��jG��4u �`�Q�]=�j�dd��i�K��o����\�K�W���%6���iRR��9G'd�T�xyx���wy�pb��)�Zsb8��6������Q�p|!�jRR��6o��t��k����dk H�$�ʳ�R��W�7}�?����� q�c@���l<��5���T���֢î�n<E� QY�߷:,V�r�`�\N��W��4#����"Y�>�*,Ǽ|pwG�����#���^��a���V��]3�|�N��ַ��C{�4>�%X�p
�`O�|	ʗn��c�E�4*�o�i)���Ywk]�Uƪ�N�#[��+�٩i7�޾b���������M��|	�wU�6W�-�T+l&ʲ*�~��(E�2��U��P�h�̌�l+0�����N׽a�`���QI�m;T=�NZ!-Mˋ"�#?I��_w�-�64	�|���ۿ� ����HpJO>sI���Fuff�Y�A)���K��]�'��$f� a�x|�T^��ԉK�(Y,��װ�Xk�\~�p�6jD}���]�l�R�~tm׀�ٟ3!�h����b�bN��yt�����m���ح�=$d��x�����y�'$��%YX�w�+V0лyЖ-f{$'���*��h���;�~l�Н�,�a5���'�5�Z�]L�����/"��y�L�5�g'�jK��dv%*�UWx>��?� /��#Y'@K���YV/.����а�u<8܇}��_�΋7��c�_h��F����iE
��1�ͯN2�������a���I$`��}#[�nT&y����\�����s+3�z��_`�BО�?�b7���#���Ğ�N�㕕>`]@E�WMSA@��{r��r�~rk������m�So�ć3�D���8���U�r��J.^n4�~:��,����Ao�r���2 i��P��G*�&]$V#���q��IǏ& +d�אoJ�ӯ���T�"�g��Ñ�i�@�uhܳAoZ%
�`�)��'@g�Z�D��_��	�a|�D�]Kμ*�Qԝ��6�~0c�8�fƒm-���3B.>�;���y�wl;["g�SI�ma�-�6�-O�\��v��(�\	.�(de����Qs��{�Ev2���(<��<h��M���ٓ�L �&_VA@'ƍ��!�>�?0p� �R~�5۶�1RoL�#�w*#���z��_�B�#� �Hjm ���,�Rۯ�Z���0����c��>s$����)�׈�?��@�v4�,a5�}���#N�H�G��8���WV���u�6���������ؓ�_3��<�Kj��<'7��l�5[��`�q 7���c����&և�32TTG��nx�s҆�2�nN@`@�H2|�:�<>te�R��f�y�.?,p0�S4�\A�	v �n'+ې����"�vݹ�L:��.o�H2�����T�����j������Xr��-G@�CE�p�+���&���&�sj�}��r�:��{���h�N��.H��U�������Wc����S����D�����zc�R,ù�Vc?ը�;
f���P�}mT�rK�\�a��7�=�k�ݯ��eq��̶'����=��#�0�2�3�ם~���sp�z����$��t��.u���݃'R���^��0Tq�����L���go��ƶjhb��	n{Y����Ր��M�MON�h������綐����&�P� �x��lM�O!y������5׏ ��e�o�1�ĄKUώّP�U*Q��7�]�V��q	��r#�\�`g��-=ofb�y`�`�s��;����
Vb�iK�y��`���Ԧ�J�5�-����J\a�ڍu�C;(����~p��a�t!�����e9� �u��V�P�{��p��ǝ��-�1zH�|,׺��I['[��Ĝ�ga���ϔ xGĸ�0�/��z��n��!#7s��ԁЧ8;w���Jd!�F����1���|S��%���'�*�'�����۴�Mhb��DM��h�21+� ��������n~�.7P�l��0��S?����j�l��
�'2��Z���ees%Rs��[/��>M�ɱ� �}4�p�#g�ޯ�#�
�S9FZY�?mSӇ?�O�PE� �?-Es��Q�*cb �qV��6�L��m9���6�z=����&,Lhx�ơb�aJ�	8/�v�"���g��� 9�۩��f�w�%31��E�`3�9�wTLt'hU���݈��rb���.j��4����A9"�"���c+�7�k5$�ϑK�F��D�w��4+zi���ٚ�DZA�	�^���Ø�um�y�ʌD�늤�̙�Ǎ������d}#�W[
��ν�ly���9��1f�Ij�X&�����U�C?1|-I��"_�%���wZ�6�s��*����M���5�2p�q��K�T_�c�b���6{�Q�������)e�
/aU��[:3B�a[z�����򟐓#�a�%7��t�����(�Ă\!������JP.�景��g�}��NW�앓�޳���O�Y��@����$9������v�C��ގ����*S��/蛜#9�{���JU�R�i�_�%g�w�'��8�VAy�GG/�86L_?"��V:�����,s������O��M(���WU��@�B0��g��n�Q��eJ��J�B'��r{��A�'A��i��U��:�����Cy�Mn<�-'=M���ت�NqD���m���_*��|�!HҶ�Qe���l�2��Ⱦ/I�b[5�u��T��2hi���C���*:`��yd0�����rC��e��$e�/����8fr�U�.�E[r�m$R*	�RcW#�o'��ʥQ����������ۏMݔ�h>�r+�}uk�"G���d���T�Ѓ2[^��'%���Rה�D�����e7�b��^1dN�[�8m��g��t�SCN#��-����I���2I��Ҟ�'��Θ����v������d�ݓ�]�l��5z]�zfh/^bW�YP��6����ϵ�uuu_���1oG~�P��b�Q~y�v{}�����+jC6�*��F5>��Z�az��J战43j:�S;2�h���i``���2Y���͡s�f�S�h��ȥ��b���vX�H��|��4�ZּՐ��8S���/�Y�i���4�C�I]	��$�ݱEL��}��8���jm�2��d�}���O�ʱ1t�����xu��m,�D�L�@�p�^���8?�C	ų��+"/.+F�r}V���yc�)��UB?��6��>A����+ŋ�VR/��Y�6�W2�����ݡCw7y�>|�|C}�|�O�!����	/V��}�0�O�o/�K͜�-�Q{�7�/��A���9��ٹX����:v_F�<�ǡlw��z�x��]���+��) ���\ZU�t.�|af���\쳨\�Y��y�+��Ǚ�-�n������"���q<Kd����gJV��UWe�C�E� �e]�q����1��:yO�����n���_�q{d����)#�܂fH8�Ȭ�!��6��6Y�B�]�*�q��#j=�!�F��=�ޥ������ ��`7�S�(��CQQ�dׯ�����$�$�Tm�Ú�4=3�6a��lc�}��b`:�\�^ڧQ�ֺd��2S�u�ǝ<���+�Ki����:as�����7�,�+8jq}9�O{���z���l�f�c'��XtL���b�Y3k[���+3? �4�dc7���A�F��o;\xD�v�ӼABzj�G�5RUjnk+��v��UtWަ���v�#$>/�Z�~����OB*�����HY���ڼ���\nJJ
)���G/?����y�U��!�B�a��{�Us���A]�j�vX�;���ni����j��/�C1A"�ԥ��V��U����{������D˪���Դk?v�����7��Aǉ�����3�N�ǆ�VT�B*���2b�Τ������Ǯ}�"�X����`����{����%�0�bwU������w�G;�Pd�ڋ��J����c�(ΰ~t�f���Ž���7����_v������T8�ځ�}�;����.�<�0t���m��*�s����'ϴ�� 2RGE����ia�A�TP�O�?��~�an�T�m�K߱���6��cP��޾�PN���[��]Ʋ�$R#s��[U�{��t��[��n���^;z.����N���j���C�i&%%�l��r���܅Ґ"����wE�������'"�N���-,F�MϞ=��!}ثfmӿha
�8kH�ª�л�xƋ��_g�e��cc���F]���V\Wb�zX-'��5J��ٞ��������{!�ٽ�ϊ�s�pU��^�����=%�Z���+�H�/��H��M�����/,B��s<���l�}dr����|��VwQi�v冽vխ�gF:BO��Q��g��A\�?t�U(7�>A/o#	�վ�ٗ�=8�JY�s��~{޽�q��o�L���%s�G�Z�	^��K����i��r��P�$��i��ǆ؉��W����׌^@��"��1Ӎ�-3%<ۭ쎍RR�ÚY�@�����r1�&��+�J��RE�h`��G�=���U�.�?���W���%y �T�n���O�lWW]��]�'��W7����2��PZ7��\���C	�C�$���c$c��������y�a�������j�6RYY�1騅{���J��z������a�}��/�ɏ�l�N�)�V�t���W���ś[ޛ��D�*zꫯ@���.�/�d{\!��Ϸ�`�󥥘�AUꊽv�Ŋ�M������^��&�%bK��P"�]
�D��,--����J4�����|���\*ب(!�bI��i��܎��f��CR,z8�@���� <�r�.:�����d[Ntۥ1� gd4Y��|lT��ݏ��YN��5Ca�ͳ�� .7W<�x@b�t�U͌E�D����l5�<!�2�̻�˜�h���O+Y�w �жoO��J��r\w����=,{�}>E��[TJ;�C�9ن��~���ݞ�����f&٨��B6(;2���\.��9].x�Tp󷝡V:�)���1%2/.�Rb�A�l�˺=�ȼkęېd��w�xei�(�U��I\I�^��Yv]��5��bG\e��^)7F�����02�.>ƹ�o� �k'�Ge#.,,;��+�ɽ1���%�ȅܺ�;�����ש_���
z�HN.E(��h�p��N[(�fn�xV`s������f2q�6�c�F��x`��H���+�<�I�n�������nBG���;u6e�01!���P�T�Ʌ�K��l���h��=��֍,G�v*;�@�0q����`�Ѣ��!���DtB�m�w�6B��p/�����c���� ��WfyԤ�^��e�{�8Z�T;�_&�q5���?�}��j�����aQ�]�8��� (!"�#���R�)!�4!)(�!� �9��H�(1RC� ���y�������}x73��^k���=3N7��xPMR�7W�=8) �:��Z�8� N`��`��]��w��4���s^?��th��0���{�O9��ӊ"��Ĥ㮘��_�e��q���K��Z%�og������z&L��)1ҍ��FUV��K_��a���LUP���=�ሺL$�[�����z����/�y)G�(^�A�X}��NN?���!oS����4���d����Լw4U�J�����'}�
���Z
ԷM����Z���n���S)+����[LM8i��zq�ߚ�W`�ssM���MՉ�?,��|�9��)�A�b�iŽ�I�U���ƀP�ȼ�1>��!V���H|���$q���5�z�cL�	��c[�����fa��#+c����\駄�����&�Ɍ����!#+�^�	}��8�_vdۉb����!,]5/4T[�Y��N��D�g!5k���������ϣ��̏�ZP!rb�rX�$τ�s*�ӹ7s{>��kM!���Sa�m/�J9!���;�kHaJ(5�� ��`{�{���1�+��7+0����!ꮑMeW>QHH.l9��̘[�-E9Zk/�����b�W���o�-;�T.&[ ^��)i���(�������{�O%�Pm��" �'�r��j��l�6��AOGWP�-ގ���6����n�G�X*Q���D\�]�u��Ed�'�'���;���:�^���F�n���/�M�Z3B�9+�VN�x�V�U@�4�ʹ�AV��SEo՝N�@9*�p~B���39��������n�pF�k\�OM��_rtt:��\0UY�ܽZ�(|�j�V��}����iFQŽ�z+�%h�'��tȪ�=�11.�Hx�Y�����N�4tP��d��5���b���v��w�.�K�yF�����kP��{*�*�α�n�#q�]�����!�����C��XCz�v�\���v��GH�f�4e�ͻ�0�=��r��=�B�qwp�;��d����8�~�r�r�f�?O�h���c��#<����\��no;)**9!�����{�u��Tx[���巠�ǔ�؅Ƚ����{s�V؁��p��4�*��Qjfa�$�M�����T}�`mY�)
��E|#(�������퓗ܕ }K�4���� ���ƹ�r�Y�E.)b�7�꽂�������O'��^�?�T�5��iw�`n���ɠ\]��6�+�
���:��k�V09�����VA�0	����B��=�t��={���}����z��A�A�x3�8�=�����A�ttI�ɉ�#��h�ۿr52���F�ӄ�ZH(XV,�6O4�m��R�{��]=��dUyhSܰ g���ߣ�X��[��N��S���)�{�q�ـ�`�����1[����<5<�=ߣ�����9*+* �-襻�i`��=���R���q{��KTg0)�����£&��kO�<��-K!��?d|-���.����64*����=T�-ju�����ͷgT]c2}4��,�#\l�ԩ���/Eq�+�.�T�*6&?��"B�'<�|��/�a�i�!K��n]���T�߰G�c�O�d�J���L�4��H��\���j!(����D5�"�,[�t�_�j�"3�F��O)�e�o�̯U����v����qZ�ʗ6>��,�Uru�nS�d}�H�����c2�+
5�$�im������Rs��f�9̻�ʿY�Q�Ds�(Vk������b��H��i%�OȲT��[��iB��@U��NŊt���SM�`0��Z��Y����G;�{/SN2��O֬Z�%����D���m��j�DW+y.�������KXn�>=�~��8�{�ׯb]ïBz]7�ߑ�c5�,�{��5�[m4(Mo ��9��b���[�5�>�#(�j��}D3�S���3)�OlZ��~<=dY�ͽ�I�#�.C���C_]��y�"?�O'����`AK�6z�y�|�w
��^�k	�z�PV0�7��r�p?=��5+�nEI�$�g8��=�C�18I�/�M�ס�_~LgaEѿn"���Y�5�X@#Şk���va�����1@�AJ���C�Cc���x�u5���Z�S�qz�V���r>tR�� G�;���
�`��"�N����7 K�e��L�8k���Vٗ��u�KC_X�6{�K�e���X��s���!Tĥr������r����i� 	{�Z��U����Rd�(��QZ���X.z����c'='� އ���R���/|Ò>�����Jג+�|l��ï��)'�9��Z���x�k]�1�E�:@�� �`�J�S�72���@��X����>��gl*u�hg�w��-�}��4�Vt4�'�>������
����uN#������D醾���� �b}Å�b�����2OP�.������ݕۋ�}�{�Q�4u/q�f��Io"י��0P���툝�5U�S�5\EÎn?�x�H����:�0.R&�^Z��He��GT�L���F�E.���T^xV~ڈp���)nzzz��t%eH��[�����O�ڷ��h��W�����[�K����-Yn�(p��� �CK�&%���xQI��P���t@��9:-�D4��!B5t�F�t�l�~�8�EaC=�K�����g�M7PmUz�}|���A�Ɗ���Q/���s�V��y��sQ-���TXg Ƀ�,�!��c>��S�{�ز��b~�W�{�b��>��/���� ����Ɉ�������f�y@��Qn s�����>��_�Rmҏ�j����t�Bq��ɔ@,ͺ�;m4�����x*�$����L�`�RTo���V9�>�m-����9�>��ܝ�0�4J�7�X$$��)'/���~4��ü��p$����AS�oZ���w�e���?tW�}�֯t�	D).2� ]����C����-s�ĵ]�Q��*���N��j��V�̹Oj+�k��h��`p��9���+h�Ҩ���	O.��}��j.=�W�ii�����ޚ�%Уh(&� <cp�5c:�2n�� N�A�"��0Z�G�L���*��O辩H�mlSSI�,�V�x�Z���(
���z��Yo$I��KN���c���sF�k�	���|�&���氵ӕQ��>iz��݅M�FmU����nE,��W�����H�q|�i@�h��4k�8���u�o�U2�h�XYY�	A�`��g��~T�PD���4z
�?�=L�&$bA�GI����]�ܿ��^
Ʈ�AD�Zn.�8��c(���o|B�`4y��un�S�:��t�����T0s�j9>�X��,P#��y0�-?�8H��S7��S���^䞯;p�ݢs|Ş텃n�Z����Հ邏x����LB>�zy�?����V,�%D��V�G�dc<�d�AE��P�t���ISrr��ک�օ��v�������ܣp|t�h���A+��R�/:�N
��uP>2'D�]����,H�N�y�8�������XTX��"��\���j���l�9i�i�L�᫓vMi��d���
 4V��#��3�1��W�!~ݧr��5'���޸���Cxx��ۆ@ۯG���t��t��9�0�7�Bэ��|@�q'''��i�)s񣱸/_@�?�LFb���ht?^}�V)��p�j��_��+��c�N�-�x�)��/�S���^g��P.3�y�5k���R��2��^�%��B{ �4� %Y�=�*��o8Q���r�Թ[��(SN1(>��O�6Z�XZs�`��F�Ζ^շ��X�����	�%"�ܚ�7���� N�k?�5.��~���M�ŷ��<�T�����I���^�P�I��צ��v��nBmg
n��K5��1�X��Y
7���6utZg�M�9��5u����CZ�k�Y�@m��GWO�kuCθ��Ԇm}���2��{F#	@%������l6Z��������̣2��	�a�<�GC���w��vv����Ӷ�!K��)s�9l=T�m��p��p&2����9.����]������d�u ���ʮ���@b���=��+;��B�P1�Z����;�웃r��;����M+����4b}����^��.ÓW @;h�����5<�3���o�}����Z������\�o�ۻ-�4�� �u:r�tr�9Fܖz��	To�}1�V�S�%�_���<����b���
�C�U��c]V��}ҋ� D@�'z��Ժt�sh~�A_Oٗ"x]��2+�I$�X�]�ߓ�5�%*C��-TVh����������w�d�
�{u���Q	�$&X���4Q�JF�^K~ʆr�?>�?�������jBs�]�f� F�ـ�z�(� g/vwdo=k�l�L�S��.&��ATgx �(~�4ou��)�n~�;dI!��8Ȗ�E�(v�ݵ�e_��rl�@ӏy�G���Md~u�mO�]t�wEN-(��;EޞS�Շuǭ���B��� A���H_���JՆ,(�����'����@1
����ǚ���3G�����4�Q�} ��9q�M�X*���e
gsD���3���Ϗ��{�c],�y03�j��s:V�e��6s:��#�1P��R�S��`���BR��,U���uٞ�\ّ�I薟�����*�Uh�
�}���(������S����8�fh|��Xw&�<�w�x���=�}���x:��ϭ>�"��S��y���q�jV����c�}�%s=|J�t�T�C�w%Ùގ���z���:��e����銐k������`���ʆ��fD�+9��ʶ&I���v<�y�,��m�B,�C3�`eo��s���'_���r�>E�Q*� �����?��r��i�:�̊�m:�ￓcu�����M�?��t.'�!t�s �ֻv���Rn�̃���[WM1�$��GU��n�޾ىok5����h�������0`�(�Oυ��`���k�%���!�`ܧ�j�l��F���#�z�gE��6����|��Z_��h���%R[.�	z���)!����"�[&�Д���A\��� C�`_�F�2`�����^G�����O*Myo�������^΅a�>���b�u������;����i��'d��f�}��wh
���癭N��o�Z=wQ���F�2""�f2���EY-U���s}�fs��ո��-Z�����`�����9!5��pYz(J��0��6^g��[��,)�-��d�1WE⾱��N��S�����ӿ�0
fU�j��+�� +�4���z�l{��M��y�>(�Dr��c�=�42=}G�� M��E�>}�he��Ve�JƛjI�]87v�O�������g�����Yx�����#��?W�l={��e�D�)XgT��#�d���FW#��J
)I��􂊘'$D�����H4ltTH�e��^�X�%�����n3�M��w����� 3�j���WP��Sv�_�	\����uBP��1U��U��A��D!��n}?\8 ��^�?����Zw|"I�+�֎�"J�/�i���9If��/��p��b+���(����ː�%��#{u���Y�GX��$qh=����Q'���0' �����Zo�)tܠ�	�ɖ�*�g��w&'dԣ�m��wi)}�&p���1�Uf���2��[���O���9��ͥ"���WS9b6ڻ����z:�v�g������X3�i����p�V�}[6���{�;��������z���1�U�>ch}ܠ�.8��+I��:䴑�d	���%�p↽�yI�\9��.��X�!ws��X;f�;�Y����|0�-i�w*��P|$
2FI�����lA�PH�*��� �7�r^��#U��P�NsrP�ąt9;ɂd��h�����,�Hg>���׫�m�{P��m�a߅������Y�q �xzѷ?�F�EM�>JD�~_`�Sh��c��B���;�׽Q��S��
2N��x��(�2;�.�M�K�L;�_.�#w;t�z����lڇ�1^�mc�{k��&�$�<���#G�n �l���e�|s�>��ۨt�w?=9ޜ�Tb��l{}�6�_	��U�k�h_�B�CJL���Q0�i5_�d�wH"�J�Y�k�&W7:��:��g�og��YШ�ڮ(??�nt2�����{��T�$�dP��֚������Td1�{ �L�0�GE�\f[�g��Rn,VH��:�!LΈ�D�]_ULL,nb�����j	]���Md�Dg����;4�O�q �{�)¦��;;;��]yY�B��6�qU�G�3�2)6�ç�}	�FcS)Y_^Rc��뗽�%GR��6i�մ�Pye�"�3�.�E����P+V"����^K���������ɱ�
 �ex����;�vO��.�Gzt�l-��)�����X|�"�-V�V���|V̩���������R���%�j�����)�'�񂕭��@��=a��Z��+�&����?������	H6��,[�[��d]���h�OLL�ߺu��y���9�_�#߅������*�<v-7��^��jC�3��(n�e�k�w6�N5����͒:��8�XN�φƈ~�wj_7��LȮ�Έ�]�>ݲ�v��K�w<��`�(MP������\TG�2U��5f����QTB���%��B��H�m�t$^p�������_�06���R�Y�����gf����J/<�qS��Q��rM	��/F���4�B_���+���xu��p�]@I��՗��ȯ�o@�RA7a�C?��#p�.����kc���>��>Z)�Ge+�2|ɡ������:tC�')ULg�T�@{G`����{Q�<@ ���6�T�� ��R��v{��oB�-�3>S���s$�,Um��4�:��+b�C�B�nwu�/Ե
C�% ���j��|��g�G���L�}V�
�e�l&;; �-���
ލZ�������D����zIƝ�|�d� �||�#Ŵ3��qY���������-Z�M9�� eF+-v��[��Q�G��(�Ł��z�����|���M�>��|or��W�f�،xW����զ���D��0�S�A����lS o��}�V��mٛ��b0��8Dk��C JH�<A#AQ�S��U� ����8��>u!n�ۢ���7�4����|W�i�t�\;&�w[�!���*v�wp�x��޼{��Y�/�g�:N�s
��=��$&���f���IK�������ӳFG)�Q*�c�%�ˇ. BM�?m�����*�GG$�Tw��o��q�0����M��ˢe�ư����3��������ΖTj��6+3R5�RϔfP���74ƶ���0j�W�f):���R��S���vJY��3�@��nQqޘ �ݛ��tYv�77�y�����[|�e�IZ��U� _X�e\i\���$�\gyi��I�r\��ӿk'�%vyj���S����C�W��֑��R9�a��|��K�΋�Y�RV������c\]�n�@�I1���D�e${l>+�'�d�4�_����B�-�;飤t�D��ؓA+���o"�̠��V��ר�m���nj�]�nl�k,�P �7z	��H��Ho\=B����h��Gbw��l!���V�~�s2��6���ۻ��D�Yo�p0y���+[l�T�
|N1��'ίѦЋ*;��xD�u�-�'Ľ��Yht�]U�t ��@��������o�8z�!�IF��:i<$�Sq�4�9��ʱd��a[�
�x�#<_�%�F=�zp��̭��:��@�^��%�~
�m�[�ō����N���Q�L2r�MD��yN�Vd���|@�,��?�ip�W��%�o3>��C��L�*~�D�Tc��9��!��+vd%<��O��;.b�$�D���3�<q�����Sf͍^�������W���k��"D�~��VoKO=��z���B��#�='�H`�q/
�Q��Q���Q�A�`��v3?j}���h���Y,�b�KW��������gP�$YL7�������ۣ��,
�i���w�C��\^���,��qf(�T�xP����]{F]����*��1��XQT�?i��ʭƲA B�-n
;d.O>�*�	�@�Տgp�+Y�銁\K\m6>�Q���g���ۧw�^���4̄]{3����:@+1���r��i��>Bt�����f�I@ʌt�Y��a:�Z$˳��c�]D<��g���i
�6����Z��W�F1C�R�6*ߖN�3�.�P-�?!W�z�`�Ü�ʽ�Fu^`$����&�ʃti_��6����`ؕ�Z9�7+ *3��X�����HU<����X� ZQ	U�ӳl<.�{��$-��������ob�L��S<���VΒ^�YTg�N��;�ZO�c�ם%�>�i�*aľP�)��5�4�&n�<�W'�!p��A�)8�gmm]b�8/4(��o����b:�td�W	[~�Y$��������9(�TJ~��I�iPYub�u�6Ӡ�(Í�Wt�@r3�6:�kw��.A���'0���sB���9��m	�Xn�t����R��Ԉ�(�uzsf�,o�:�u��Z\�\���Zْ����!��V�z��©�.d���S,0f}ԥ7���^����~���i��5�p�#c�Z����(#U�AF��t���K�`�h
���8�]�c�k�߄�):�4����q�F�`����i27#�����Ɋ�PضG��P.DbtHH���2>�UK1½LĎka�~�t�UV�]��3O�q�sy8E�߽=�+`9�����!��͟L�Y�ڧ������q!VrZ���M1r��oM���i`�+J�]%�5���}�� �ԃpf``�FH␄6p�]-���23���Hw�~5�������v�V��$�x��A|�L�-�l�Ь�wn:�b�w�e.(X����}b��}���X|�wW,7���w��[�}�{���5�*�g\(g�E��>!B/��o����/���Xڮ��]�DPzw_8@��>Kx�&�Ѧ"K6���/��@�K���ó��X��)��獣:�#,�1,��j����;��)(���MJ�����uP�7�[T4@��Ï���^~ڦ�S��Å�����b��(Mb���~8z��s[�ʬ�{���S�4xzt�ƫ�=թw���Q�w�����콷;a��5a]q�`�]�VlOG�2���%145���{4u���S�b�Q�Du�jar\o�H�8��C58t����"ˬH$o%�{4sB�b�J�*��cH�u|�y�F�Vc��e/� ���V+fb��ݕ aW;[Gu��h�z��G���y	��	��&i�ӊ fr ���ߌ8[x����[X�	NîsN`��W"Ia-�tQﯶ=�\�M1ٺ�[ӳ����ݬ���T�A>��*�mur"����oPL�U!�cn	�s��~ybC�����Bǎ5/�o����v-�����L=c����e�`eȇ��[�z�l��ě����u�fn�~٧a�%�f�J~c�_�q��0���>��SVt���P�2�Tq�Lq�P��?��^�#K��=ZsI*�v
R/k�~���qB�;N��������1r��.�͚��)^&@���P�x:�p9�@��R���}ԫ�D�ymIF�BL��������RǕ�d� �J�5֥��̹{����I��{�v%�\��eo�j��r���a*�`�\V�
t!_6����j���ԯ������O���l��X�Gh�R�1���R'��
6��[�n�p��<#F�N6W�xe��7����C��NĄ�I[���X�XB�몰�5ٞh4����R�=��V�����$�ɗ*�����K']�=��=���My�*���/ONV9f1I�����c�o�K�*�>}���/�|0��X�K��
6������5��#U���rs+�8�E��B,��֏��J�9���"(ب�۫֫�L/&�w~f	���|��U��kK';E
#��t����e@�skDv��'�F�}����o��/&�B>��5�A��1�oҳ��p�/��{�����?��+<�'A[5:����D�<���]b;㥽��	yV������{E���JQ�e	y��w8|}oW�2@�c
��[��x8�k�N\*���!Ʊ�7iY�����_ã/���?��qh�栩}��n�����.�{�I"t����?���ɉ����4�?�B�b:��������c�y�R%����2�M�oS����/�\�p9�p�I�b�}]�I�3�!���8�nG���Q���޻k���LU%˾��߭6*����}+4�'�zX	ò�b�[���k�QTa���8��i�#����7Eu,o��� +mP���]���,��Y�m����c��w�:�����#~r#<j,!�j�t�������*��8���Y6Ҽ��$OeP�@��<<r�M����c�AwM{�/G���#3U�ķKy��<^�p���Ehd<�3"�죴�u�E*V�������� ���}b�;���M��Q2�s�ɋrpD��h]�s�8��wb&f��_u�JM�W���3��5�P4�tQ���J��=���kϱ�٭g�nE.�-ּ�P_mʻ�I�"�M�e��Bn��(��w�	��Υ��c�����$�7*��F>�\����Ɖ	�)�x9�͌&m�R3�] �����H��,Y�r���w{8������zo��3\;�)2go���:.�j��D`��2�{a�w�r��Lets�r���rw���V@�z��y�y#�C��5�bػ\����x�����2���2M�E	���ҙ�hYݱ���eާ^c�LBJW�f��t�׷��M�m3���|4/�qg꜏���v0��n����*Z�1^�B�E��Ñ�MW��(��ʿ?�Vv����F�F�(V�V�`_U*�����;��1J��^*��+y���=��kq�-ԯ1툸L~�W¹8V���)��0$`3Y�Vl�>m��ag#r!X����~i�g�Wٽ�����/��HI��9����7��Ŷ)�~U�O�61RL�}X��u�I%��2kٴ��R���\:��b��_�Ӯ˓��T�9��O"S��'����Zy����?ڿ�˭���u�*'�9)$�%Y��J
��f�D�������K��"�H�e=@���z��×�$ױ���E�_�3]\�n�ccl[=jQr���Y�ȰM�]��R�,�.��ׄ������G
![�%+N^��/D_��A�&W`P��W�&<3/��L�<~协�F�K� s� d˾*��Lu����<�~����K�Ry=��~+������ྀ���Ƀ�k�8�W��>>R@�O��rY	[�/t�3��#�!�9=Rnyh�X�� :^��bf'Y�M`%�mkWq&�ѹ�===Ɨ�Ih�ã��G��������c��o(wAo�l���3';U�������Nʓ`�(r�i�4'��K
w�,�IA���(4h{�� �!��>*�z"j�.��.�0Y�覇[eƍ�.�ׯ_�v�E�.�m1+���p0���,�Xn�e����98Ȼ�Y�	����vHe@&��6���]|��v��y(�����DPB)�"?�a�h���,���?�:�A!�7�s��5�%�?W���K��W�O�0�V�x{�s�gϞ��A���4��}��]=����K2�nCVV�RY����H, �����h)��.�i��L�G�k�[���?@@�ܓ;l�z�R�����2r'/.Y�[O�����aQJ^��x��z>E�
y��z�">�:�q�5}Û��4[�\۫r�[�?�<ݲX��s7���H;7�gg�S��k�O���g��4y��W$�i?~�~�G�ҫ��$��u�D��[�%��<�<�<�I����Tv���!�������#@~�DE����Гp�s坹���<�V	{�:h&���:� �̜ѓy0_�s�lO���Ԯ7����	^��A�6���$��[�+�9P�!��k�5ZN�%�y�I��{Ue���2�� zE�ܕ�������	ѽ"��%���9���O{y,���k~TT��t|S���ɕ�Ҭ�����	R*8���Z�����	�3������^̉H��s;,ē-i���V�{��@�b\��Uz��وu���.�t)3�T�-@B(��\������4���M>'� F�/_���Z�@��J���-�LU���j�I�y�� 'i��0�Y!Ǚ�����v���[��!������|?e|�@U�B���7���ڂ:���VS�UY�~+��)�1�o����d1]���9ܳ窇�F?�q��2]�["~��犔x
Y�N?�� �����}B-�Ғ0�����'zc?��H?[9]br���,�"�P>�7{��_J�C �aH%�k^�}�׌��T~�۟�Id�f���)I�3�//x3��gExX9��^��s��ś�
T�U�/Ɨ ��~ދ����M�c��w�mg���5���c��x�	��l�%M�s�#��w츂��rK�{��n�H9����|�GRL50��;ܖ��Ol��]��Cڼ}�ɷ�p�������gv^dv5ΫU ������7E�r�G�������]�\���E��0-��PE�k�o3n�p>�$m���|�P�#�m_ͤ�m�< o7���O��(7��W��u;1��'G�Ie��Z��更`��)��|����%��W�e2�O6q��A^�p�.�6(�W��ܙ��|����[��Õ������Oo5Z��?�K-v�ظ�2�t�a�Bܗh�t�]���}�"�/y�vg���� �v�/*����k��3��zSh�L��*t����y��]O���Ϭ��q-��$��2�(��:�T��ɋ�`�we��"���0D��9ي�1]}	}bG�n��A*B�L��>�ΰ���,�׎��$5B�+���U均�1�>׎^�:�AO��L~P�L�C����/A_V��ƪ�W��0*���U2����fed@�~������はM�3���2`$�`�������Ŧ#t5�fc�~�W���ϧ������L��)V�<�%BS&v!�����Z�z��yf��������=%ѝ�t)��!��b��;���X9�,���z����R0R�5�U�k�'���|'�	��C���a����h����w�n^��eM��<9>���}�����M���aA ���H��|�s�3u���s.Nh���u�)x��D��yO�]&� ��

*|��	�AŮ��\<�؋>B_��ZLL�V/�,����*������|����1�5Q�#��IF���S����P=��o� Eb��+�+�|�,���n����ԍdD����c�ԁ���;�]����y*c9*S�X�]�*S�%��d(�2ce��R^NfU4QYZZb6[�Ӏ����U:n����go�.�=��6x��r@�=_��g��CO_�*�Q�g`����B�X۟H�[ڜ	kfd�@ީrǂ�w��r��8$[��K.`	c����Du���_HE�^<�i�fӉ�\Q�0��Dc[��Z�`����:L���W\���Z���Iz�CɼqϏC+��M�>ۂ����؁�Ne�j"Ǻf�#񚆞�Å���nk)ޢ���Px����hd���Y��~�'��r�^����<��l�V�5�U.EPB Mm��%�o�~C��A:#B�
�P�������0�_��ua�@� �d���
���QRd���%�3��'n�s�8]K�T�0���W�OX6�I���6ѹ=������hټh�I��KS�9|�<#�3hN�:Z嘃��|� ذ(R꼪�]���o����bF ꖗ[��.��+x�Ho��|�U-�V�+��.�d ���F��� �	�#A[SR�g����@U�!���\�H1Iv�ho-��!�i@@L�k�U�<��8�J��n/��[�c�ECx���  �����WJ��������X�cz��O8�#��-6U�@V��뫶����|P���y#��t�>�����X�3ˬ�uy\5�\��J)QH��lwo��,�P~,��χ�|���&��(qIO����uN����m�Ήr�v�r�>}Ϯ���!0D�9��DhFƛ�������0�!�V�����/�{{��.�{M`aaFc[���MVe� �4�=�V'l�]\{����w ���E��t�楿/:j�d0���*��Ց�8?]�� �c]�&��ҺB�n1L����y�[ރ�]�Lx���tжŰ�-��pee%�`�!�I0�����,��k��1@���;ڿqM�K�����C���8�4I?��L���� �� �_�w��n� ��9n*�oN:*׼���k�)�չo��>���1I���d��������ggk"@^�	̯�7S5]1��.�k�]�������gN�O���gĄ;���^���
 G�bkGE�f�
�?D�"�&@ُ:ۉ��më,t�c̀&������� q��T%����X�ݭK��n���LT�O��jyFCL:�|�]7��|UC�q���St�b ��ul��j���z������y6�:
�x����E�?��2k���
'l}� �Y�26Ӊ�|���?���Sv�t<T1�HU5h�-�ߋ�a<��[��T[������y7��S���y�H����4)׸����8��j��,�gI�%N�2��1F6����9��Kt��t�.��Ժ:�(Ŏ
� 9��[!_�7Lw!W�T�$���^|����߃���Ͷ;3��J�u�$ 5����Ą�>��ޔ����@���� =�ǭ���RU� ��QT�|���	�T<T�JO��m/C-��d���f�'���z���Y�ߢ�C-��d	�G���#��˔�hDDL[�Ug����,��~Wױ����?]�2#K���2��Ʃ]Ȫ�f�ɝ��)��&�M����,U�e�#���]5G>RH�V��P����|����*l��=��U��� )/�W�q��]�0�oh9���� R8���^���b���y�)���/h��r\Q�f�pG�'�,2ml��=*Ma���m������
A��d,,�r;���#��~6������(�˰�)��]&������d�|�G�ʽ�Y ���{3Egz3-l˯H�v��+�K-�w���b���(-�u�A!*�D���m�{`�1�u���1wP���W���r��'~V�P3�F����<7�O���,���T�H챫܏f��{&�E58������Cp�ſ�-(�D��w�G��S<�E�j�5����I	ob(B�����RV삢e�o���B`RB�`�^]%V�H	 _>�m�����͛�v�kv��u���h��j8��\�YH���Y���-�������CU�>�TVT��j����l�w��*?H��>��L=����+�"p�����>����p���Ϟb�^ �%�>{���0�۫��\���۴�%�2�#@�0��C%�j�������J�M^p�me'�����/����'��F��bzI$�6xZ��������	p�����q�M�+Z=l�ʄ�c�<X���.�$U��r��+�����@�L�����
@�F��Dr�^RwS�[])8rw�NT+{4hQ웛]<���n� ��z�}�2�ϳ!�l� ��$���K
	�9p�%���8\��(g�7b*{�e?���tL���u�*䴆�d%p9�����;���\�o{�vhӔhH�
�˴�ֳ3�(�F.9�z��M.Sf��s~O��Z��?�it��J=[�6�]�~-|�f��v�>��o��%nb:J�{{���/��\���%n�Z����w���?T��9�;#��z�9�ve>R�y@l���g�˿��<ff���t;�{RL'Q��$��E$t��?#������ȹ�rP��RƂ���SȊ�>�+��+R;5J A#4��1㔏�5w�~+�]�=Z�em�8$��z1��X4]���b�8Q��d#(B�t���3�S�����v����s��4<vì�BЏ�N�.�jҟ����6��Q��ܯ�4Ⱥtt��;�.�\�ڭЕ����J��=xHb� �����c� ��J��@����b�w�ݨ�u��7<�+��dM}Q-c�~8�	�r�aTT�z����Ԛ�����̃�)	��~��l�L	-���S��� �ާ�w�S���������M�<X ��Ja1RIE��-�k(�5XZز�|�O�K�����dR��] )� R�ja�f�)��Eqٛ�N��c]qm�n~)�P���(}�ݸ�D����÷�+�z>�P���_X�KS=�M�6�fN�A1�j�l�@+�)�4X�kkk��v̒D�L��������3��:u@���nzk��צ�B�x4 �ǘu| c�)�T< �%%tC�8󉎰#����4��5�)�G�s���9��&b$C�BF=vC� ���2�_���U#��[�Y�JG��@e�������yOpƣ{o}a��a�u��"�:��L@ ����U�ޑS9��Gυ$���4�����3�,��X��1����~�Zu:@�6��#�

z6v����a�$;V����AL�ݲ��-{���B�˿9���)�u�K��A%`�eBi�p�H��� 곲�z�c��
"1ו M\�����<*J�\i���$��AǨ�x������dПw���V@�͡��!`:8>Ξ�Q𛮙v�¢�񵍍F��'�:�?�#@�蝴���đĉΑϹ��Rl�=ޫ�)�${�<��<�����b��? ��If|V5��?V54,b���
�����l��e�ʌ[u�K���I7y�s�Z�b����i��7-��PB���C|�lD^���|̍����OFhD�h1�@�H*�%U��/.�Ł�4b
���������V�@ʬz|�	���N��{C�@��Z��'4P�7��pH�
R�� �>=�-�d�n�Z}?v�/��,dYo�f�2��&�)�y)/2���0:�2�ӿ~�2���}C_V/��?�.��R��K�����Y�3��{aw���9�j,_ߣ��Bw<��\>��W��E �`�,Xﻓ�v���.�N�[�1�����������X���)t�sX�0h=�#�L���������OD?�hFn) �Zʭ���&5u?/{3/�p�	083�aT�#&vqPR� )q_?��m�`�iH�<����*ya�jߺ��8`)���H�=ʀ�7��� ���&A;��,4[? q�R�;�7���o~S�.U��`��Q������o��
�K��t
�
�\i�ːJ �qe)a=���5�����&�K��j g�2S���/~(wk�p��@�v��
��%�!����a�n^ �T@�%Sd�^�f���s^	C%�?Wa<�|�j�ov�Aӑ��8c\�Z�9v�-�X�̺�PƆ�R�0%��8U��{w��П�F�b����0�����p#IhE����/JHI��b�+l��� ��
�t��T����8��[P��LU/b�KR�C1i�X�&��}Ƌ��)��w�a�a돤6�F��Ԥ#���xu�x�v�k�r3y�{������$+�X�1�c�jڇ5=�6�r��t}	4�mԶ���@B�B�P�y.S"�p����<dh"N$3!�1T8f*���9�c���?�8�����[�]�w����}�{_�������K�2CU�����b�d���-L�0�^]��Ax��庩S�'�!J ��J	$�Z'��'b�5p��k:@�ɣ��B�+~]�Y�4�J�x��c �!�u�T/���c�������A������C&3�n0������rO���x�t~��G�%[�.,�#j�]8�t|��٤r�?��ʉc�>��:ـ��w,��<A@X#���>��_�r`���w�	���Ue�F�څP�i��W�U��?��'��N%�D\!A���|��5)2���`���*wSA>���~�4�	bS��N���C�A����T�+_N,mSgh'��q��FM䩼���a\~W�a�_��ۉ�������J����"��;�9g�vaq<O�4uͩl��bl�mhb"tCF��{�Lj�c-,,h��3XsTw���"C���_��r�Rg�����Գ��?��V�Fi@z{��}y��,��f��ͩ�r5ޘ'ŦXRA���%�sl۵K u�vV���I�"�¥q���O��V�噀d��:ϔ�/C8U�f�ѧܪ7�Sf=�11������j3�N���k��8��C�6
i�R��BA�r�^�:O��RQ�!���q�i ���B�k��!��@8x�a?m@ �	���K*@AH%�U͖"\�FV�ѨI�̄��B�`��w���D����W�	�=g|J��U�;����{�_C)���W�`7D�|��Kp��{tQ�!�9$34�5{�mG���5�os�RO��.�#��Z�3��D������	t�aӧyy$ʄ
p/����b^l��L
{�/t�P���S�}4�����מ8�ckX���)�Z�Br~>�S�K�kC��4ueF��j��+-�8�O��;ߺ��@:�z���ݻ����V[N�i�I��#]����LϨ�CsQ���f�*��;���f~��N逺&�V^H��D�Kp`�>d_���_�7�Ib�b���-x
� �h+�E�9H�.�iE݁@ɻ��Gǻ	q�E���(Βêt�/,��O��G��Mg\�>��}'O=��UR���3f�S|322���Z�S+^0��(��ڴ�oP��$:�M�ģ�	V*e �)�@��,��`��|djsF&~�#��\b)6z�ށ����꾩�v�A�4�<mp@�o��(5�vAE=� ���r��Ⱦ��3㝂(;����w��hI ��u�C��rL��,v��� o�
�=A8�>�j����M���	R��ڬ�f�*^�+V)C���)X�rH�q�	�����| J5�Ρ�W�*fg��P��R����Q^����Ry��qq���r�!��lV���O+;�d�$�"��5�Z�o��~$�hTѓ�Mf.\dW}�@p$f��Zd�W�g3߸޺pjh��b2tZ���;d��+���� GpvnAv�'�iC:�z�<vL�Y���;��iL�3����wA�ֺ�/Vw��2�W-�Jҹ.I�����`n�}�Էu<�	��2�S��3�/��S�jQ�����ʭ���_�(�50�27#H���4�ԉCj]*xd��=�N�qZ^S�(� �6�� ���%#i�q�JS\A#�Nr�BpW)�4�K�֥W�/4����4Vݤ�޶��?�Cc�W�;�\b���ٯ9��ߡ�ڋ�%-�����/�P@�3��6���™ѵ�i7v�IާCv1|se��r��x�q�ImE[������;�1Aq��I"j�u,Q���U�@�T��3?qi�5��Zj���y��ẓ�-���٨ �U������v�������ƥ7k�2f�ب��MG�S�~�E��'�}O�Hu��pJ��%g� } 2��w�1`�X���������¯yrW�+#%^䨦p![��CۈWc:c�빶�ըٴ�	t~_�шw��A���u*Rh����>�)�Z��[���E9)Γ�>={�������G�O�n/\_1�^�Y�!��KA���������N��gk����iyb��o�(�?@m"���O1ہ������Z�lǆ�7�}X�GCL��<��Ŝ*�*�DKvp�m���zy�X�xj���z�"��z��66619iF8zK{�a���V���G�P��=�2�ۻ3D�	t�`�A�;��S:k���~<�6+��sD Q�WB!���])ר�J�$�ɒ8n�zh���a(2���P�:�����;���(�Ly������R��G�5�G˖U���)[(k�`�c�.���?���ϯ��퇲/�\�hK��/���6�?��2Z�U ��������g���O�5)�����C�^u�V�x5���I91t�>y�$G�g�M�o�}# ��P��n�!�S���as�O-i���l��S�C
4#����J-��o���!���>�s�[	���"�s�o4��K=sV��6v�?{z|���]��w�;'����xļƬ���[��83	��)�s�����N'XS��*ʊi����n=�cO�d��-{�#3��6R�6��.}�YB�^�w��&b���0�Y�B��Zf��<���:7$G�|��+�k���Q�eYԭ]���t��?ud<
˒��XM�	W�{�8�����讆ٿg�0n��5�q0�N��z��X�w�=�r5�7I?�+�������G�6�1f�;(��A	���AY�@"���_�7iJ�|PypY�Ro_���G��2�8}Ӯ����`��8����H�vܔ�
��k+M3����� �m��L�E`L��A����7��P��9����/u���-��]���{)���p�SF~ڬ�aR�Aμ"�^�T/�^��q�qt?��ha�9Gݣya�v���q�р�C���鳡꛳��,g:%�^�Rלh�����1�4	����|�(e�p��7v���i!��S�y����5�}��;�l��[����>Fh�Yխ���u���fN�	�U0'����>{+-&-���T޼X�n�蔴��I��<
�����8�O��/�HD8��Q�Zk��2c��/��������0?��%� ��wM�fB|��*մK�g@���{�	�:�RJ;1��?)	��u����<Y��#k���s��;�@��!Gai������9`�V�������L��ʣ�#`����[P��O֙9-�Ͽګ\"��T�����N u����U��֝W�.���N�L�J��1R��y"\ �9���*�W���9���cf߮*�Z����,pڞjF��������τ���2��k�!��i�����߸ ��W&��c|�@�U͟RQ~��T��1��l�Yq�+Ρ����҅�Ҟ{6}���x�������t���|E؄�+w�L��DQ^�?Z?F�)zX��m�5揰hp�6��:��|e�*�b�j��[cmQ��R�I)����y���Bâ���~�"#no�=^�
4c?"���;���3��C����7��0u
v�}�Dg���@�r��p��vw̤%��6c|t�Y�R��2J�Ϗ���S=99�ő9�"���}��吹˥?�\� �9/V���KH@h����\��5j�܏М@Z�@?G�R��+���Ԣ?o4�ff)e`�Cv o�F.�h�*�T�����J��t|���@BL�~�/P�f�����hVZ��ly�V�_�;O(��̋j7�dk��`���N0J���;~'n��ḨG���3����)��O+���=ڪ��ѧ��G��Xo+/b�	�.�m�OD��Rr�;E��؆O`o>q�Έ`�Nr����%�����qo�E���j��Ɛ>m�B���C��3.,J\ s�7���x�N���E��w�V���T$Jt�p�ڀ/��{*�������^F��<�+hx�$�9��E3���a�d<�ʆ����e�B[o��D�Ѯ�����ֲ���ן6/jTF���2��Og��~xU�_58��e݂�ލ����F��ٖ��y�7,^#�����Nk��(֞"����026���[]���D0~�(�<�S���A�z���@�{(�uP]���@)���JN}�L[�!̚

O�.?�S2p2�$KǄ7*	���K��$��,)�Y�W�;R
@f>5�n{��}��+מ�
�#��T�椸lǉ�����1w^{ 3;4�
t�9����$z��?��Uԭ��՚�����L[�v�_�VV|6T�G�&�8�K���{�CԓE���c+ ���\}�������Q�8���*z���T�W���:_]����~&$C�o�v�Ģ��d�4fd�T���o�dpl�3�K�Ɉ�~����N�_  o)�������K�	�g��KJEQ���<˫ �����M�=�+���hk)<�'���g�׶�$�gk��,S�s[��!������w3[�&TI�h�*��&�y<=#$eY�F?�L]�/�':q
��b���ۿ�!ǊXo�s��k7]�0(�?�q;3�Ϊ9��.��=f\Ą���V��,d�jm
 ���1f�I�����;52=Fwg� C�/�Cc3���C�H�UB�#@л�ol����֌k�\�9�Ty/����ܭ�,��B
͑�z(|Y�R��\uBc��GE
�<F�(�&��*�eۯф�j9e$��$�sGz�K�/����	Ks����՚_�Nb��	bN��%'���Ӣ.O�߹��!��kʖ�=��I������~	6Z1���ABq�Y7��������5"DBO�ӳ"�����S�ІOKa�31c�c��$ �Hٗ>BX�?�v��+�?��Z��EF5�"E �z�m3>��Ψo1�?�u!��m�[�lqv�l�]�ym��"�4�`�E&���X=�0w��� �X1����
YGaS7������?[�r@N��Tf��(�oI�ǫ̫�o�f32�2�_�xj�����6ѓ#����⫴0+
>!���"D�T������f:A�G��ޖX����ݧG���\�����S�)�b��9̙���o[�E���Ƙ%3 7��1d�)))1L�66��Pby���h�Q�ؘ���c�tAT����C��&�:>WT+[t�˫�G�^�@����.?��0;��������?ߚ����P� �1K�9@�Ҝ���o-�&�p&H;R�&N���UuҨ��1�]�� &UrPt���Y[ �w��4�����2���2�/(�������+���c�������F���^��a�r�C,��
����13s�T��TZ[�����#��M�D���Q�����vv������g�^��?K���du3�����#�[4Dr���%w��,bG�����I�~�=�ؗ�G
H�9��C��|���r+4J-{y��.�B7L�����6u�Zz�ˈk���l|o~<~-��t�����?�3L�5���D�n�uZ������N��k��u;�z��V`߳��R:g��4 ��1!��j����{�N��6�$U�����Cv�m �������� ]�/�Bad)��V���d�w���*r��*�M���1�v�m���% ���Uk����`��&T�%z��M��G�I�fF��&�x^X8�y���Zr��x\>hr�*�$�{TW�R5��3�f��f!"E��$�Ǳ�#c��(�2�SBC�$<�������`�%�L~yjw�$:7J���5Vi4a������m�uVG�O�z�̨�'�Rs@̂D�.<�H�XSzy�����f���2o�a�Σ�+���J�6ݖY*�%_�D�D�4�2���O��%�e�lq/����r�����S�k�M7{?�`+��.���n�3�w��oaDX��Ǵr�V���ܦH%y�x5x�P;���`��766Z-��Wl��s�?�Mϸ ��D��q����C�>j���/60���in,z�߽��3U�d�2�<}�f&C�)�����5=VBfH��k>F> 80�j��	}���@T�#�u��J�Y�3!�@�!,�Յ��c�>'�{�Mh|eQUzW�$o�5)QM0A��O����� �=�m�_��v����u��p� Z0�����h�~���6:��_�(Q8��n�Ɔ ��)��Dɺ�]9��ok���FS��mӓ~�Wrd�c�Z�0�g��s���g�v�e#r�Y�a�v�ٍ��L$ҐE)���}H2�];����\���޿d��hn�E�Ѩ�UW���Fj`��c��$Lz��ww�*b����2�Wͱ3$9�.���+���Ϯ�[�QK�iyzbZ�/�:.
_S�^��h9��P>��X�3�}r�<��8}��G\	&��1K$K���s�y�?���'�l���9gAV�:)�-m���کKScR>g��#��)�,�<߭O���pJwB~Iq�rAQy�t{���;
=���<�㼯Z₸��D�ZFUzdǭ˃�Y�<����j�w�WȲγd!\�g%��v��SMd|��Γ׬G���x���,�%������Qg��IO��N!:��H�-�peͰ��	#$�R�K����b����[A���j
��_.���Į��+Czb�R1`|^ '��,yh�h]((,{A!��49X@��C|������y|�;u�oE�~-��8fǱ�OT���^���������"�q\^��x/����{�lc�Vg&���5�p����5b��y��Z�W��Jg[���3kUSo�L�pHK�'{���O��T5�G����!��N�E�9^�q�R��TM��kB����C�W�	cX���g����r�Z���
�p�۳�s�y��(������$n��gJ��>]�G�B&|�QVNY�P�,��R�ڛiF·�痆��s:��]Nvx�T�ѫ6Ad���ס}����ף�s���}�fr>w�/��u��� �5R�l�3�-D�L����'WkiT�+;bBG�=�3����p��=/�#��D(4�9�5�_�;sV��o�����O�a!wO9���޽��[+�f���M�`���[p�X=�Te����Gll�afdD��"�ѱ�7N��E_S�q"�������v@r�oU�V��Y�o˧C���B$^?W�"��^��.�m�=9���j�.�W5őJ$���:΍�no�]������lF�OFi?���a-�-3�$ ��Gaj2��CB|mI3TH���_ɇ�^"��H��{�n���G�����O��A���m�Q�����P��M�odYHp��g�\�Z��D!��,�2�I����H!���?Q�Q�*-�m�w`�1��5�Ͽ{�տ����E�x�v��I���H�(4�NfS��9+d�nIi<K�.���f>�ʏ��G�1�#��A��Q���O�����8j�y诵}!'}��)�g���X#D��H$wN�����T�!�kܤ��&G5�er��&+�� ��>Z#� `r8�S;�.W���o���Ӝ)&k2� ���z�&XCT�_�B�J�H]�m7k���Exݼ�"�������\3�V�Q.��Xٲ}���I:w��Ї.3_U����$�|�w!���
pʿ���O�[}5ꅢ27k|�z�ȗA�ƪ��q��b�|�L9Iq.碆�}rr��4����}��$l���Qy�(*K,%к*�a�ڨv� �E�s��H��PW�SP4%k�5�Du�<��Yw�xqRcc/H냙��F�7]�񪫫�Ix:/���kh�S���8>Q|���>�z���+�d⽾�V�ȟFvy+Yon��@���g2_�j��M��g9��[�[.}�u���'"&�O�V����n2x��1r��e����u7!r<��3�����d��~/7���hV}�`�$�����!�Nr��*��#�����iU'
|X�M".�B%���ǆ?�29�+;J�[�aN� �G����dY�D<S����{�yr�L��'� �ld�T�Ϙ�o���T|�ݣ*þ����9K���@GI���3*H�5�Xf1�F�x�mb�v|�B�@@5�>�Z�D]�����r�3���q24�&��\{$p���[�$��IU�#��̷��m��(q�A�r�L��ީ��Nb0e�R���Jm�RH	+98a#{Vj��v s �ǈ��\lHTNn�|]=�2y{��0��쒁�E{5|щG��������*8��b�bڞ"W|f?�P�/"E�mX�Y�S�L���T��J�J�$�-���6�l�;��q�� h*�B���9C����z�U�fԸ2s
/�[
�C��Z�'ʤ9�{�u�s|��f\�ڴ�µ��	5U����V*�	���]c2 ��EB�Y��@{����X/�Y}�9�.؃��1|�8Y��f�f���h��ѷ:�4R�����9զ�h��B�؈0��K��L�s]Fو<���$��v���S,����X���uaa��Ԓ�v��1�F�[A
�L��N��2[�a���͗f:_n�([�1��p 9K|���܊
�p��<����:���݃D#�dL��#.�@�w�������4�zY'�@Q3��- !��\|�A��Y��_����Q�4᫷�	c~3gǍ��M���h��@�ن�� ?����fF�c?����邡k|
�ʄ���S�y�ACuu��K��3�E��P����e���������$�2I�\T�_9φ7���I�2u�TV0��V&�rLi��&��Bz)L�b?l���'k��'dyܱ��)�9hیJN�&�>o��
|��m�a����B�\k���i��j:�>�ʀ(���^�R�bS���,���a�|hh"p@����?����sO�e(�A:E��:?�V�\�!)�-�pE�l�!����r��h�
�4s��m<􌿖k�5������,�<�9XT�X#0�b�����f�&����rvalk��
:�O�:�q�4�3�! ߌc�믵����|Gǿ W5��!�%���S��XJB����q
JA��q���j���B Jo�O���V�5��a���1����K�Pb������Fµm�&����\N>_PoU�������G��C|{��"�^�D��۳����P��P�xU.��F_�#O>�.���q����"cO�������� �u����}�RŜ,Bʖ׷_�D��O�y~!��S{��T'�w�mŶ���LT=Q���Z�z�:�sts����4��5 F�W��aj|�Ȟ��'�O��F$��E�sf8Y:��`n妷,��nL!8����g�?'��¹�z��,u�u���g�n�n����7T��Ӆ��x���<�xU~6t��^��g�^)���Mr�CIpb�k�Q)+n��|�ʳ8�Y���H3m'�"�,��~��D���/�s*�S}d���A�����Z��|�����s��������3�B_@��5+wl�F�����Z9[K���q�� )��M�!����l!z�|BB�m�(w|q����n�#	5:4p\=C+jp���w�ښ�7�_�sx���w�#ђN���]Y?%�4������Lsiz�m���W������u#\��A:)|� %m��7�|��ZEq���뤷>�#�5���pB\69J��KHDD������\��5n�V�~�7��lUq�c���S};D��{�&�����������WAb��gT^ńz6��N�T���F���d;���k�#�ZBH��{��H�X-}�$��;�"��"���g��I�|/MG�k�N��u��߄<i��T_e��s�n�(`
�VA���R���v��p'������~.#�1_pydn.��Q{Y��D5�ZR�#�.Wt�+�*����I��SJ�'�E�f#���� ������t���Ia��W��Ӻe��|��dl;�=�Ѣ�����	tZ��?J����:��18������30d��;;�\�ݶG@�8�	e_4���QS;>
���諗�/B�BM������'��v�Hm(; ����j*]�׎؈*^GhN��!*���S9���n�ﰪ����B�_�f�f�`�;E�  ))��8+�;P����K��l�"�.�c곖vXHc��L{��St�Jxom���Esa#d�%Nf�_%�_�O�ȶV����뇒���'���׿�}L��@���e�+��+G�~��7����/�h\Bτ3o���dY�0�:�%����, ��{Y�n�v��S�d�FR9�ǫ�m��+v|�2=w���E�R����1��9�DAx�d����	�1�R�x�I���z���Ud ��N�.(���Ӑ6Lp�fs�[��9N(y�i^p��/l/���?���UꀒvI�MiN�{%� �DL;�{hHW�/�g�G�	��W~ϼ��u�N�q����1A�|�+��.�ײb
��a��B|Iy+wG�����mkS]<��W��(%��^�z�&o�������n3)�F���9Фx��W4�Y��J�^
�|B���-�rښ��0�����-���"D��3}1�O��� �:��1!���R����Q���vC�$�z�]_O���!���7<�AX��=#�:զ��j�B«�wK/~/�ܙ=��D���80m�S�9�0_�:��X+ .M���~�������he�?�%�ly��t8*�����U�����I�I��_���!��J�m���9�e�w��ش�E5af��W���!]5,�i��zbF<���ـ�	�s�7P�b��{��̑���>W��ȯ�1}|�[Uk9Å�s�
�ƃX#�{�"�����}�#��JTĊOo3'��	_����Y�u��һ���'�:����Û(�'�:��y-)���C��Ϧ:��LW�"XT9b��;�cϰ��F5�O�y���]c�yǛ����Г�o����ב�s�_d��f�s�U�P0������ci�8�-Y��$D�C`����1����ZsXQ�1������\1��'-���(`�A��E���X��7l'`N��l��r������^'e�Y�i���tx@?�R��E(����]�֌4��)���5v,��~J��k�]Nԑ��m7D�������b����)���h*˽W-'6��m�jk ��ex��5�j�tW����!���7��J�z�Ooo	��=B�\�֞���/���H~�G�o��v=��+����4�b\��O��iW���q�����It�l� �V����M�����q�l �~���y�&
��#1��|�p�?�0�d���*� 9��*���#���F�fB96�C4V��y���m��=�_��~��kկ?<��m�.[|��ʪ�$�F�-�?\_�=x�=Ц��'�l�xp:@&�qq��X����||�T�hF�!�w�=��g1���1|�;�I�����^2B�S#����[�T�ۤ'���	����|�;�є��Y�9<�:gE3��;�]8N~*�f�~�_�䫜Bc��$��.�5q�Q��9Gp��ə4��~6��)�S9qz6B!�{��[�	؄~u���Щ���GD�2%3z�{R��<��w���|�F�[(��S.�[����K��������?�?ޕ8K"?݌~T�m�x�oZ7#�];��굄�'��2�˚#5<����I��y��n����νY�M��'8�D���=fU��$�<��RLd������F���75&�l�J�1�1w
��M�b8�"'G��	�Ċ]���#k"�,������;*6�/��1,׮4���(���"������.�?j���Eq�����@��i?j�!ƒ2#~��i�0�����{�N�r�s��:�E����TGJH�x3�k
c��箔r_�s�ò�H���0Y�����$�:��V+����..F��_���SSO��&t|��!�׍��G�=�2�{��ưk'@�vv���Cpl�K3�	��_��O�6'a_n�pT�RB�e�j��Y��Um�9iT@�K_l�Ö6��� 렾)H�|�ú�&V@���P���-X����g�2f�Z �Z�s7�u�{s��،����Z־ID�����rK�ʊ�r#U�eҦ�~u㈛�g�I �#�M�l�Y������v*6v�G��q�|*<Z(�븋bu��r����sc�Qɍ1�4gފ��օ:���+ߕ�%��`3�+�7\���݀"L�,�X8@� CD��@0w+���K�6������	B7o�RP��3�/=�P��V?������6��o�k�LJ��T-o�v͊[v��%I"]���yg�՜uJy`K�;H��3Yc6¯���(m��w�����՞n��a���T�YS8�:��9hF+��u�]X{?F�H���O��4���F@�[}�
�@��s���7�f�~0��S�-���/�g��(���@i3����pv�iJ��ޗ_�H՞��"����ѭ����$��?u�ES�N�a&��~N��B#TH�٥�{Q^w(q���o^G�Tf-ҚF��B,�/��G�nc�@������g?���n%�\�/�-eO�j=����JY2��!���`�ej��� �+c{ <J�#"h��蠧�oͩ�'�YaTą�{�T�=q4��0!�d:V]���X�n�M���?�&Ng�qD�&$��H�G� zu5�'N��5y+��֍KC��v�O�[�;��
��z	��N�σ��h�w��`�%���[��v�]������ /+5O;�U�"3�C�G���I���n��
6b�kˡ��K2���v�Ip��b*��xB��=M[���%�CR�.���q�T)�,+�4�Yɍ����D��볯��C��&��B`ր���13wOz��KŔ���f��Zk>�x*���v���S��kmy�wӶ�}��8	v���=]ћ礨N��5��㤖��G�1�����7�&��%ٛ��V���(U�Hx�����Yq������R݀� ��F�>�وR�w���E�Sx��ŕ�U_^�;�7�tu�X����|�����F-��[	7U�����(�|�)P�zw�b�R1jB�1�J�7�OH��a�(����1�2�H�,o��Yﳢ�x֑q����0j*��)���
 �&F�)aA�l aO���ņ��)�1�����0�$����򓧁�ͯ��a�4bk+-LsK�b��(��w�U���^u�~��i�U%���93��2z����(5�hz�T����ٽ��&č��Є�ـ���e��)(3���J=�8�MH��	/z�l$�7HT5����,dp��v����}�G�Ay�X^��XX�_�Y�W���*?L����n�cm�+h�u���g��*�ډ0�k����$@Z��:�k�Wv��36�[��X�P�r��	E�v�	�O�^�|�#������ڤ�M���{R}�̻'m��ل�]�9D��MJ�D5��9���aY�#?E8�(d��}�ʖ�>����`ǈ�L�Q�[�:�Cs���\$��HZ΍��:�vJ�yM��Z�����4L�#LK���<��m_��7ω�		مJ���V�}�O�#��e�}�*��Z��ov-O|a����n3{���G�á�cn�l� �M�R���{(]�\:���R���c_ �7B����:���.�$_���%S�P�Ž�~�"�*@���i�Z�����ayts����h�s�,W|v����a�����+W�������;evVw@%x������FS�q��f�iqEX�X��Hx���M����ut�#�븦zHYC٧����AWN����cU�^/��pF��^΀�f��(�ss.���? �>3�{JF8< *�C�qj�G���,;<3�����-��֔��;�E��uyM�Qt3e,wr'~)�`	w�3�b{S�P��|�������ث��xL"������9؂-sB㇅H��C)�Y�j��Z��������m��[�f䇏G�/;Y=&��� ��"p���I�/D�W �j:y�#�i���3 ��ԓ?f��'B8������Es�M~��c� �6R���n��JI��[M�g��@��6/Oh2�=�8�6��K�w�{�>I���ҽACQ���{��]퍐�!��)��p��#���d�A�alU��3׌l^�SJx�[iH�G� \{�u̜��|�P�P�II��]A6��A3�{���,Z����*\����qk� Ĳ�_dhx��2Xeq�ւ�=�����L�c2Y���=�呿_����'��4��g(�������Z}6�C���|1ٜ��0`I]��V��c�;���/L����Ya�e|��"ɓ����uz�YL��+F��R�_r�?p�?�(�/�QC~���50��1�Wz��u����,Ï����=u�ox�b�	u�`u�8�0"��\�W�Ҋ�V��A�=rI��q�����o7���|9x�Ro�Û{�?Dז�P�E��*K��:�A_ţ^�����bT%�G/Q���s�&�-�.{���8�a�eL/�x�P��Bq����ͷ��l�����r��n�7#�=9 ���hS��ľ^�ޒ��S��*З�Z=�v��r�� 8���T
Y�xI��>�F)����luc�a��S��"=��J�s˩?Tw��A�w��Fc�;�t��*���"�/f5��&(P~� �V��r5���i�s�3_�C]��*M�v�(*n��j�S�4��9���g�����u��-B���,q�J!�g�F�S��噀�93��@�Y|`>�+	�CK	4��>4#դ��Wc������_�^-Y�6���"�e�m(7geŖɹ�YB���l?�8���B��m5����U�ُ@�����������6��&"��m�V�����c���M�фP��ó CS����z��nj�������
ꘕT�;�y�m�NT�=׊��� 6��C�9(ľ�zn���nn��t}���w�<�m�ǰ^j��m?f_�'�
�z� -�-�����|ˑ�r���D�IC�#R8~����tȵ]�/�&��z*�'{.���;��(���������a)i�<zVs'	R��}E!��9:�J�����T_v	T��I��x�*9���Ai�ʐr��	�oT���H?�wOOh�����D�#�[�'wvل�ߎ�Fg�Er�ᴈn�ZH��oy)���/�È/�g�?,�(bNAC�P��f�pS�&G����|<K���]a靿wKz?�L�8c��ݎ�������Q;Y`G��x��}��B��\�4�vs��V��u�qERhX �wz9C���9��@n�8��AН������fh���M�&�AF����v�4���{x�x�{F���J��l���X��̬����+@:�Ӣ�� ��j
)au�Sm����ETQh��L�T��������2֥����HF)#셍E�Q��䫱������d��w�TAA�M��zn����᧡��lw��RA[[���n���Д�yC���':�d5�C|�\���4"q��g��o�G@�0�#���@p���T�z�26Q�_�I���� |��:icl�:W��W�K)�b�1G���r����>�k�Z4��a��+b��&��ꋀ�#t��o�!56�y�V%�(w���N�{�E
�)-���;At��,σ�����w5�U2f�<x+��Zfv���ŷ���<��ؚ|џ�Y��=e��&͘{h-Gd����kiL,���z�r^:	h{�{ �T�L�	S���ŶM��V9E4ARG3��O�'�;^hV�=
��|�7"|�
}��u�����R�:|F�o��Xf�ҫ�@ x@�����d��(]��v�%-��k�\HI�8�JQ@|(փ�S��W��SZK�5\��F����2S�^�bݮPjUMx����hp�v{eM���i{�G�]���߽F�m]�0��{�hԯb���̌���Ӕ�g�C|���~���I66]�~�J:T��L��C�ױ�~��^�f�-�(%����?&~�a��Q1��tA�y{R+e�\���I�Q��Fz��/�8�3�_Lp8���b�W�Y���כ�;=��'���ے�`>��g/z{�3�Nz��IZf���vTlsuǄĈ`N���P�%cf� [ʀ�������op��qThȱބ)`+I�h�c�$��lh7���֭��EM����y=㼃�/���H�n����w�(@ؓ�!�>���&w!2���/�"��9_"�:B��
<8c��σ�i��[�Tg�����qW:�v�7$��;u%#۴j؝䵻��;Um=�Mق_98-�G�H�	��� `u����j���rU�X���Ng�P���3ٚ�~�梔*��n��G�֫W�o��vcY������+wމ͊��}q�Q�t̕���_�OEL4�:,�cyN��{%��s�	YO)�1#�r�uw��{M�[GdlV���T�]�˖���m��`*"�$�F>�xܕX�~�E+�0Dsۓ���E�W�|��ÍW'����j���B�>Hf?��)��c&���_���|��D��N���D-��_GE���YU�|EA���,~�ԓ<U�wx�����\B$y��_�\�f���-h��:F�C�R����mb�>�H�s�7EJ}��`������+���!�>�/̠�ѷ�7˲B�	y����oQ��'�->�\�g���2�Uχ[��2�8H��x�)��C�$�X�����x��\���75k���K��5Pt�/Z��	B�m~��\��*ɗ�+�Ryۈ��<E�������+G�(2e�NX��T:���Y��f�
�r]�Kb̨�k��p���V87�����X����q6���(�U�w�'�
�]���yqk���<v[>�a�ʂ�k�W��z��ğ��%y�נ�y-�HN�O��%�^�"���K|�����W�H}{�x*[]� f�r�x�
C�G��� B
��"r�_XXO��M�	I*��8�6]Lp+��'d"��b(�3.�j�冡*0�뵛��A�EP��E?��R�������ͭI��ҳ��X��^������:�����N�}�qӢ���ٳg�~�����$� �.�p���;3�~B�}¥wW��#�	��^\�/���`�_T����
��E������e�ǋ��R�S)���Ԁ�f���[K	��]��/R��߁Q�����0T�{ ������nJ}�k��4<\0��0>��F�xM����|^�>2�g�Ikrs<u3�5i��ҘߓW~^^n?O7�˺�'4�i!zR��y��g�x��F7=�yd��0{/��g\�;�u����2���z�e��ޙ��IU'�b��Xdq>n��I�Y2#KÉx5d��9]®������T��8+N$.`��>��ߚBo9���m�86��S� �L	#&�G����`������ ��bn���^,9�_��U��_�w���!�'�ԭ 	"�E�?�"�]�gv�E�V��*�;�x)�{3Y�����7	�0;Y��:�<� lM��WZ��=�j^mUb�t�x����w��dN�����֚7�|M���[<A�g�&���,qj��i��VS��lw*VTRƞg�$ދ�w&$�g�x�ܺU�����L29j�(8�>~�E��9K��ظ�>����t���כ��v�MG�?�֋c���=���I��'C��T��'���A�W��q�Ԭ4;�Y�n2����~��ht����v+�ݸ�Q��������~p�9��یv�^Yx�^�����L�p!��Oݾ�k�e7��ڟRJ���g�v����?�~�Ƶ9���ʛڙ�K�L|���I��H1���3�Ƨ��E)�v����K,\}@������ɉ�鹴86�AP�2Y�ՠ�\n���K�>U�v��><q�.a��+�g_)y~2���
竫t2Yj3m�sp��r�ٿ�S�R��?�v���h˫����-�\�ok���ߘ�O�i�k��*6_�坸�l�]?¤�*�DO�>����c;;Ox�~}�&iӈ���m6���q��P����l�
Y7�%k��U�P��d��#�X�6e�hQFc�[���R1��̈́���������{~�<8<�罿^��sfLY��������m�Rg�!Fn�"	׸�U��|�z1gda~�o��#��PQ�T`P�������r۟b$��ߒ�=��x\/J�� �� ���A;�6�bw+��zfJ�*�DE7�9�����:D��dޭ����_^��4����\��t���>j��� |u [׽oS">;��s��Ω饕[�h�4-�D����I ���6�n|�N�+n^�\����,���z��C��|���I�̍��{���f8�o�����Ȑ��!��Պ����9�Q�䄹��Yy	 Y%Y�"���7�<�|m:�<�z��U�Ǩ@�˛��G��ɰe�@�ac1Ǌo����ˈ۱�~R *�_w㹋�͎����O>�mJ�����W�JO�m������C0�[-��t�!.�0K���5� ����9�m	�A�J}:v�~�oh�HIS�T9�?j���/[�g�PL�8;[5w���PaEa�x&�0�r�W[���Ս����l��rO���pf�We�}����K%��e����yJL����!���j}y�X�o{@_*�;�կ>���ɇ偰�g�L��7�H���.�tI-��Y��9��+e�C�j$#7�#;��ך��p�������*�}M�|l�_��xK{�'� ��	\\C[����%��݈>Ǝb`�@c0����?��ZF��7ed�0��`���������l��~�� ?S3�GC�A��l ��)���xޤ��!AY�۫#�vw6�*t瞿�\N�����3ǔE�m��3{4)y��Y�Q��Y��/��:Y������(�c2��1�$�l�A�92����f�g��&K�ѻ�kD���|f=CCZ�G�y���+�B���e:���1pG�
o��W���g�;�����7�Z�ф�<�5�p����!�M���*�{3L`x��dCC{má��������� 0<5�K��ZaU��ސ�7K̾)5%�����=���,P1�P�f�a���r0z�-�@ �W�}�X:t�b�Suu��?��	�>��O{�+�(�K��T����M��]����6��@��9vYӐ�m�����$A ��t/c]N_pض��])n����W8������`%�6����=������d�����n]!�u)է콎P�������3���v�5��t��Q��Kb֦8z�}�׻@|'&�䶎ĶVJ1���g�sPuΦ�U�|~s��P@�x��z?�?/}��.���~"��c_4RP��� (�|q�p��Fk𥉟�_�0��ǭv�#�O4��,���N�B�E�W����h��uw�0:�^��Y�1��T0�[d��ŦM@
X��k�a��SU���"��@��%��tn�
������A���G#""�5fD�{��_��CdQ:������
��
� ���ӷwɖ��c���,��D�3����aW�C´^0�02�ӯ�%���ֈE����i�1�O���^�m֜1k6�5X���Q���FQI�2SE)2�$��/�I&�)�9��xE�%�ޤ�;ON��D�̡�(�Ib��%<b�M����������p�`�F�l�{���	���G}'�f��9�E�X�	<��ؖrIc�_���+���m�+S�y�z�sy2{�J��TnΩy�����i�����4��B�HX�$��=�"��g��r߿ �x�,�\Wc���$,���a�Ծ9o&�W�r�%S�/��#.M, ��o-��}�o��Ȑ��j�0��T����<�ҕz���b�(,�� >)j�
��
�}�3��n�L�o��Z��k�<ֺa3�H�fH�2%���Y&��f)P�.�*���DPf�;�wsU��#1��|�؝ۓQ� R&�Us*�7Frv@b��:���6��3"7���H�`k����m���$jƞ }�Έ���?�Z)����#y�iξ�r��}fa ��]elK�ue3c�}�b �]���P/�Ֆ�����Ҋ�{���%0�ii)���}��E��;��9�+W�meXX�z�>p�<b�:q�|q�%v�~%�5s��{���ƙ��[[�#���U�_2�����$���i�$�n~�~64'3�:a3�����M��ʕ���(Y��*9�!/V������_���
�⽕� \ON<�d�� 7��Y/8^�L�n��	�//=�"_ؕ̖��8�R'8��x�Z*=ݙs�_�F�> +G�N�-���N�.v�L�����d���ʓgOk�>���ie����A����?��[
�7����[Y��ٲ����{aN`�d�����)X��f�`�1���]G���'5�&+)�:62a��[o.=�:(xp�[v��^�5Ǡ�l��@�� ���V�����-JB?wn�?{�1�L'�{&:��� ���_�5�p|,D֥9��Ρ�T+�K�[U�|�����hS�"3���������R����B)�5D�#�m1BS��ȎB�������ooH��mX*pQ�N�'\)iϪcd���>ܓk�&X�Z��ַ���%��r�W�傫�~w(Q͜�W�CX�t__�|�Ubbf3��C�����76��T	fK�Ef�`;c�]��Y�e���'1�	��������aw),����})��ks����,"�+��fMg�I}�i1[��ck�`JZ2���1{N���9V�u�:Q&yH�'ih�7��������g���8M���(?,?�*X�0�Bp��4-y�U�ND���D��Ḳ�/nC{L��y�D>DF壆
�������?��em^޷v.�	\5��'S{��^ȓGPز��E:5&��4u³6��=c`����!��9��F�Q�@ "�H��!y��t#��I�=�>��ٵV�hˑ�Yf�{ն�Ͼ���e�?��rPpB-����r�x�3T~�����f,9���W#i�ELU��e4�<hX%?"�p���+/eoަ��BiȣWƋ9콁� �É͖<�ð��{76��2�����$r��ʯn���V���2Y��C�n�kAwj﷗������r\��=�����A�#�c�ж�P�Ơ�"R.����>��v�g�YT�k�2��b�M}me��4����-ibv0F�%������@x�WS���T��俑i��I���Aǎ6f�].;4����o��03���*Q�R�J.ua�G�Zp���lM��n�S�Є�/�Pw��|��;t��b��;"ȉz�9�r;�6�}2*���wS�p�G)'� �㬜xEڪ��݁ߩ��Ho�&T����"�ƭ�!�&f��b |('=��&���1�fZG?�)�,6ӝ`�Ek�J^����1>ah?���I�����Qn�[�䝢a�0�٧��"ߝ�x}8�rl���DW�=|-E�
��?FLhzs\�d I15C>UCڠ���$��F��j�� �:Ϸ|"��4�L�6�E���t]A���:���,.w�('�^D�'�
*R���	�8i��l����)B{�����)��%��9E#�SҠ?���5��Βnf�L�"\��jy�vi��D�H�}؃���x1��C^kZ)�)-�ٱ)T��qtp��I��i���(���Q�*����nAj��VZ��-���������;�l���	��V� �!��,>����pr�� �^˦�� �yY�)���!����@�{����y�0�P���]��g��D�b��/��/�7�g-�,�F�;#�1�����B4�ԙAv1�5*=ƶ�a���CTN��b″$��6��G{�|2N���f�I����TY���P��E?��{�=Q�@��q��O��{��֥h@�!�>��Eq�s��'eɈ��d��uW����)Zfd�/���V:tFEqZCǙ̡}�_m�%9���H����Y�6���N
"�:O��[|�����op�
�� 8p#��>zn�	q���,�����������u+���-�P�T1�M���i��������[_���lĈ���	��]B	��&LGRj�*ޓ5��r]�0Z60h�<WN�k;8�o�\��{%�擛���c���Y��	a֝:�(���烣P=]���5kky�.CO�3+��C~�`�ƃ�X����������	�2�x�!"nG����k]�!�$-=�� �Q�Jy�X�V*
Ol[�/��*�4�-tp#͔�%���@(-5�����ʎ3:�"CJ����䵛�bN�3�Q"�9�#��얇� �����4�3�fVX9�6x��䨣�Ȗ+���S�u&[�\��c�+��ii|�;���-E_%��4
��Q5��r���C�����c�28Jr�X]ѷ�̖���Ё��ax�
6(K{��
�KT���Щ�܃�����\�~���HwV��U�0�tt��""�É���:�9M@k�:��q��sj���_D�F��cF����ǘʹj� <{h�����7�" �q4r�[��������5p݅P��Ҡ����_�"��k�,�	h�t�P�=���C�"$Qr8u����0#Y.Z�x�]p������TY/=���|�"
H����?�=N���?�Y.��f4m�T-0�i����ᇼ�9"N#L�b�D�p?��t_?��6ϣ�K�����44JV$C������a�(�� ��/�cm�_�p˗�7���r�����Y�y[M
,�i�����{�Bo�;��d:_������9C�a��DIڣ�d2I�"㔁�Av��9�*G�i�i0*Ù���y��G�Eg]@� �t(1g���G��	m�P��n���K�nبP�:���Gi����DR�Knp�f���>��}`��1�H?�^����R�I=vB	�7V������@�
l	�O#��Q���A��O��=�����qi�����^S-�)�d��S1V78V��������T/�2�l��(�s��d�
5G�O_�rr��<K�iC���S����gi�ڵ����"�W+��� +����lt�#��
����;�����8&'�O�\v�B&[��hs�k��I9�;��op���e��GR��bxAjolث��↼I�^�Y:X�Х-�Y��'=����&�C���~��*����a�v��B�o�-0��L=E^c����"�C�$��I��r區��d'� Q?�)��n�v������8�<,���*��� @���KF73�+fv��y7����P���E׷�͑)��b�1�&����a�0B�FJ#�}ۨr�a�8� pX�����em�.���[#��e)?��MbGO�&|!܏q���m�M3l��i��O=U¢��`9�����
պ"2V�a��Ӿ�?�c��Lb%�&�3,`;8,�A�\1�Z1<��s�*��><bo���km���o9��7wEU�=B'�g�.6Yt?g�@�u�r��������~y����ʭR��bթ&�u�z�rR!�8@{��/C��n����|�Fs�v&��wƝ�/�H��N��U`Y�,_��%|�"o̝���D��z�y��Z P�\�^}�5���5�=Z�0��S*���',�A��z51U|]��O��,��>W�<}U�j@h��l^�"���l��Z����U��M�k���B�.&:4�_�м#\%���곘N3�������T��]O�e���h�0h}�;���H���'@���{��\�-�������~o�t!Z"�����kM�n}[�a�����c�䓷�$@����f��BX�,�/߯��r)����u�h�E��6�ԿڡD�|t=�AOx��*Kt�ٲ�T$ԯ���r;���a�V�{���J��kx�9�}�	��^���8���c���7�����]���IO3�@��e�M��+N���PK   ﴵXJ%z�� �� /   images/596a7037-fb63-4077-b806-d059e7ba626d.png "@ݿ�PNG

   IHDR  v  >   �U;d   sRGB ���   gAMA  ���a   	pHYs  �  ��o�d  ��IDATx^���e�U���9tuN��h4�	!���`�`l��~���ُ�~�}�{�[6`c�C<L�DPi�43��$M��Ωr�����o���9�֭ꪞ�̀��W�}v\{��{�}�=��+��O��v����Z���?k�Z_��U.�ᚧ��֔��:::���::��I�0�y��Y䵵FX5������C"x<��"�jE�ΔI�ɥ��u�I?ed9�U�5����.��Z]��պ�kַ</������k֭����ɸ�khME���XWW������Ғuww�IWiNT�N]]]��.�-����#a�$�j�p��ą�ʶ��ю��pq��'��*�&��E#��W*^�h%��+!�ԩ6���Z�^��U���c]�4�V���u�ZW������J�����#�IҁJ�/�+\[Y^���Y��x����L��Ԥ�j5�_X���y������_Q�Z=�U��"�e���5�.����^n6�E���G��6�R��21�гb]ZI��X�|[SVȯ��llǄ�;p����j�\+622b]��Q��	5�n9��Fȁ�)i��Wx[����缉yNi�3!��˨�)mM�C/u�c�-K�����YSb���d��S���5���9�7�\�i!�>��<�q�>P�Y���twZ��B�{)����+�A�ݩQ;��y��$z�k�5ڭp���q(H��Хs�Ĺ����ӆ�r��VS�^_�. )o���$Uv P��g�/[>/O
�A7[����
;��[��seٹ[`�#��V7��lu}*PO"r��G�ԟ1Q�4�,~ !�������k�E�>�rK� \/E�^sQf�Z(W���(b\7s��W�T��%m�nr�K{qo;@.`X^^��,�e�@N�� o����r5:@��4�BȨ�ܪ�&О�x��fgm��d�����Ң۫���A�萀rP���O���1�b���Vz%K�fZ���rV_{=b�w�uVޮ��KZ4��6�p��"!�JǨJ �K~�@pŖ����688d}}}�M��p˱*�s,��o#�9E�w�bl����	�6�"�� T���^�W�uPUB_��ȤgI��Uo_E�$�IU���e�B��2p�Ox}�8��"L@/&��U9����}Y��r��>G���4���F�Ţ�:�_�{ۥ����)s�.=t]���ՐI�+5W	�r	���#�0�Z��Iհ���P�t��6��̃�zXp��/Gm��)����b�����Xw���ĩׁ��	�"�u޳"k]��,k`�� �Gg&AHM�ԉ����X����_]���2�-ʧ/�� �+�Q����)|E8�wSx�� ʯkP%���/t����b}��{r����+9`��Ů��V�e��zM [a�c�u0v�1�� ���OOټ�s�u���쌐s��줡�$���W�J�L(l��_�H�j�E���!=�6P9�)�v!������N#`�;_�Xw#��,X��;�ꫯ���!۽g�[oO�묧�7Ԫ\����S�X�y�'{�^B;�H�1|J&�ɲ�֠�B^�p'L�6�/��;�:�*  NL^\ cI��]N��_-'�[������NW���dG�bet�2l�!�F�	ړg^_���'o����u��z�W2��)❕��ڻ��]L J�կ�Ef�Qa�A*j]T*J5,i�tM���D�t�K��/*F=�����@�[P�|8�D�һu������Z���^�Uލ�^_�~�{O}Y�![0�S�^���0L|$�~d�[R�hC����J�lExC�:�іB4��Qn�-�H�2b9)0��}�<�cQ1.��)`]{X�� 9ֹ��i��䧘w.�2��w�xw��YW_�u��n;�tfj� T���ҫ�_�җ�e�,��t07+�s`�,�H�-�:��C�^u���Ẇ0v�I)k��@Tgn�C{�$�z�.��<.`d.�1�vP�M�����;x��GFGmbb�����oZȑ���KY,��h�����WՇ[���-	�ǿ�Mvq�Q�����JQW��,�e��X�N1��'���J� ����O~���|�U��0��r��. +���0��&�S�[���)�4��C2���h�\�oN�\ѶГ9���n"���H�-a�3Ɠ�v]w���bg��Δ'RPPs�UR񅯤h#?�.�9����_���Ƽs"�W�\���_yܯ���9A�u�����Z]���X�U޻�(P���yIav�~�L��'�J1��A�2���ry<@"�I.Z�k��?��)��NX�'�όԁ��'�|�E�J��� ���tV��X�<;���9��.�> ��5�9��w���L#qC���CyU�/�꣥�i�/����:��>kkKK�+�(0�����l8���أ��{ Q �}��*�OzBhW��K{;��^U$��>
�y�>�K�ў����]{�����؈�߿�� uɄ��]�r����4j��<�_�%
p�_�"k�_�ϵ��0qӢ���.�}������j��:��W���!�1/"Ml���)fy9*�;�>���֫�zN��c/y��#o2e+YA~Ֆs~��M���4e����ǜ.�-��O�U��������*"���n&l/0�	��_���UC�u�5��{����m�w��i�rܧr���p�X��[�����t�<�G���0�P�5 ���R�۳�l=����fWV����*��������x8�DX)8*����R��?����$��m�a�<"K^�_���L��'Uy;\.]�dY�c���<���k�MS�[�%ͶL�.�Rz���t�*��}D@$ˑ*C�輦|�2�v��º4;�{��E��c���k����T*}X0�{��!+z����}񽺋�� o��M�<�Z��c�&,����2aa��>�V:���2�,����8�O��a��#�clL`'��#�Ɣ�R(	�pJ�<}Ƶ�D�Xx[�H�}��r]��F��W�qݏHE�H�MO�c�𻅍�qu ���?�*-q����"�9Aר&@=��Gn����I</e1��L$vy���q���oS&k��9�y0I
Z��
;y�E~���D`�U�A�'�����wq� '�w.-���-y�R7�e�������_.��F^�*���^���*�p,JK&��A>8�#_Ga>���.�z�T�j��rDwa�w���t��5���q�P�#��Y�\o�"d�Ü]��-�)��T�gX���t	��zn)SDi�s�9�>w'�N�>NЕRҷ�#6\T�}}� �z�9�À=V_�V�.<䏽��o�+�9V7�y�����}��X�sf���9/��P�@w�P���+���+@�U��vi�E�eY����\���<�Q��<ήw/�0��K]C��1`��~����6�s��������ط�z�!��9E��#�zuu��;��E߇oԍ��Q;��i"���a�g)�7�Xd3.�p����u��.�"cK����.�3_��q}^���(��=r��g/=�|P��e��Y��/�<���)�G�Or�$r7؋����[堢͓�YĦ�NT2{��;��<
��nskݑ���:��O߽V��|qk���0��"�mtZAM�^�c`���Rj��RaP��-��_�(k}x^7�#�ŹDh6�$�x��5T��zӠ�U���[�^M?��k\ �^��:��V=�/-��wI� I>������'��O��$��dj��nK�l��9�B���ɫ>���.ޔV-��erC9<�z1��.EZN�@�N�.`d��햺�<��8 [)U��.����a�__ᎲK:� Q��]=���P��^uųY�K���Y-�+���/��:=}����\�5'
�|�\X��[��cz�4X����vTy8������w�z���,���k�*�P���l�cX{����پ�{�k��;a;G�ld�����5�K�Ղ�.-*K�U��裟W��w��z�]{�K�e/������"�1}�/�T�W)���!����ŵR�.Ɖ\�A_�H7.�o/�<>�H/<p�O���e�.��?s���߯���@s�#;�,��7��������J�Q�Y0���վ�#���1Y�����q����FS'o�'�nm�{@��qfr����D�^Q��
��ր�H����v��]��׹�s�H���&ik�Ls\���`��n�e��A���&��;�,*_� x��?�{��zH�����#M9�H�9���AQ^�X�Y�v��}� Ђ��[">>T�\�qn�p6�	��S1O�_�΋�9�s�K�~&|���u��	 �~ �g���59\f�Aݔ��Z�/�P�s�p�̚�E���O�&[0�����_hr� ��1DxY���|����I��y-���(g@k�h ��� z�h1m����>�E�����'�oC�61>n�js���=�y螵�ǿ`K�n��SR�,�>��ڃ6?_��-�v~�ۮ��s�n۽w��v�D����b\e�BU?���V����%�'��"]�k?���"�x����N�����>&S���ё�ț�!~{�����SN��u�l@��H�HG�Q�>��u6��񲩏v{`�B?�=��J'��0=ܫ��*`�w1y�<�
�Q��p/�%N1����U�Ͱp���{"4<�w�A��A��9;e��ޯ)��y��n�ݭ	�'=u
�*�����	<��AJ!���A��%���/�H��}ʘ�$.y�yJ�O`����4��Իd, ,�J����5���H�|2��"V��`�K>�0��.��0K=��������u���>�&�J�	W�u\bRw�L(�<V���MP��"}'e&n)���dT���]f�0�|��\~\�(��������X�F��s���w(��$�/:lpt�:�F��l��}��N{��lx`І��t�8kO<�a;��ÖgO(��vL����<����:햛���e�ܱÎ���=��O�������۾��T_��ܹ���N	�CG1�X<�n��a�V�=��iNO����C�aG&Q���г�1���4`a����JW��Ma�A���*�$U��R��؂�ԍ�mD���*Uˍ2Bw!��u��F���(3�i�=���(g�Ǵ���-��b+F��=�`H�[�� �V^���D��jTMU���=�f�NÛʐ�;��"�2E�ݜ/�|<X�r1��=����8��V{GY�=���pqT��{z�'���Vw!2)���z=���t��E��$�f�|ϰ�.R�t!9��B�\�]�^�Ex�
�8g���W���2��������E����J�����0��#�K�J�@���T���2��A�z;e;�zq+��� �䖐JXY���zWV�EF,s�f���/S�Gn~����;���^Y�kjyYK�������ŋ~��/I���=�s|��M�������u��km�[�;g�]k�c|���++������m����g���>{�،���>b˫�v�m����뤺^�#�rK�WaI���F��=Pu�tq�D��O�~-�D���F�J�?��4��(�9��D�g����c�-�D��y�Ou[1��v�`@��D]���J��ғ�E�ԟ���-��*[��З���C?�凾੕|]׼�k���C�E�v�+tc9	�S���6�+򵆓��i\�2�w�^���c�P��z�~�E���r@�O��t�;����;�c)0M��c�G����.A������"�cBD�F3 �����U_�K)eJ+�s��a����t���̲R)��k����V��`�J>ϋ�8Y���ߍ�-�̺@b_Lz�Q<�j��[���`��'��]�J�������
4��(��E�[ֽ��C�;괻#�L(���_����W��1��˻4F�����=]bN�tۀ@�4��=~�P���!]H��x�Ν>n��[[��;n��n��{�-�؝7��8;c�����I�͞���S6�%#�c^ctN�OIB���{e��۞�}���=�ۃ?.��T����i:���c�kQ9FZI�+}S_���4!���#�G���N�,�S��Ʃ�4���XQF���ﴂ2��M6%�;��� �|��q�17d,�5.�q]%�HSR������H��Ro3�,�E.�-�Ő�ر��)L�B�����䂪�6�krnx\��"m5}����i�6��uv��-H�� �UB=-W�U��A���'w@���	�:�/ ��Og 1��R�敆�`[3���L�I,�;��0��)�-�PA��ۤÚ",`-�p��l���j� s{�>͉�i��g��.�&-��,�SX�+\eq���_Q:_ �(�:�+΀'!�'~��	��=�Э���T68�ư�R��z\*�?�S���J��m
S ������|p ���ĉ�:ހ|W�@^�!�@��޾n���^�Uho_����}:X��$$�0y�f�fmfv�&'/ȝR55�Z}٦Ν��'�ڱ'�����Y�����Wgmv�r([w��s�70n��[\�ξ]��6d�s�����ڎ;mO>��={������1r��[Z�~r{��N" ��?���Pn�<]���p�%c��ÔI^BI�+y��h��.�ղ��1��r���Z�8���7��Mp���o�D�Yo+�~����LW�-���`LnJ����*O!����]�����Z�%�
���7Y�,.���J)#�Z�nU^�ۻ��y�7�0I\�5�n�yx���f\� �2)8p_������Wg�V ��:���Ez~�B}�Ȁ�����n��jW����S^�J��[�����!�\�C����.���S�x������jk� cp�}��E��I��^�2�{��k���.�����oEq���0�]���%RK�Bg4�}U��~;xsM�b��x�s�&����KE��q�F�h�]����B��,��]v�^������F�������~��Y�k���R_���Ѐ�S5+6y��\�h�Ϝ�E^�������)�_�p�N�9k�5�C�yר���E�m�lx�z�=d�..���n����c��۞y�Y灾>����U�J�:p��&^.M����e�������z�^~�}(�T��$������A�uԇ��G�^_q���u��u�~�C!c{r
"�F�ee��	��(�� ���?]R/�.����"��+��i���	(t�xx��	uY ~�A���0�~TN����2��^%1':�j�z��V�i�5��kHm��V����7@�-q�kp�~���
YY�~I��,@_��X�~HSX����( �q��Io<LtţG'@+B����`�Ї���_�V�O�UV�"-mw_"Y� ��҂���z.���@�l�ot�m�!�}��% �7����J�6C�h��j� �K����X0t�P���e�w蓉pKN��2�C�珁 u�A�K��~�iݯ:�����T��B�*���h2�]�φ��x���-��ʞ>~�>��Oh�eY嫌u��7٤��M-�L۾ݻm�Ȑ�*߷{�N����!��C���,��5��}��Ю�l�g��;�lA�ϑ���1[\�$O�=�'���/������m�����W�ʾ��ou]I��B���}�4E���u�9�<��!s��sP���]Q�g�Р�u���J9"6�/��q��y;�1�Ři{9>�Ԛ���y"m�	'�n�\z~�,�ǖS�� b�^��Uz��X��u�]_Ӱ���!E�t���*J��s�4�H�^Q��8�Z��Ni�S?A��zE���k/��=���bx����~�4@�_�g�W���'�J���<a]�ҙWus-v?J}A.o��v���KJ���+*���S�5VP:8����&Etl,\u�m�����*���S�~���e5<VAj��.W�^�����WxG
��~t����-ܞ�{��S��_P|1�BI}�YW�������r��ǜ�E$�z���^z�AQ��%E?y�U㮈/҄��WF4��;%Z����Ҳ]P�<s����c�����[�Lr�t�krj�fggU:_���7=3g3sK��eK�.L[��ޱֿ��8p�M���>aKk��X�a�vu�8�s�뮷G}�.\�`;wN��¼-/.ڈ�={v�-2BT�
X�bQ��Z-d0�8%���1k�9���	���MW�=]\��Mq�>�� ��_$(��U+C!n�3�y�".��9K�I���-�����%m�U�F�h�����8Oz1�#'��TՑ�՟b�z>�o���~m��ϟ���Sn��HAg�p���:I�H'�@�ƥ�x"&k�jV���g�L�Y;ʑ?��Ƶ�|ay��"�����9����'wH��H}���}~[��"d�k�S/�Sg2e%��A�$T��*wl��֐) ��.���v v���\^����N@GFY��L��h+�s�"�k+���>�R�>���E���~7�V�N�=n���&�ϴS��(��V��@a����}�mP���|����ٴC�����q��]�� �Gq*�C�Ýt�pG�O�#@� s���䔝8s֞=uڏ?��>/]sR"�h�D�,�pI��=t����hAc�d�޽���=�v�M7ݠը��L�b��!����S����_R�y�!#��,x��i��>������k�g�^;'�X8o������ɱ���G"�����ؠ�����v�M=D����{�(�w���}C`�X�pj�
�rЋr=}Z̅�noN���ǸeR�-�6�#�������I���V���&*t鵭/o#�������:�Bl9UY�&�JxǗ��w��h���i{tv�WP�����6��U�(�=dAQ`/��F��cm��ԇ5Q��싚B�R[�TLN!����S��D�bSvt��R+���]l;8uIڭ�[������{o�R�:^T��/�Y}IV��8x	�C�溒�����=�ت��*��,X��E�
�/<tc��#���~���F����u����[NHJ����2����ܑ>)�(	抱_��B�*/Wwm��	a�.����>k��_p�_��lfYV��h�(	e��������>-����~��v�mv��a���P��f���w������b��$�4e���0�300h�e�������K���o�*o����u�گ�*���VR+�B��7��3���]#�o��0V<��ND������V����B�ŗ�3��q��li�]Q>T1�D���o�2��l��*8B�:�ZJYSP�Eۣ��n����}��*O�(����,�mYO��B��2G��ɿ_���j� �P�w6nш�oTY�3�\BE����֎Ke�`o�,�����6�@A�́}Y�v���pm�Fk�
 U���V��x �˫ ��ū�(�(�%t)��:d�ͷ�䇵P��*���Z�u�b�����U/!���v�[�����l0���b���(ގ�i�\�!�����џ����������J�r<J��u�ER�K(\tr���V�m�P%?�e���ɐ�n�X�N9�+u���^Y��$�a5��B;5;+��3gO��ӧmv~��k,�ca��Ȗ]�9:�Q��ٹ�v���Po��������
��ԯ� Jm�����{��|�իl���|����(t}[K :95m���K�l�Ξ���%��7�u����#v��~ߞ�w��u[���ӥwk�wb4g亟p�[}�,d�j���E�S�T����(�B�{�f�L�A��o�r�
�u��S.�P�;!���z��CQ>��Rm"6��6�&��L���(�1^���.��:ӧ��'V�m=��L��)T��T�@GQ[\C]W��k�坦��k�������rR�'/��پh��F@P^���[>Pc�y[ˁJe�r�Ug{X�Q�_�.�t�C}@3�t�-�/��h�p��'��)���M1@���!���J���ɽEeP�2E��/\�	��u�����זt����(�|I\�Z\[e�Gنѕo�,/�K���p�#OՐ���*@��\+>�f|��BŻ�ặ`F��^'~�I� �\�Qɾ��u�2�ˣ���_�*�p	s�~O�ty�uW�p�㾨��&� G�J��ih�:�k}�� e�`��#O��3�����������)�UsO�@�U�����s�Gؿ�n��V�������3�C�&�ó���p�Q���^�;:4h���gb���e����a�ذ�������5�/�u'�}FwoK6}q�.�;k�����lin��ϯ�������~-�A����>���3[F���vY��naldȆ%/2R�.sg�U.mgZ�z5��+�N a�s+��~/��O�.�����.�c��r^3���	/ ޱ���kb=�.s� SQB�����׉i�?[`���q��i�Ў*���q�]��?�SkX�{l�IPH����-�DY���vTAc�H�k�C�kN�����R�B���
�恩�akK��>�I:R[��ڜ�c�w��[����{�L`՛��U|B$�P�%(�[��![�
����uP+n�˯4|�ӷe4��j~�ӫ�a!���Zvmn�Vd�����)����Cw�\��T�֕:�ۑ�KY����T�%��u�"������ �!��bL�p
�;��G�o��<��Ex�M7ƚ��N=����|EAJ�jQeۢJtӭ�Tcrb�ֆ�lraA�?�|����'��:�e�`�����
nMwOo�!$�Dk�5۽{����/��q���aۻk��@C��A�e!Q��������2<��i�ߧ�a��N>[&�W~@����˹09c��_����m���3^���c?�����Mo��N�x�=iT���(/t\�	��0�:G.?俇�߿o*y�����_�.�a�^z\$L��ES�;m��Wq�Ϙ
9�=�D }��/$c����i��O�fV5��R�M@��2�/�T�Jr�wc�a��F�v����<��$�[�i�)��p+�z��꿫_�5�bl�:�s���)¹���z#.��It�<P��D�P��Z�XSX�faI%�C���L�?0k,{��wP�?N�_��n���J�[ |������yg:�`03 ujY�������.�zp�R�K<@O�+��:�� -H�����0��]��߅cp ��4�3.9�������8ɸF��Q���d�ٙ<&����D����Y`�+/��~�SV�?��_��a�^Ş���Zq
�C&嫎� �(�w��	�zA��d�9j=��}�9z�_	�ȉ#���e�Y����oIW��W|���G�پ��즛n�QY���ڡ�A]ۈ,�1�ćd	���>:��V�NY���Z$U���qW~^����
��-����=�����O�5����{�i�Yw	W_}�U���ئ�X����T�����/�s�����sW��m��������+���C�[=~d����c�����o�o�|�|����\ޗ�8r��q�� �jo�+���yV��Z�p�H���:���0�#-��]%�A��2�O���J�2��)Ra��r㭙 �k��]���A�č5t=��u;��д�	��I�W)��_W޴�E �r`�O�:�����)c�lN���n\�&q"fpE֯`�w��`�\�R�?��+��)sˍ.F#�q�D��`
`_��2pK�KfQ���t͹�v�� :�o7)	`�/:��� ��,|��/_�Г�:|�ɅB��ǠwXn t .@OZ�Q7,?����{0~�
F��1�bd�d���rݯ@�yP/:">��u��4�\�P�O$(�/�E��F���ㄘ&��V��wY�ǟ=a�&����6u�--,��\�t@�Z~��\�$}�����Fl׎	������.Ӫ��qp�-�a�%�����~۵s���1��A��;:8 ����"���N�U?=�C��0@�������ߩ���?w挟��:?��u���� �6?�c�;:?ʋ*բ)z�lQ�5~�G._tp�?��gY}=�Zl|Ѣ,�Dx�����Q}�_��0��.�[���U������p�u��%L��z������ו�P�M�w�d��E��,7�R�nP/�6�����2�E���~�>��5_�.:�_`���j��2]����)�`/C�~�oę��WE�E�@E��{�rU�
'�+�$G� ��8�k౿ާ�:$+hP0�.7��-��]��+���� �$(؁J�"����a�V���"�c�ϋy@ʗ�I��0g�9��]@#������S��	%�ɖG-%�/���-�1h�/�Y������gRRܯ�
V�u�M:Xu�4u����pK=�S/�J?.e��˥�\8b����/7d)�J8�����;�����}r���T�C��`���V�
������ry@�6[/h�&�"�-��Ps6��=&�m@��/����6���lߞ�v��W۵��C���z���~�j���,~�Ie�jh�Z4z��!@S�߽����(�Q���Rck��=�������v��#���Q;��tݵ�~Pwt���/��Y8�F�@��hQ�������\zq�Q��嚟���豝�ó��y϶��-���lq��2��2�� ��{E�1B���^���,��q�-�j���Vf��J��,�J�0�G�^�g��'V�E:��*E%��\Dw��근0���-��L�޷�$��E�ui�9���:�nu���.���:*�z�c�dX�e:eq���g@z�5a�1��Wgib�:r(~�Ad�~��	@5�L]ǰ�rV ��?��_)�X�<]�Sn�ғ�-v�ٖ���i��Jyʏ�~�+QV�a��l1�:�ڎ��ʫrc��~�dZ�ÿ�w�T�������ה�=g�9��Gz�|]�O�I�Q.w�}A����"\���<�V��ɜJI]�BE���գ�0���J���3�d��=����-
D^�M.-���g����ڱs���ܔ�5`�5���r�J�2��nimE���!�������u�}���[�z�����QY��v��>�{b̆��5y����U�x;K�-��E�*l�x�U�\5A>2o���)�"���ٸ��E�i�8q�A������c�?f��CWV�kۼjxՖ��bݕ�=u�)�8rcWjc�����cK��R�8�z@I����ŖV�`_��,�%S���Y�]�J:��/��do3%z'3���q�x���D/��`�T��3ڤ���N����X ���B��E$�}��8��%������0�A�������!�$,��2�<��[��֨�t3U�*�x�d�P�ҭQ��Qw<���U�iʰ�\#,���%��_ջ�d�k6��h|��K��ӭ`:K�����l_��T5�eqY��� (4���UE��Be����ZZH�πV����4VP�!��ױ�(<X��>�ۣI��{��]@@���6jѵ�bи̺n2]���k��X��Ol�j? � #5.�-b��.����)��x��D}�.���j3��vV %h&z8a�"�r�]ѺF;�K�}z�k�� KwI��}����SOٳg�ک��mj~��Iz޻�`�V ~�,N����cW_u���e/��~�ou�*���Yo��ůq95�;���*���h�H.d�Mh'��I#��rG{�L����Ӻ��M__��x�;�ʊH��ss|��f���g�~���}���/�k�}�������뚝9s�h�F���[ �V$�hx�����}~�����G�闐=d�Y\|���{�:9��$y��b�97iӳs653o�˶X[���-8��,|�)�vh�]>e�I���*Uqc#�� �<�Q�md�x�=\�p�͌���i(7����Qv�'�a��t���b�x߫�p�_����^��;?��k����@1�^e���S����+��-�+��k ʌs�V w�6�<[[^vw;�ڐ}�/�m����j����p�jC���e��cR�vo
�Hd@�� ������~|�{�O��娣�����X�� 0���z��uk��n�MJ��+�Jʟ�Sz�jDlc�>�'1pI�.p�s���!�PLV�l� �~f��Nق OaL?��>����X�I
1��o���OX�,C �E*)�
����+�E]���݂�{9>^d�s�/����䤝���#�N���Y��g��w �/�� p���tQ[��>;t��/�ݻvځ�{d��y��;T�7de�`��	B��+��IA�s�Hzmĕ��j�q�:=3�8?���|xq���e���Ԝ;'n�9j��?�c��bx�;�{�G��?�����>���ި*d�^�������Q[/��!^yN�Kw"�CC���v����9���	�O��l�9�u�j�v�������E���>{ў=u^֝Aw�:pW��v@^�++?�mc<��"MRs�P��{ʬ��F�RN��p��qKn֣���O�!I�12�_Q��J,��ё�E�!�S����,�Q�u����յuN�p�r��VU�V���L:�vT�$)� �.���`���+�� ��|�Ig�A��ѹ��ȎD%�q�9�����/��Xy�� ap���a�GdX�E��� ��`��%p�KOkw�ũ�{�����r��Ԥ���J�iY�J�q�����`,`�_.K+�Cz�ҁ9r}kK���R|˫�+�_���xXI�amiQ�5�O�};ĜA��b��)G`�}@�X��Jϣ��6��p3�B,J>�����:a��6��X<���� �æ�18�cSSSҭ�Շ����z���[쫿��lyq�8�B��o]S�⤉�G>�3���UB:�����MJ�o�5��B^��4��$����|�{���F̡�,]�S�#Xu`�����������}�#���^�u<go��/������wلUػ}ܧ����}����{���ޞ8�>1>����Sbu��5}
F`2���m.�p�\�OڑgOk�t�-N�p�>V�|��������ӥo�;HJ+j�/C�s��������y��)�F\FhR�� �%����*�凼\e�>p4�B���7�x��B�M�ҩ:�Wn�V(��N>(-��.��N99a��%���^&�.��uj�2��橾�s����⩯	��/��V��'(Vi��_���!~�N��M?��9x�+�-����� ���b?v��jN!��r���ZHH?!�����1�XU� rK'CY����.�Im���+ �X~:9��r���C��,/�HV��>�`�R��!�����`
"\�7f���-�L~E3=
��t�aER� �ӧ����vV�v��Y;v�Y-@]:t�~WF�k�~W��5��.߾�_j��7��풕>>:j}�~�/>
�=�~���g����9��PC�=����F�8`ޯrO�<e�<� ��?����0�w {·�!�U�V��v����t�����{���Zf�&�x��8`��-�,�&�(�a��A��Ǵs�o�����GJ��}�Q����T�@�_��P���n]��ٖ���Ý mg�Ĉ˨��Y�s�m~y�N
�/N���h�j��<�1�����\C.�¨#��J��|!�ʔ��Tm��Qep��(���AD�IG70h�>d�^�3O$_��ė����>�c�$���o�џ�q+�S���g-�(�*ԥ�lL�Kޘ֗&ryNi4�v���~p����:X].2�|���>Q?�3;4��\�N`'>n�qprs`� ���؋�7p��¨)#����O)
 '0�:�󑛴~�AZ�� %��G�n�89@���R�jw7&���fM &@ٿrb��4w���% 7m������������Ô�0��!M��\WJ�[_DS��`��=���ɤ� ;{�\N����x?n'Ξ��S����ÊTY*����=�Պ��	��w�]w�־�k��n��V�M��J����K�us�,��!r���I 0�z2ה.~�_���y���ܝu���EzV��X*�ˊ�>S^���c�y^�[�����ه�GRs������#���bgdپ�o�M���C��!��5�#L`'4��>�Xs�Т8�'�J�g�8��9׾kׄ,�A?�ޫ0����$y�;-n3��n�bq�fu��9�~�"�0U;}�0�U�bqc3�[q�3�P�a���'(ǵ�x��!��ɝ����j�q�U��'�����}�d��G�,?�f�|�A\D��#���x�G>�Ư��+��ED�m��_�H們�$o5��AQ^�σ���)�N�o��*:W�r�,>��SV1@�ߖ��S;1tN�`�������RQ��5�N�(�ݘD�	p����"W�z�\��O�����i��R0p|�� ������$��ϣ>�|^��U��sT�b�Գ\���&c�3�W���	q���V�|�F���F��k�A���� ������}���y�1;?y�&�K�̝���X��{������]�S'gR&@�}�w~����שO:m�⤀j@�oE,�r^�}�G��#�n�.;ܐ���;�n�� �E^���oh� 0_Z�C(l���[_��^ ;��	"1�z��qB��"3�:�� 	?)�|,�J*�>l�؟ٯ���j'N������7����Ν;]n��E���j���⥻�������"��rM�5[kJ���1�;^r{���)^;��d��h�@�-��sai��5?�����=}���n�� �k���t��R{�;��OTRĺA ��v�
ɱ������BW�=ג����Z��HJ��cQUuK	��5"U��YN�����k��7���	QpRkC7"R%{9ECB�[#�K�}�g۠L޺g��� ��l��:�?�*���d/S�깦D(���߁K��s��oP���+tH���I��a}(�;=���ML�G�"Ep31as�FY%�\1qT�
$e�1�}�LXn�ƙe@5�L�j�0�u|˧(?R�BA��\�a�3��� 0�W��E� �PZH�a��<=>6fG�>b�����>h�Ϝ�m������*�/��H�-/̙�Y1Y���;l�{�k�[����nUښՖ8���8�ف�V٢��IFq�3��ڄ��Sj?^��f~K�f�v��W �J�r�e�[C��q. H� ��7d˪�;4��7��ū{��~Վ;jS�SƋ���k��k�+��+lalH�{U���i�����_x^ =�h�� ��C�c|T���G�G��}O��q���ϓ���Zk+,b��JG'N�u`��uW3/9݌� h��ÅB���Ѕ���A�F_��	����^92BDX�+X���+B�͔%�K*�C!�+I���Z����~BwΚ�E"�*4��G�Ʉ�l\u{
9bb�9��lM_y��5�ME����/�>�[���6���0%��B�<�FYA��a��y�������`/?c| ��*ȷa��l�<��U�����2s�G}q�V$��*���sA��B��b{�p,�2:�*%M3eܒ,A��o�ّ�����6 ���Q�?��?�O~�v��9;ἀ[ȭ^���, ;?���\��!����$��_~����^z����![�����9�S�b���z\�@�U�4�8��Ƭ	�|�[r���rF˝kb��Wj�^�Oub��r0�l�aP/���Y�7�����>䵾<��>���j��˿�P���₽�5������o�����96�Y���P��P]��B��}!�J�t�;a����C`�g�w�������؃��������@?���)Y�K�e{��i�85S���T���<܅:�����9nbn�+�T)�@!哮��q�<��:��~�K�<q�L�\��.u����捓�(�lm�u�0��>�[�^�����9�V��l���Q�d�U��;=^WE�mPl��U@"�Y�(�I�������R�%�6tL�A�I� �Z	S����B^|���@R�2���T_1��,�]�H�XDH�)E� �+	Y+u)o V!�+�$����L��,ݷ^��tl��qm~a9(�X�-��;e���9��G>�!�%�o���Dqc۠Kj^�>h�����x��[o��&vN �[�l�`�
T�8ɂ��S��K���& h���Qє?A�k�P���EE� �|B��2o�G���5Ҫ/<��Rzd� ?�������;���O:��`�r�-��������i�@�/h*\���]?n�&�6ǥ!���r��V��d�*o���L
�w����̾E��$��Cb�����<���E-�|�N�N�St��[u_�En'!�咱��cMg�c�BY R3���(ʇr����������.���w�,S�OJq������J.PQ�$��o.jC�}/C���}�ʎ���O��\z/|N��)�訚
���u�q�?�iؙ�'���A����m ���?���V",���(1����D|�����Ԑ"%�<e�%)���dh%����W8�E��??�=66��?e?��}���G�K��e�fgfd|�����ܱb5Y��jFG��}�k�[����u |�.���\��Vx�:�T���.8�$�I&Y�:��P����_����a�q�[%��s|�6�0�߃������B?��g�3��_����+5۳g�}��~��[mdd�N�>w&o�b�O �'�z�ߟHf����5���B&����A~tP~?�.%�@��J��+�p��.�_n�7�����������ѝF�&�9�Ţ'�Nrb�3�B�BZ����������T�񸐛k�7�~چ.�Fy����}�A<.e��Ɵ�I���B'�A���6@X��D�a�����@\�����W^��:E�h�+��a�u���֛��*�����V;���	YM������R����b����ˎ�Qv~�[D�$E�ܞ 9	�I����>�5OP�K�L�T�kN��(�����zT8.Ƈ�S=ٶЏt�����9�����������yĦf��}���^��Z���Ȁ��C�E��5���#��Z{˗�e/{ɭ�c�n	'��J��6�J ���Af�@s��a�:�� ;x}pbϘ��,4��{�hE��a�P�I���<����zy�|X�r����C�~@>E��#G����������j8%�_���ַ�U:�g�}�5v����!�F�^ra��@��'��| �_�N~�,Zٖ���C�̻��� x��S���j�>3��/��3+���������,n�\�y' _�K_��+⠲� ���VXX��H�|elf^�C+�E8�JE���j��,�J��'��P���0u��Rh���	ZRC��"��"C�@U!���Ǖ{��N����W֙���}D����eW��Q�)�0��OHv���i�V�e�d/�(����P��p}��?���%�VS8܊�!CP3x��[t���Z�*�R�NXqY�c�"C��]�p�Ξ=+�:b�����=(P�V�؟��Z�\:'������������^z�}׷�]{��՗����h0���1&�滻s?�)? �E�6~���N�'�-�8�Ÿ# ���芮��%1& ͺr�j��`��!�R��o���������a����y�}�w}�۹��t����(�g)�nA�D�/�1�2�<'�]6�x��΀�l��c2��(������-.:��
�o�_N��W􅟺*d��'�[ �"܁V�	
9IwQ�pw"�<r]�މ!_�_�n��2!���8�~��y[�]�{�0������ �ŕ��{!H�O0hoc�6$�u�����)�D�f�<�!Cv~Pi_�"�E�Z�v��p�K궨%����uT;�ѷ�����*�))����Q�E=A�s}�Uj�W�N��1��OJ�gV�}��g��;�k'/���I�5e�+M@���J�|=_��a,��~������W�y��w�b[^�6G�l�HϪ0����HXF�,q��"���au�cɇ��*/n���JKA	��i�Ÿ�R�T��D=Yw�=v����wۉ���@�]w�u����v�����������8D��*�E�Y������a� :�R��=��S����R��`�W���[/ydo�d��uF-���4��̜- ���+i�WimƯP��~����H��p��u���)��ׅ��5 :��Ej�A�wO������/]��e�l{e}��- ع��f�Hqy��z"��`O����PmD���O_Y���,������z�B^�r���/E1�"�:�e�P���U?�fx�6�RV���?�ov�L��5+	.eU��\v^���,{����x-�����3��߰�?��	����'OZ�,x������◣�(����+��/|�ۿ¾�+�b_�/�� tʌ�_�J� `���cs+��B��Qq��l��`(�$��6Wٶ ����Uu�1�mN�f�(��|���4J��k�y���x�}�3��_���-��-��_�uj�A��aT�OP�V�'�I(�n�ʃ."�E����Ti��, F�����������$#mA� p�#��e&�HL�{}��.cF~�]�"�]�����lM�V���q�Pt^SOX�"oc���2�\⑁���r����V��}��U��B!��&`o4�[��p3.�
UH����U /�E�v����b�Eck�E�M�I	�D�,���A�2�n�oRs> *�@W��V��>���r�#c+�o�r�@Y>R'�^7S֌��zE�Ź�ks��&�D����-�'%'Q��W�X�?�3?m�=�������+���L(M!���#v������y�]��7�ew���61>g�Un�M�[z,+�9�u�)�����ޮ[鈫��� ���D�� BP�.�G�vzR*oSr5_r{�q������������}�׽�u�����\��=G3U��Q���[֗��f����?��iu�z4/��y6���,��<�X���ss~j��S}{~��Vu@8)�~+��)�3��MD�h/v�Dޯ��&JA�.S��M�0�dq�i�"=c�A���VP�+�?�V@���)
&�J	Ϣcp�n+}�����$�V����_EY���ۧ\X\A��\�|��'��*����Uj�[�a�U;j�o��_��C�უ(%������5�z�$������2V�?�YL%����_~�\�|���������_���d��t�.���؆�a'�ҙ�a�_��/���{�z��f����E�ƳO�X�G(���<�A([3�H�P�gT�M���g�&6��t~w�US�RQf��(]s�(g�2���5?=t���ٟ�l�ٳ�v옰�����n�=N�4�Nk�J�F�v;T;�4SsPhÉ*�?�3�-���������%�t/����,�qQ�C�}̸R�Z��駀���<�hC��)��R�w_�<�~�j����LEX+ex�0���_�+�/`���:�N:�:��D"�K2w%@�0
����lA� �*x�5��[���gb[���eÞ;����D&e�ſ�))�UɯЛ��S������ϰ�F\ᇪa��Z��sL��.9N:�rk��2+?.�m�8&��N������P�E�I�.�=���H�o��o��3<$�A. �5rMr�(Ψ�uu��#�7��[����/m���J��𹲦[�����Wd��Kx}����f�g��zO|�F�`��I'���뙸`)�� *ؘQ��t������R�L���[o��������ǩ���POB�/��
�㧟䖱�)�%X)J��Yu)V7ʍ;%��x(���,k�=xY�i�6�,**ְ�q�m�$�2����M��1�0��9�ϸ��j��K���Qn�����.>3X�jW���1�b�.�O��@/�H���5��5-�!��8'�S�O�b�U*'p3�gX��?�ۑ��<����f�kܭ1L�q_��J�ϸ'���F��'�Y�&���yЬ�Ojk$�[����t%�u5�S�k;��?ケ�n� �2�J)C��uc�z����◓�O����I���>�"�A���� ��#��5�4I� ˋfw�v���[�Q��?������y����E�Ea�ͻJ�;�S 9�Λ6u{M~��E�O�h�(�8�D ��k:�vM��|g�,�=el�i�#�a�`��cS�M8t�ǹ�b8p��}D�X��ټ��E��1���TՔ�7�o�iC������f����b~�������m�w��}�B���'ex�a�\���5,Ót�߹H�q�yJ,�o��hi��KW�׷� �"�����d���o��AKP�ʆ���Ki�7�qA鯆��i���$�m��Ά�ŕ�%��/�ſ(����\��0��J��ne(]���*ex5��uR��j�s�MK�q.6ۡ��1�c.�]���[bX�ra�����=��U{��g|q���5���O�nX�;�w�ٗ�u���o�����{��n}�}���#��h=XZ���,.��΃9,F@&�SO���TD>���󟁊��J�>7�u\^�K
�T9�X��B䉻� ^5��O/��C�{�P
P
�K��+.�E��BU���s�E&w��>��o���tEZ�ӉK#�m���E����)7��+pC"��{���Y3��b��G�HW5����}��U�9��(#��dN��<EQ���yW*<�a2���oW�5VZ�7�)�c�"vy! ��Ւ<������2
.��U��TD�P/��8B!��:]�ZGr;�Ƶ�I�}A	��˹�ߌ#��N〱�֠g�j��^��i��'>n����o��n߆!�" 5e3f�<���^�ҵW�o��7�?�'����׸u3}qRcEV7�@���\�:`��4m�z��6 �ogc
_P���7Yh��8�T�Qó��"�㔆���|�I;~����ht|�n���׶똿��店��O�BQf�E=��~'�.9qGG��?�x�A���{&_��!G��[�0�3�F=���Lo��SW���:���D�x�O)
7�hߞ��v�/�"�g����Q��
e�� |yK{��+��",y3*��B�V�_���<�.�[�]�Z����^i[�J�CU7�Q�ͶBq],*~]�sQ��˼�Bհv�q[��<�ɻe{�{��;s�l�7M�)Y�G�<�{�ı�2��t/̞z0{�u���>�ll�����W�~����W����a�л���_��R�u�kn�rԓ�(�Z����}f]��
ǘ`ll��:\���6`g��2 �ʡc�}���~���|����o��J�n0
S<,Z�7�*������!��(-r�؞�|��q㯀����3�W%�4tXaC���>-8q/�B�����Í���=g�଻�qD��ۗUe��j\��/��V����*�A�e4�F�Q6���u��)/���e�9ɶ�U.�N���v��Q�ގġV�F�2��.]Rk���������Jj��ap��f������я~Ԏ<�����7��//��)��--N�~���������U�������飶|������^�����F�-�v�?H-p1����RW[��'I��� c<�`kܥ||�h�#��0 ���������Y��q_�$���^��'R�oƛm�a��_�����x6��	�[�����x8�z�IyM�u}�2Q���]�7����E:ڟ����y[�<y+���Ve�C)kT�np�U��l)�F%y�+�U�ך�5l3��o�i��f�eD��ܪ��S٪�VM�`�EPR5T-�5��@�x �z�,.9�/��ڎ��K����|������ߡ~��I�֙h�{,�Ֆ����4�|Y�������O�����Mq*A^7���D�w����:݂}ۅ��l��g�:����H��s�����4��_��&�J�g�r����[n�n��ffg���7�Zxd+����屽���m,]t1.}��a����_\X҂�R�Q���R�|�8�v��W�u��G�j:﯂��jXkX���^R�LVwq�Q#)Õkr{�W�Pd�� �L7c|e�ۚ�Jy/�[�]]����'e���[�_��|W��=\�(��f�8���?���c?�c������d=r4/o�y;#�B��?:Z^�_���������{��;�֛�3���;ܗ5�I���W����N���k�~�ׁ]� �A�i���/0�7��#[��8�
7�'d��I�H7�$m¤Q�8�ht��8�`;&��I���eN�>u��A��٭� M�։k�qۥj��Q>~��?e�x�N2��Ug��Eɮ�\J[-����r\i*u��2n�Mm�BK���I����u�R ⒓���V(�:�n�����-)�.�bNE�1P�����������l��]���ɕz���v��1��?`����ӟ��=q z��jU�\��eYߋ�;1v�~�������n�A`5��k�W-k�,|c����KAt��/�Z+�G+�J���A�^�
0B9��qY �6��T�+E����6e��9�D{8����W_m;'��jS|���9�9��/��+3(��)WʩR:[M0���� p�ś+y�;���-/���ޤ0ַ����D��-�GΓ%ϥ��V�g%��6nrR���P5�v��N�-�<�;��[@��~�C�+.��Bюf�Զ�ok����qu�pa/����������������Ka�+�@�cE�9ʨ|!L������oz���k�Η���wu�*}���[V��9X�	��ūZr�ݥ�L�9~u�K�V/���&�@����=����6Ӆ�����v��A���
Exڠ􇛋S�n�ۥ�v�����q�6DQ�Ҹ���\�rQOP����P��*o��F0D��r��K����}���"�v�JU![)�m[ Q���7n�U�:?n�6ks��`O��C��U��*ex�ٌ3�F�ڷa�T�G��j#���5;~�������}�>��O�ɓ��|?����M�+@_��_=�	�W���ۿ���;��N;�2��6�g���עaؗd��V�8#of�%��(F� �����H��9S�?�U.t2���7%e���pP�ez�18Qr�7��'��Ҫ%oԟ�ae�o�h[��q��q\ ���z/\0��OPO�3>9�
�/m�搼�?�a���N@����T��f;�%������i�)��r��?3�����1��J;���[�,�}�|_h�q�������S�'=�;:WuMM�V��:�f3;tp��o����w~�7[mn��w�+��u.+�3���+R���U��/
ؗx��.�������S���U�o�V�>fTKR΅�0%��K��'��v�7cy�Z�O���꫾�ݹ9�	����rDY�a�Dٌ�8��H#��_� uC>�`����(�m��m;o)U̟`�n�փ2}3w��Vv�[�U�vqϕ��W�K��X��M���[�ꂘT�ƥU�Z÷��J�ŵRky���)�W[e(@|�`���[0@B:~X��{.���{�o��=?�����x��2�̺��%�o����?�����p�k��++5�8U�[�0�9`>��\�������.��\:K@^��H5V؁<��6D{^8�0v[�`�\�E�?!9����x�ZMwE>��3T��D�5|sj��%c2�)��%�Z� �8��?m'��t�A�\n��Fxj߾�Fȷy]�$$m+{KS�c���K�4UjM���e<_T��|� `:�>����yX��r�_\Cqlp�&&v:��S?�Sv��9����������7�z�̾�;�`����/��F�la~ηm4�m O���-���WV��z�U���H}�'at���< v��÷0�n���3�C1�=���cO�$�n�u�pLot��?Tڱc��,Eo@iҧ�?�A��"�R��}� �t��&�"�c�=X�m�#/�����&U�'��])J��Q�EgI�r�����s{R��"�O�"m��D�/țS��fir���������nN�\�uG�7{����N4�����#�4r�}�䔍��������������=�e7�|�[h� �7����%[�髼��-^��;�V$O]�*y�@99��K��HҮV��*�����x�\���6`U��,%е��L��5/ÿY�I�ۈ2?�[�n`"]V)?�Q=��[2\{���z>\J7�9T䃢䒿��hw��hkuQl���z=��"A�P1����V�*e����1�&�K�b���I�5��^�,;�/��{��R�Ϛ�i�U�����=��>,M9Lֺ��LP�n�����׿���6u��|_�����5��Ҳ��ٽ�=�ea2�`�����%�8P��CƮ��h3B���C	ʩ��rӿ�8�%�Ģ���?~��YY��n?me@��.�����HW��R8�������C~�c��J��A��hN~]p;J9q7�*�ukx+�����2*�w7�3��R��k���U��8�\.U�l�v��]
}���>�:�������P�����i�x.����}�4�Ϗ4�wII� u�/�P��S��o�F�����j5���ܜ���*�A�V�*���]���$^�+����UU�^�?�QkRضeh{ι�n�n�J=^����
�X�8��m ���섳X����}Z(�x�WF�n�����B�VBf�OW�RҒ���[���K���B��-��6Dh�F�M�J��t�Ukٸ<-���lRyƤb6��^�������_�C�b�e@�8?4:�G?��#��ڒ&$'_( +����7�͞�_���ڿ��ܺ��O����B��]�RzYܫ��fߘw7vk�b}�>n�%V��GN��!\��ܖ�v����� �E@n��n��Hm�v�_^aL?qݫE�E�����J�m�b���CaU�RP����g;H���A��:ڑ�g�[�"O;����ׅ�Z]l
���
��4��I���
7���W��}I���r�7�[ፉ:���];mn~������_�o��S��eW�-�.6�ժd`dk��>5{��M���?������>X����:�����`��b�@��*[��x���2�\� `����]��n���Tυ�����p�t�b`�����$ʝ����q*����s�,c���ynT�M���)ҒY�;��ǘf�Z/c<�J#��R��^��z]���F�����o�:�a����S�O���z%�jX;j�X���%������-e:\���	3C�2b����ĸ�Ԋu
�����{�/>�vϽ�����m��Q���*�A]r�j 15��p������V�?��/m��	?=3�7(@g}��.⯛�-�m���ut�^��{��sC�	�;�e�%���]���>��	�'��C����l��߲���������e�˿�����d��*��C^�v�m��m�|��y�u�TfEω[p�3(Sȗ۸T�j��R���]_lbӗ��G\s����s�v���؈���m�����1�V:LXs�e���Í��O�����##~N�豣�������{졇����[򀺱�-@��}�V[2{����v������ku����ɋs6?�D�kK�.[XZ���e�����ǈ�4,u�t@T-�
O0��Q�.�*ؖ_T����8�M.�"�������ܣ�W._P�y�{��
�� X�C^?	�@N?��}�ƵbS;P.1`c�����v)�6�k#��:��(7�q���% ��+AB�MF���~��`�X2��_�K�s�>j��TXu��	�׾~�S���?a�ȇ��y���`�n����Y�F$�&�y��k^y���w�~�����aCã��7bS�5[X��*_V�|���G|�,��U^�%`�4����:�@x���՗P���Y[�1G����p�����K��K����Ǒ�;���P��T��Ș@�V;?p�lAlÄ��\�
�oD��(��e��^�T�nm�:]�0�Mv��By�_x+��l��S�=��weYC޿������[P	ʹ�+u�S5e2~�}#�v��A���ٟ�}�C648���=��_�&sFH˞z�/��ӓ*ke�~�_�_�������~��y/���>[Y��b�j����0��;�����P��ۦ>����Ծ�S���(o���,�oɢo�9���ۡ��<��p�<I�(�ӥ6�v�T��p�Fe�CX�]e�V)��P��z��KP�h��V�R�t*�C�[���� m� �!���UX��G&�v�4�Qt7|BIw
|! �}���_����/��}����mffZq��a~���Rwk�OU������&��_�/��W�����lM��Ã�>Q�
�*����Rr��u�X��ޫ..��`��#��S�&i�h��^�`C�֖������Çل�u�H�Z-�d(J�"��S u��� ���.��:�!T�I9F���0e�ވ��f��pO�.��b/�?�	_-*�T�Ɣiʲ���Jeu]'���G!���*zo�j�����]Ǚa�~���'��O�u>�644(�RnLF��'��]ᛤK�e��2�~���|����;T�,��);w��-.,j\
����"oe�[[�������h��0�� ��Ĺ�mĤm7���I�-��:C����|Zy��cG���3^��_g;���]u"g�Ѫ,�^oޮKQٞ��đ�C���H8�7�����p?���v)�����h;�z��Ͳ���4t!��^u��v�{)*���[	���n��NO�8/~j޻��|(�/��s����R��^�@����g�g������g�5-���>�F�*g�يa�l�J��������훭ol�֦\vN��!βSgJXrH�a��|��� >r���1�G׌�b2(�i$ތ�2�K1v\Ȇ����D�[e�7[gh��S�����tQ����6�c\wU+~]�6�.}t�&J�I-o���N���;�ϸ䊣�((�y�����2��6���+y��U%T�w5*��	Y�KŶ�͈zʺP2+�(���vq��-RUw[��Z�g�'��$P��(%�4
���~pVYL�L��������~���O|����rr@����C0?0������x���w~��������W��lq�lIV|7{�Ա�_5�J�#����62Wo\GT�K[V�����xh�RW%ho�W�R����N9xi�ɓ'�'���:��648�n��LP��6�/c�Y�n�!_��"�]�����y�j��R�U�̱?Wʹ�|���it��V�KN��[�+s{u%�Us苛����bs���I�B�ׁZ��c� p�ui��-�'�����b<�C#��''���O�g~�g퓟������Svs$��.��''��o|���-o����e���&4�U~|������5�_X�}y��ίT�[x3z�_�@+(@�gچ?����^.��/�W�r��.u����?9}��a���!��D����+Cяp�wU�֬����zy��QB6�Zg�� Ѕ�_��� _�A;~1��
"�7b}gq�Z'U�ϙZW�\@Z��B�IY����Iه��X�	@�ı�O�>%��Y���V7���3�{���)��W�����٧?�Y뗵���ۏ�%�wwk𫺁�^��^�ڲ�?��?b?��_�ַ}����ҙs�w��xP�D����\:�0嗦LZucqJ�=UP�/��G�+
���sb�?����x��^ �\`a��������w��ܹ����)�kܭ�ߌ�d(�X�(�n��*�S�ц2m��V� A �>�����LQ�
5NBE��Qn�Y	�-����p5n���m����RE��Z;?r�[ q%�z9�Bٹ�m��L�|s����ba��6 �`���%�m��=~����&}��r�1��£������{�����ǿ`{���W���(��,@��ڭ�/�����;��v�Kn��i]*�����_y�T]|!�w�/���\U��p���ֻ����'�7�?M`4A�h0Q�ě�#CiQ���U��<IbE�*�_��5|t����}�1T �U�|e[���L�t��7ab\�N=��[��p^Sץ �4ț[0����������(�G�k��I�$���ƨZ�y�9�R�E`ß�=
���eD��Kty -�
� d���(���~�ͯ@�����m��cn�3�B��.&�ޡ���}��ʯ�����gǟ9�[2��sV[��W���On�I;N��%�u��������bo����ؾ��/����	�
[0��K�%�v���&e�ƃvH��۔�c���	��9�X�m�!��}1�T&�^���Vj�q	~.T�*�o��#j~!���C��2�|�����\:U�~�{Cj��]�����9����2	P�6
	<�%����ƺ|��q�=���+o�T��>x4���)A=��ͩ��V�V���V ������b�P�U�������#v����m��n��NYB�v��}W�/k���;44�&����M����?�5s��>(:�:}&�����2�xY��J���&�_��w�-o�r�J��OQ����fT��To���	ol��|��u�y��4nUDU���?p�P�wG�!h�G�A?�{](<���Z#����9q��
�	��y,���C�O��O��Ӄث_�j���AO�sw�q�҈_��On�P�w�J�`�ӭbR��&x9b�ī��e����������Yb���X�7��2��emd��v�1���xǻZA�;��蓸ʐ��Ԛ�3�e]M�e�m�+A��t%iM�8ړO>i����{�̤�ȟ��{�Y�̧?c�v�k������Kئa���石_��߰#O���^��α��뮀�Z���5�V����~���}�W���v�ָa�`�����T�,�e,,���v� ZK��y%�� �O�c���`��C��)]�ŅwC�o;~�P�%��j/E�d]@�S�~��i���|D��[�w�y��x�M�����i#)���U+y��k�8��~��~��btԹ�H��x���LГ�v��e=��h��i[cRnϷi�e�rkR5S��
�o`Vn���]J�K��!����W=�5�0����-�C?j�����?���O��fO<����~����������/��[���c����k���#K�[x����65�{b���5������}���+�)���9U#pg�I(y9	�����Ż��פn�k�(���Ү|�z���2<�`eqK���_g��-g����nґ�o�b�U'�V�r`N+=i�Vu�s���{�h��k�qw�Tn�뢔%�"�N;Y�T�c6��W��+;�ù}�cʸK�v��^+'eT9i�w�[����^]�R�M܈+<�A�S��k'��~y��KOm�r9T�_���308`�܉��������_�̺�5a��l``�\>���v���ɩi�#��}���������a��!u���UϮݻltl��m�ۿž�������[�KB���'� b�A^�+a��	ؗ��l��d��#�!�58�=�#M s�g�PO�X':n���A�U)tV���@�o���~z]�~�g?k�����?��}�+_i{��)�u$o�<m��e��т�������������9���.��e��G�z!.GIͺi.��iJה��L����*Ǩ���+D�oe����]B�<�)��=��1[�]-�\��NY U@��ݼޖm���62>a�?y�~�~���k�n���A���ށ���~8?@����]�llt������ȸ���������#�5_�mv��wخ�n��WY��N��A	X�W;%K��t��~	Pg�ähK�|2������M%O&�jQ�����W���5W���g"t���}��,�',��r��b�_![{lø|��z�yA������ϭ�A)o2�l�Xq٦�%�_T�RJI�"�u̗�!�L5I���5q�y_^�x��~�i{����v��NY#v� S{�<��]� ������>����[x����~�s�O���d���������k'�>kS���>��^3Y���0�d��u�_�$ww����)�\[��l<��M�F^��5L}��Km%�P��ou������؆����1����߶�k��[2ύB��E��M��1G��X�9��C~�Q��c��E�
]l�W�(R�W.����{�S1�����;a��W�/��Z��h�=�%�����%��0o�CCv��q������{(�hވ�&�}�7#j�t�Q1�<\�N�Ly��AE���c������
5F�$��ԗ�%�<Ʈ��ڿ�.�;c��=võ�ؗ��۝w���?0d�.N�Ï<f#��G�w�)&(����>�:����4U���yh�8&��j!�F�Z&��)F\����yM[&?�QPDۥ�͗���K�I�P����������?{��?�#?���ia6���y�=R_ec�m'i.��d��LE{b\u�L�r�����q��y*�ᣂ1��W)�Y���Z�]�U����}_���r�D�7�����'��.:ן��oc��r�t��K��=�O�?~���=����ȕ���S;=� �%������6&\]) � w@��D��o1)����{{�41�]�������N���/��ؘ�zǝ��kv���6:6a��m�����{�-7�����o`�'�,4� �s`�5&u��P\mY�N��ʠ���>��Jp�M`/�|lom,V��V'c1���|�� ;D����>�A�o������v�UWُ���g�?ٿ�\ޘB�1Bh�z�;�9����v�����(�1��~�&����� ;�k'ӥ�{9}V�sky���MO}@W8�b��r3L�~�FE�)�nDMeC��՗�B�'Ɍ����%];wN��>�9{��\�L6�����xȭ�.���~a|�&P͖�d�ů� h �&��gE�_er
�?ٖ�M�K�u[�g"�JM̵n[Z6��Y��Ϟ�g����Ssv��y{��3��#�ڽ��o���g����|�{�I���a`��w��/ڃ?l�CZ F��v���М����_��෫�:U)�m$waۻ?����d�t�m��"�����u�{�U_��c�(�g>�Yݝ��;�_�����Ȩ/� ����mIP�l�,��܁y={���, u�/��b�1�r�z�#/q�`�D������S�Ԯ����Amϱ'ex�%�'q�!�1�]L��ֺ�6�%j&tꖷ/�p���C��kSN>�{Ͻ6(˗���W��<�G^Yi��
nGlppL�h��断�oL�w�0\�`�6�H���bn�$�)����D%��>~��a3��v��[�w����>+띗}���*^����%;w�;q�~�1���>f���_��_���Ҝ����3(��~��iQ��P��1��A^~�h�U,&N��^o�9��cS�D�s7����7��[-���ElA���|�:Eyp����;���Q;��3��O}Jz��g'��]~�)JE�\��וRo$}	����h��_����� �9�!�G_��v7�JB����O=��zm�?�BQS���Җu���|W�ߐ�a����*����$|#�6�%
j���{�lI��H����l~~���O��_#��|B�W^&���r^\����.M���s������%Y۽�X�J�I�Pv �ϖ� �(�i���m����y;w���m߾�6�c�t�r]֗�~�[�.�&|��U\k���+����dU�E݊?{����g����3�q�'>�I��O�9�eW���y��o�,�V����c� ���`�2&�Lm�8�?��<���#����?�Q���r�-��c�l�,�����ӂy�����=gc����7��b�ZB{��HQ�RQ�Wm[Ÿ�ܛ��Q�g~�ĳN��2�ƅ���0(rI�z�.w�<��+����sV�<��B!e��KЖu����%�b�iv9Ԛwòh�6�%*��U�oLt��윃�����Ye|�hqa���	�>)�E��@s�^ﰁ�Q��E;`/��Uv���M^�UXQ�J�;�t��a�dq)���]]���vvn�n��&����w������;_f/{�+���svqj����. ~���r@Vۚ&7[0��;� ��&��,�%Y��n���Y;?9esj���g쁇��ʎ={B�����{��&v�31������-2��b��8�1�\��yˡ���-W�zXmm��U(��1>ػ>{��s�=vR������򔭘}����U�&�y=�nKʞ�n_�x�˝V�k�s��;+��������h�M�rG��j�)}�ݨ=_���\�6Es`��jӨ\����Ԛ�R��Ó���\�}�)�c+���)8�������������Y��'�>w��A��w���4�׭eX��Xm���622f�\s�}������';e/�f\�FU���W1��_�fXH�0 �=���%�������wԼ��o�����vP}�'m^�O��*��l%"ʂ��
Pp����ag��KaɌ��ԬM�/۹�i{�g��Ԝ���o����>Y�5����3�����u�~A���/k]&Y��)��\!m������*sD4��o\�1
��A�������_��:�K����>;y�?{���855�c~�[�b;w��c��I*@�ǿ��&��d�RʻQ|I��"���\C�]��;+���a�W�!]�7�q(�i�v����[�m6aC`o�f��Ӏ��F�����s��)��G��ۘ7��>E ;�_�����{��G��x��t ԓp�\Ba_`�u?#�h.��3�����X}������؛��mdx���SUߊ��3�8s�F9X`<�c2>��3����}Hqv�-�ح������C�W�S?jyr��b����'���d{+tU���X��� ���W}��t����>l���~������*���%�ѻ?n�������������(N�9c'N���O�ɳg|߿���es]*t�ʍũd�������#�LNP1��oRy%l�X�y��#�>j���g�:fێ#�o��7پ}���}x/�!Ws])��s��j\�t��6�Bx���r�*\��u.�	G1�3�¤�H�j6���AQs�7�-'��
�y�!�~�Mt�ne-۬m��*���������pk�U����O}������6���)���l���������۟�����MoX����<���/����5N%W�mf�n˵Y�/�׾�k��;_��u���&k��=�Ƚ��������5�������u���/��u�c|L�+� �t� ƒ_i���[�:����ۚ��C��v� �&B�Ϸ��j��n;��ܵ��cll�]8�q��׾�v��O}�n[���-Ν�5-@,*otxHm����۽k�_o���m����3��_s����g�{��;�}{���H� hY��\�+�d����-���'	�:��4�"m�>�~/�E"5ϻ��n?aT��ٳǟ����������/�c+���8TpE�f��g�,��&�꼲"���[��28Vjn�0v�!;�2n[�R^���=e���V�e{��O�{;��N,v����R��]����bЋ؟oyJ��S�ƤSGj��ea���w��m�Ν�����v���س�v���=n��Ƅ��@����c�W�z}^�t��h�?p�}��O�Ҭ۫_�ev��^b/��N��g����{�K�=�kV�"��RY�=n!�Z`�k��ܾ���Ox��6	A��zl��-s�����ES����W:�w���5��(�{���%[���/���֟w���L��w��V���*}��V�v��y{��q;r�=��S�ԓOڣ�<b���=���v��Q.��vX�@�>�;�H{z�������Bf�IK_T�. �D��M*�S�����#o�#�;v�m���/	K��qS��eJs�B|p \Y�? բ�]����wRR�?���>��$c��4SY�I!Ŗe٦��bwB��Y�96�-&��ӕ �+	�ϻ��$Ƅr���'�5�&}�����FN5 �7� x~A��������*�yx0 ��H���A����_&*�66`���'���J�k�N]���	�����z����_%00�����}����`�Sys�g^ei��b��*�a�f��%�U��})��_���?>jBC�<P��O�z�a�<*��w�\��Ҫ��s���F}���+�C}v��)[�ɪV�S'e������W{U&?���X5v�:��֚d��hQZ�խC:W��4��ݥ����_oc��v�UW�Cɱ�Q���g�U}��̸�=>V��g�1�\,��g���Ч�>b�]w����!���q�w��<�V�k�-�:REqߑ�^wk=ݺ+T�覛/��rA�;G��0�XG�)G$��{�qq7�l�vh�y��[��Z���
�P9��o��K��mC���J��*��uh;�NZ~�I�z-~V==;�@ ��: ,�������������� ;�����L���u������>Aa����N}��z�Gf�������^�&�T�����>�ُ��YY�X]�[@�&^��b�&.�ń��&������N�棩2��<����R�)���]�7@D���M,�ښ����M���dXq�tx��.�9)�^��ÒMONŻtT~oW�JP�U`w�@��j��bA���ZH�? t�?֒�J��>�x�q��x����v��<c��v��������bx��5�^+����� 4�>���6��KM ��S�X9���ŏ�؏�M7�ti`�t�7%UT��+�clũo�����ڨ7���.Jc���P� �U��FU��H�97����V�T1����9�CU�a(�*D3Q�ƕ]�R��
�W
̫�bv��\����F�O���{��'|�r��]n����>~������}��G�
���bp/��q��!��k��CK���۫�ï�M����k����^��x�>x��9s\�E�-O
�T����PI6�ݿ��֏�V5��J������Z�x�pLb�+�|�9�G�)�{ђ�����b�������#&�PydhPV�������Y��ر��7�V[�ԥ,���e�Z���9[Z��$]�ݨD���d��q!�Yp���k�!�����#}����M�{�/��m�������W"��ڠ�'�չ|ir�)���7�Ɓ�:y�������O���|�;��0�P�<��O��}l7�m�YLxxL
αWϩ���䨫o�BrϏ�A/��m%_+���_�z�����JM*��^�^����(s3
�t_�U���4����}(���=ҟ���j7�x���c�!?��Ą=�ȣ�����E���"����� �
�j�Ģ�1�#�u+
�BcB��%�1	ϝ?k?��M	�w�
�5��C�k�5Y��h�;���(�ļ ��__�{���2�C���[��?�8���CþM��>__��8��lQ`�IP���x��ԴVr�	?Ƀu��~�tM;���J�><4�7Q�{mx��p�KK�~d�����ĤM^�hSS�6;?�q�ysƜS:�������������V����]R�6S�P�k��II|�A?�γ )�q�qﾽ�Ƞ���k�d��W��_@�=u����"�w8ޙ>�xHZW_D��W�f0�1Ҵ����J��t�,�������6�ܖx>�ۮ U��lIp
��+b�NN�w������O��@���������+z��p��ȷbU��֐���k���۱&��ah�
�:����EM\Y����:) {ʾ��K���Gm|�Ϯ������.��������!{轾��V���K.�w��!�>����Y���G@�)�w�;�BW��,��NX�ض�=l�Ы���p��}�A?P֔�}~¤o�)jn�0\����7c�m���� 01M�� �'k�����*�y-
<�L�l9 ��Q����S�)�������K�X4�Ȳ�#)]�awۡ����븨1�����^�t�m3��5�kׅ��G9Z��*1��1�.%�8&����R�*muk'�V�:6�vqU�7)���3�r����
.G5��i��?�� 7@����,�}=v��Y�����/��O�c�v���8i��'�ĉ�n;v����$�v���R��)�q�6l�6Y�!���9/W
��r_e��U���ngm���g��#O�k�|���O}�.\8�Gw��Y ��:�`�528��Lo�D�>��~w'@[p��`�^�e�E 2_n�wy΀<��Cם, ZL;:�c�b���jg��u�`�9�X呑`��ee�)���_wC��a�ie���L�!'9~��g�?�1{�' c�j��V����S�r��2wPܡ�ĘJ���C~(�����u��+@=󱯟~(�ʪ����I$ߜ[��7ц�+�w��;�n���e��Լi���zY^xz>e�P.�~�u�޶��ey�-t��^{��/��ﶟ���lK����o�7���v�]o�����m����M�^��,�'�{]��w�r��;��J�J�(���u��� 6<Ej��>N��;d�ۢ�ن��]��T+'F��_w�ם�z��]LX���^:��W�j��n�;��j��Vlxx�F�'�}�|�+�=o^�뫔�� ��,-�����ܕ��9��0�o�������xPJy�x1Is,q���O�?.?c �Xw%ʟ2��&�؊b��D2�����%�����o���:y���1�1@{y�= G4��������m!�8~ʾ��j7�p��_�]�t���!t@�����~IOr�.�~� ��:^���~al�5N
��j�����/��t����-�N�+w���ݳ�j�"��-)��t��x���*��)Sօ�Vz�1���6�Zv�ޥ��y����]����-��s�ڎQM��nM��������W��&vL�q�������O?m��_�ﺥ��ri#��@��8��֒��:(�[׿�뿗W�K��h���������E
�%	�`-����u�v�l7��Y��9d�p�U�W��fv���G��Ð�T^��wﳫ��٦kvaj�x�c����E�[����Ҽ��\��/	�~��t8	S�l;'b�Kճ㯮�L�9���ˤ�vC��i=%��������CtxQ.u���{��X�����e/��w�w��KdN��������'Nػe(����+�����?�����v��U�<�L��;q�� k@�kҲ`��P���f��'�aK"���9�������*߂/ːॼhoE�A\GX��p�K��A�kOպ֗��H�ȡ�16���+.6���[������X!��(i�"�F����/5u��(U1!�3����c)dzzʞ�m������.h�a��#���y����{�w}�[=���d��߷���������I���|��JaM�f�q�"L�V���q�LҼv˰�t�#;���AB.��b�[�d˚܋��jku�@���
������;�?8�"��[0b���+��F�֗~��v����'���.�4���ʒ��`vN�p���T�8j�TeX�5�%�QS鍝e>�]�\襕�Ӥj��5k7=0ra�FX�����%�����i&gmt�/�\ ��z ������3.c��{��{�v��Y��W�ھ�o}��mۓ'N�3��G�6�����-"���S�,��ظ�ڽ�n��V�����!,mgABV8�,���|n��������SPY'�?�#9���L�iͽU�R7'R7r(�vh��� � �6T��bɶ�ʹ������b�Wň ܤ��Z@�ϱ�{����f����=�����t?��"����n���Ln-� �߳k��?��/�{��+qk,�ANU�-�1��M��7|A	H�E��_��r�x\�*�)W��Vd�Z�4�_󏳃������3�s֯���;�2�}�N�]�!� i�rw`�D�]��И�|��m��מ=�r8�(`�wqԲ�$@����I��, b;�.� ���=N��yu�!z�x��lgs{Kj���o�F_��!��*�'��>��F�Ms�&V��~6`��m)�o|�}���A��������~'��A	�x����!N�D��6a��|��X��v��ᮻ��n���~Az_��'�����Q��W��W��P��Q��X�#�zI�j����I��6JݜH�ȡ�/$�w��;����ib��-�Ũݠ~�����h"&VL]����׎<������){衇�/���x��11��]���w��n��fM,&���4��ۿmgϝ�IX>�*Ym�:[*�ڝa!aI��8bۧ!,J˒����)ɉ�S�[]@*�;�ݲ�}� ��!ځK9�n�! c=����ޞ>۽w��w����>�jz*����kˋ�'-�l�(��*��>���@�(�T�T���5������?��.j�Y\)t�@\9q�Űņ�����홸��8��(�Î=s���+�1 8e37��[=��Ü���k�����d��B�s&'���ɓ�J���ϛFGu7���%�8��!�R'E���fJD`���و��m�Y9��R�M[,�]�7#��X�}��pR���=?D'����|���ǟ����߱/<����ޱ~�U?���ۼ&ۅs�6<8d}<X�[uMn�U��?49q�O4�p�4Ǌ�%�O�`: �\%�-��*(�TIY>.�UvhR]胉�I/  d�4\|�z
�\v��\]c]�mX��x�����Q�-x�~�op�&e��8����C~T��l4���pa�t�����!��+��!C ��[z��;�t�1�$����ϸ�����k��1��N��|,�X��Irh�}~���_��f��ﵻ�[Ō�y�x�hk�Ϥ�ހ�L.|�
#�fY�9��� �4���2�K]��S1�U!�SUȖ�/%p���y�GU�����]�p�>�a?���������e�b�����%g�1<b�.zַ��mv�-��ׄ��Iă+�8Ϟ>m��[�%kl�jǜ��ӷLcw}B���/%��ﾠM���Y)s=�?�h�����'� �����ûdq��1Dl�x�J'���,�p�+�w��5H\�,v~ �-.�����{�E�l�5^��[ ����`� �c�6D���ԤÂ�+�!|��o���6��B�=;��
��,YT��~i��� j^ Ws0f|������tMe;E�~w"כ%���Gr�6����<uℿ���D{���m$M�:��m�bq���Q�nE�F��q�����@(��({>S_*O���@��l��Q�"������� 	�p~���?g��g~�>w�}6�+�[�Ґ��5/��n:p�Ս�_�޷�.�=c�����e_�Y��s�����K�����L����5�7n��c��?�	y�2��Kŗ���y���
��j�uw�3L�L��ß����j����CNe��ˋ�O΃�85S��\��j`���������;��ű���{X����JXr5�t0��sk� eg��k���"��V@[9�G����e��TU�ߔ_9Ἓ��P"��l-��Ȱ��.���S��~�~�wזj5?��9�Ӡ(j
n�lZ;"�-���a(ܐ�5��Tɳ���mh������Lk��|��>�r�$��F[��Z^�7�L�ߒjd|�������'��[n�ɦd����\��~�f�>[��;VV������Wِ,x^���3��䔿��W�����2/P�$���LT$���o]�z��G��̈�r�)K�'zA�8�Ѷ��f�8�t&��䞾>p*�(�^o�k�a���SYԴS񰘭������%�a�"����� )�Q#zą���^��S�����^�����p���>�P�}f\Սv~qԥ:�^�3��:O�^���nX�j���s��:ˉ��]���?p4��z<ۅ�-)��#O���[n��i,)����V���U�Bŕ|I)�F�}�P��gEx�|�]�^t���Ġb���퓟���x����yr`��h�]�s�u/��CW�W]m#�6$�������sg��iq�γ�E����p᥈��?N�O���!-�LLJ�k���D�I���1���T�1L���qݟ�j�[��
QEQ��j���H�0t�h�v՗�/��vEv�d ����tx[���;+,�/��+�Z��y)� rq�5��z�J���e`!�A����~�ߪ}����J�.o��[����|���"b�R� ��n#Oǂ�0~E��O�=���}K�����^�u�/*u����>���/3mh����v����Z��:.���>,.���ܱ�G�G�o��o�o��o�EY2�������ڪ-O�؁�v��kl����b���n�{^\�-=vR�����g��O|��4���L.&�����uw��'z1q<>ڒm�� O�4��ky7��2�XU6��HWO�,�W��!��А٥�՚ �}rE����=}����g5�)z�ڕ�4���c���@.�s͖W�i��0�+���z��xկ8�	�WMSdr���׎2|����+�J��p5V
�������:�f�UKl��ܥ�R�(��H%Z�~�i{�ߨ�/���W�Q���*�*s#.�\`�D=&��۴���Óo��۔K�W�<��)��C����^C1X�!,&>����۟}�C���}���#�1ܶ��Ό�%몭�5���PW��p���I;yᜍ��m.�*��'����<�I�I(�	�r�~�?��c��uǤ&0�G�p5+Y�����}X�ߘ��ռL��"�y�
�w7�bԳd�q'-���fF�)f�Jďg��i��p�׶��� �Bf�<&�'�K12��H$�C�i�?��V��R��^~�We��p\��+qqR�_�F��� �ʯ+��_��꠮��̺ ����u���S2OY�Q����kߧO�v˜=���Y[���c�(�8~)ϖ���T�`�t/�k)���!���z�^ɷ@ەf��v�\��y�)�&��rq��@�����x�q�R�v��i�<���>y��C��\�#����ol��.���6�<��v�m�ڡ���%坚���?�y{��/8�7�P����':��ᶄT��Px[��u�?�=lK$�4�t�SO���{b�Ȟ[�E�\R7�|[A��_6 ��8@��X����sQ�4j/������'��v�ٷ�~r#�����u�}�a.�8��
tn�Q#^��E���Jw#"���.<qtV�`0з����T����|9D�~�<���.����������?d'O���z�_w�y�ٙY?LZ�C��N�6r�9�݌�)�n�G7�o�<�5��\�jy[�/Y��C�T|�s�?���c�ٱcG�}�w�����[�Z���c�0;��!����^�94��/^�-���_k��z��L촚�y���AM��'O����cQo�) ����K
OXx��䖤���p��GX;*�`#��j�K��ֿ*�����rQ6M�x����:�Qް�����^Y���բPT�?ʇ.(��l^��!`�A4����i����l {F�l Z�����8���,�G� ���-F?P5]5_����E�C��׹\�j��)���~Jj[�{�_鸤�	�ȉ���!�4�W��>�Wp���﷣G������1�QN��G��O�L[��6f�%5t�-�)��
۞^����������D��廥���?�ȟ��\�R��{�{��������QǑ�A�18d=����2�|C�vÝw��k��.~��r��s�Gd��MO�*> J@�ʏs�@�&@����2��"b����@��䬀T����)�6�'�Q�
8NPw `v�Xk\�xj��Cug�e�)N��v�@��3��3�h#�=�a���O3��@������L�+��'٭���q�ny�K��Ro�!/��xª�.,�[�iz�����^�г��EZ��M�^�}�x^�ݝ���ׯ~����-�/��H�y	/&�=4K���={���f��v���FԈφT���J�F����_L�=�ۥ���eW�K?�8z����������������&}���~����=24lgO��E���6��P����}���u�XO|]k�/�`�p�=� KL� '�.� ��ª%�"ol	� �aC�j�\�-N���5��+@.	r!��`a]�CJ�򩠉���i;�F���}�o�nzOo�l�f���� �A~�%�mj͵�5*j�-�m�"K)��d3�N��n=L|���k���k��i���7.����r�#7O�p2��4g���0��Ո�r?������}���p>ڭ1�1_	
�%��f|��[3�Pαt�K�l�`XRpJo��,n�T-�r�_	jWo�\�b�s	```���y���v^�z��[����O�8i��3�?�Qy���I~���8����!���y����?����M|r&G��.�/��թ�a�S�[���h��*A�d�c'����gB�e(G�RP�#/[Ez�E��o�@��o�rdt��	;|`�ط�F��>�Gm M�����V����\�?/+�-8۝���!g�M @��_�Be\�[������}�]"Or�k�b8q������V%ǒb��%��q�r�8�㊫�&��%=�1���p����>����^{���W�h�v�)G+�CU����[���m+�]B�L�W���7����"����i���������ܼ-���U{�Y���@�m^iz�u�����6�R���9�0=i�?��}��{}�=@�UN +����&��,��9��;��]rM63`���[��b,)�r���|�O(�kCq}%�[9	�@{�s�6}H�]��y�נn�F��V���/V��� ��`�������mD�6ˡ(�or/&B�V9�fl�,4����̙3Z�}Qw�W�=�@�<U��0<�H����
fq�� >Q�=닩ʫ2���Hv/�NtFs��<j�'��S�q�>��2��r�f�n#��R������s��b���r�L&<ۖn~t���sn����o��o�����gfl��y{ӫ_k��m�a��=֧~������w�a��tټ����E;?=e�=��=q�j'�L1���u�귘z�/Q��%Pd���gM@��Sp�Bd��:M��$��kqXL%@PG."�Չ�]r������� Ψ�H&~�5��g}"��
1��a�<x8�*��mP�ֱ�q�"�QZ��!-�KYN�-�b�"\�����֦[��Y!˥�����'U˄]�B/�_�^8wο��"]���^��Xgg��Og��EP�Gu�?�v��?�#�1��8��( P��n�Z���}�/>k5�ݚ�O8�8^�_v�긩�� p�2����\�ZF�_~>	��!ѡC햛o�c�����:��-第�AY#O���_x�.�>msS�~�ed�����l���V�(~���,*oA1ib�&�hr�dbg�. �˿��K�����	�'�muj1�]-��NY�\�J绤 zXg��h-�:��ޡ[@�
(��FZ9����ˢb���u���(��[U
���W����Ã�ܕ��_�?Ļ�{�x��-�tsˉA������$�-7@����-0c����J�j��U�D�I�[��R�8�S&�oE�P���rwH~7W,^��;�;��ٳ~�%eC[U��I�:xS��I2 X��!~��A'��ٳ'Oٟ��	;y���.,ْ��&����/����A�R�~�� �l�iN�d�uޑ��C�ѧ�ا?�I��_�{F ����v���SǞ����]8y�l9���=<h�o��F�Y[�%!Ȳ�SG��#G����S�r�:����`��� ��,� \@�&�^�@�\~���˶����^W�<���[޴(�q���r���rKN��.O�����9���<�7O;�y{_�c�Ez�T�,�?k5��G q-�r����67;#�z�?@26>n=}6�k�--�Ȩ�JDv3�*B<�Ix@��I��ԴX�`Դx�K��R���F[W.!�P�{�j�Aq�����v�&y)�и_;�K���a?�©�r�����;_�B\����K��n��v��_ܣBV�x��\��m*�<�q���y�����F�[��w��e���{��Jؠ��RV��J)ǆt��͉�[+ 4�U�^�+�������[0�*b�!;:8r2���ә���K�@�����5�������v��1�0󮉝~��g|̮y�mvnq�Vu�=<d���^��?��pmſT󲗽����ﶷ��v��!;p�*۹w�[�f�O�Y"q��&Vyw�u
8��T~��P:��J��Vp���	'�I����I,+Kr3A!�������/���\�����d0���NJ ����X�b[Z���{{?��ٙI�����e�K�c����ٳ�Ք}n�&k b_|t���N1g���j��U��e��ZS��66ا;��/��Ȓ�֨�NH���6�?��h\S�7NDD���Z�J��[!����B�E%yn��VOW_}�]s�5�����ɓ66:�����⒟��z����}��g>�[1���/y<�t<���P��ǕƗ�FjI����r��\|H�n��֍�/��/�~���)G6�-R��ˣ��Vț�e�^�/Y�W�*`*;:�'"�J�3�y���]��~���k����s���~� �S�.�䅋~�wzi��t���vwQ����	;z�}�/>���}�����߱���+��/�2��a�A[��=_[��yR��u�ZǠ���1��;8d������������gd���*��(����3V<�H5+��@շjdYŖ��5��Ę�=h�*wԅ���grו ����qO���S��݊X[X�.�.@�U���vx� �.���yչl�|��lǎ1۵k�������+vqN����i�\T� �e�_���>�'�Rﱚ��u�Ho��vڎ�A[��	��[O���@Y����9��U���e�Q\_]>�7W��p ��o~��*`?t�,�~��w>��/}28Z�3�Q�%�� y~���E�d1��z :w��CGNƾ�,"�?�ͱ���~�_�S���G �!P� صs���\a ��T��R�6]N'�m-o�x����W��*|�,���<3m�,"�S19��O(tTց;>6f;��}?����?q숝;u��5��P�܌,",�;l���٪,�.Y�K��gd������=����7�կy�M��+w��^���'��ӧ���Ϟ���˶��l��kl�klߡ���ʪ��e��_����n�	�&4��v��9�7�ɪ�����
b�Ƿx:�t�N�3������a{gUw�8��X�>\\a�VL�X4����j�,�좾j}J�"`��_Y���U��o�F-�� �v��)ª�&��A��%7�`�,w��K�|�]���󓳶����dʽ�x�1g�U�,uӢХŢ{m�v�خ�^���cҏt&��������M����X��ȼ��;��JZ(�mD��oG���Q+~�;�x�k�������/�hn�-�={�to�������n�_����5�{�/�x�|ٝv�7�dx�;?FʶR#�2P�˃���0�B?<�y�;=3-��/{��n��P�ȵ5B�xN�N�[!�n���հ����rA	�9����«�r�4�-��P�*�VY�#U�I '@ؿ�a Gd�?08�I�[V�q����o�7���~~�aYH=2^|KC�Э[��^��Ӡ��������W��~@���C�ک3S�D������g�5;'�\ݵ�F�{���6*���m��;md�n�#@�u���{A�4i�XG��{�=�a�Un�,{^�5<1a�##����y)ap�^�W�k}C�3�.��aY���=|��_~��|�7�Mj!���mMh�}��U�e�������������(��Jw7�.��n���)�	�o��Z�.,���ge������7��ˬ>{�^��[l������SZ�jZ<��쒁��`���]�E��Ö�V[p`��t�����w��@���3aW_}�N��`�s�~Z�w��j@�W�7�Ep1@
�2�aUj�[�J���Vj�[��|de��ꫮ_��&��(P�!���8�O�v)&vjHW虭'��{
�[�9�t���+_�
����Jb��:w�`	�߷iT����l��-���P?w��*�=�@�_ '�ř����O�K^kx/AES�H�K��N�ip�F��,�T��������miX��Bg�p<��`��8�����O�ڂ��[�I�w�M<j���)Y��\w�}�7���c��5��i��u;r���Y�M
X�����V����>��e�S�ZX��"gryq���}]�L�P9�Sw��~�
���&5������,ע�ú�'lh�A�۱�j�/�U�jO�u�ZG���d��;d������=|�[�[�uM@^cB
`V�l�z���x�n�?��S�*��)�k^�*���}��|��68�oSS������#ni�����̒�=b���o�c�?`7\{�v��c'N���/ڼ���ѧ>�2�[/B+,�Zm�V؆�/ZGMwuY䋫6&5^�g���)��ӝ̠;q�Μ���G�{�}4�a碿|��Vbe�0.��D�ª�'�E��JY-�Pu�Q��8`;�mD��.7����a�喛m��w(�-,�A��UW_�����o�_Q������@wv��ٽ�t>��Zt/x�����Z(�����{0���jEw��z���a��-#�����ړ$�_:�f䵅�T�|���ԗ܊i�mRk�-m�lB~{��ϭs�y�-�a@^R�"��czO���}���k���s2E�^�����Z�ߵ���_X����WɊ}����&��{��W���I{vrƎ\����v�V�I̜s얱�	�Ȣ�AmM�4=i=�ұ���U4$Y�x�eߒ�@�W�W@޵cºw���}Z4Fl��7Z��n���%z����yY�+��!-;v�b����l_-T��W$�j� ��yd�:,k�˺+賳j��gNX��Ã#�0�`;��i!��&/�3�ݢ/ʢ���J�۽f���x�-7����� KwK��=�t��;0�<�⺟��f+�G2�c���/�I-���-oM��ִ���[o���ҥE�c���E�hcۨ��n�+c����ʸ`�0wb�ƗD:�/�y�8�QwL���֠��:�_`;e���x_:�o�d���� �Scq���n�(��>|�/
;���<���ɕ}����'''�駏4��L��)�����0�a���������b�]wXE���4�u�Dޭ�oR�%i{�����V0o��V��e{n������]��xD�{����=��{l瀀P�Ǌ f��ܷG@7l�ɩ��;핯z�n��t�(��gO���?w��ו����s'�s $� c��,YU*�*�j�۶ܶ{x�{ؒ�;��q�������1n�֕eu[n�,��X�E�@������������ �J��]{�{���ߜs�R�*�r��t�'�WȒ-��͈�!Mdi/_����6�Q�t�э0ڈ[�dpۭC}��b���p�@�d�T�@|�{� ��'3�����&����ϰ��idg�183g�bã�dq&�r���a��z�`O O#�8"#�1� C/��"hӲ����?�}�c'O���`q}]
�.����K�
��0~�羁�gN$z��Y��qsu�wQm���L��i��F�(��v	��N�`�&ҡ.&�|�����j�G�o��l� W���&��u���˜����^v���s�d%��w�1zѷ���!<Pa:����G�{�ʪYZ�7W� �Y ��Tm}�-t����S� iM�ոh�� ��/l�f��obb�4{�o?r�5�A��-j�Zá�Q}g�-*�eFeѽ��x�����ӭ�B�y��Z����	�4�����D_�����}��>�=Y��?�O��<��ԟ�=y�x���W�4!���������'Ʊ��I�5��9�F���N$՟��$ӶX�� J����v��;�"vH�E2L�L��k�6E�6������o��%���}�v��DZ�ڌ�PE����U��-�o����ԈAͽ`(i���]�L�Af�j�0�|�fz�a���	�i��� Im.>:���BԺܣ�N!3���Èd�Ћ$1I�O��H��{i�j�U�v��@fl�f=uE
��r4)XV
�P�Z}A~s��)<��sX���V�������5�UC�u
rE�H��%��VC�Ї�����p�0��@s�����`ƺ�:]�V6���m0\K�Mo4�	D���́�(ݱL_c�oO;�P]+��w�q��?��\�c���LXW��0��|�iE4�ˡD-^`�-�<�wh��^�)��_ �	�5s�ڸ�2�0����`v͜Q<#��_�|ׯ_��?^����\��J�V�J��]΍S����jA���E[q��}zj�Z;��?9vv���Ƈ��\?���,�O�"��O<�(?�4O�{he�g�*�{^u���7?�����a��߹�ƞ�д��Ǐa|v� T@vf
��A����J��ٹy<����O���X/����%,k_j�e�2J�y���}��'�w�%�7��׾�e������,j�-�\�dS�4W[�Nu�ڪ;���Ҩ��r�rh�1��^�V,@o�4�&�L�3U{6&�k� Y�|v�����g�i�L#�F,;�����zth�@?�5� �C(����B�߶)8nolb��b��3��S����%145O� �7޿���;��0��8ꈱ<A�)_� O-T{���y���,,�af$�dH]f>���v��]u�[>lm`o�B`�K�i�A�'����nm-ot�f�����;�ɧi���� �������h�ũ��߈G4�P^��9i�{�6�E�'Z�P&m�^�봺�A�8 h��E��]�^Ҙ�U���ͦQ��߸a�~p�w3���0@׽�[uG�l+��x��y@��l�k�t�ӕ��x�8��1?7�X�p�)����ɜ����Aq>n��Ǭ�q/|h��B�~�+�a�������?�����q�W�oW�^��������?~,�y�-��LOmX�%u���k��~��[��أ?5wбc'���/"K`}g�� ίm�۷��E��J�I�m�l?�z(��.B�����T����?�;��3���Y�O�����{(S��1e*k�0!�'pk+���*�a�y-�b�pA0�&Ѥ��>|���u�M���^�e�J�C ��E��I�?C�?�`zuc^�-OR�
��H�]�?��K�^���T�lC/mУ��w�e��{���e)��_'�H�5�_��i��B���;@�u9v�$�I
�0��u-@)�b[h��˚����:�#8� �)`,�G�[C*��$/�dk;���W��{��5)�"h����1�����az����=��yx�~����Q<�9/>O!vޣ�!������6��ܠ�+��i�3J�M�"XJ��w���Ӏ�V�Z7��d�X^Z���i꤭���g��r�mڥ�@e���3�<�+�O(h�L��_9�U9@a4�I�ԉ�o�뿃ɉ�ǪW��}:^���םS�>�=)���-�?�i���>�C����^`�4�t���%ܵJ٦��D����R�
��?9=�3g���Ԭ�������b���U�њԞ�]I��v���uPG�Y��t�Pq�������ŕk(o��AM�Z)bue�4�Z�A�;O잱�Lj�ej���`9�b#3B`B���[����Ǩ�k�}��|�QEao��PQ}��1yt�,��[
�\�F��Ⱥ�6�.�N����O��~����LT�:Ԟ�@���n4Q#��w����E�R�
F�(�D�S%�7kUj���W	�`�T~�B�j[����ƑL���K0b�����I��2.]_�;\�5ZN[[�0�pte�G���;�K��4�{ �0�:p\�p�Z���O�o V���[�ѣc���J}�^~�&hZ��ge���N�{׆`��'ꚑWXy���H�
�eS(�H�Q�ƨ��(��)J_���1pW�k5�u2ϲ�2�$��?�x��S6��Y�?��y�X����ܟ�+�Ӆx�9>9�����gW��ᡔ�����6�L���V�5T5�ܫN�ٗ������pP,c��)��#������U\���j��=��UzuF~LC�aI{��������@��Fn�-���pt�@�J�>�a �+�abj�dܦ'����d6j�6m1D@%ڶ�D�D0���� �r{W/���[��Z][Ekm�VG�5��p� N�A�&��JCm"N�ߑ�G���ҵC�b��f��\�B��<Tx&2�� �����I�ǧ$��>@�D��X�u��gka��އb1�cI����Eh�Њ�*Vp砄�R��֋l�ZX�հ�o�N��(D�Ң��~�)��-`����pn^��T�t��	`ėƛ�EG�& ����	�%������^�C>�Ͼ�����{�59���n]D�}[��g:\Z�i�E������&�m3�������8^�Ěj��W���W�e�!�zk��dh�����'��)�%m>���#����45誅K����A���	�G:�W��ǹ:|�P�Z����������v�&�?�����h����:�pw���Aa��|���ɼ451�f�O�^o�N&юu51D�N�'�*��D�==>�n4���<>^Y�R��FR"pTL-i�}&w�n�PC��W �g:�J	�a?&2	���~'z/��b�#�s1�U���`lr'�:�25�|��&Sh����;mݖs�q5}r������Ct�\�%��;:4��Z�I�²E�4�)(�uٞ��
���V�Z5�AL���5�O��Hڢ&�_���
뫨��XyԢ�`,�]ZA���˄�_�DA�M�R��� ��
���È��L�����ӈ�M�a�0�[;E��W�Z�`�D�Chl��	t( �P��1
/�q[�y�6��D5�i����y�M���`��\���m��t�ɾ����0^�����w�?��U�r��%/����7�{N�G����}����0��(u������gv�%!�d�)9����'������6�Vu�he��r����`�q�+Ї����Y��𸛯�9���0�t��	��W������O��?5�{�1����{Rw~�8���u/���q^��b6�=_ӹ�dfRáo	ĩ���n���	��G1v�8�ol���.������M�$��*8ן���e�
���f�����ZO�M#`g���OS,033���:eomn��O�^k4��K/�导�͝*ul3�v�T�C�U�L!�\�������ds���ĩM��,��2�����j|�R[�z�o�Jxol�3X.�U��s��2�*@T<��2O�*�������Vӽ�EPx6X箝�ĊGx'X��s�H��"29��c��Ev�2GNb ;�Nb�H�O�����N�":9�of3���O��`��=�r��@+���7���ա�{M۔ud ��h���6���|��m���Z�+���S�)�����Y=�;{�zw��t���U��m��<�<����n��wڌK�t� +/j���2���]Y�Rt���u��R�>�^��&i�j�=�[(�haV���(���N!���~{m�F+���,ͥ������G:�����YN�>�����yu�Y�g6���1��Y�mU����*߅�B:� b���}|�b����:��_?�=G-����q�j������h�m��{/�ȳ��������J(v}�	
Z�/Fw�nE�7��U�)}i�:)I{���c�(RAj��Y*�ujAa��RC�Em���~��8�D{�<��!�GP'*�^ݤ�[�-���V��ZP=�g�G�Z&�S:i�d�5��fK��F>�Q#�©�u�h�I�oϽ�+\�pX����	mpJ��GD���6����B�X�r	슢Y�B�\%�L�c�������L-�-0�
��[�W,I�4D?��82�N�?4�f4B�}q��O-�����C���q�y�",*� �G�&0���@�Z��� ���b6Y+����~��]�\ˇT D

�[V�����ay�/�6������,i�;zů�" Ӽ����-!�va ]m'K�����{E'��)/� ����+-]�2R8�\�����"���U�Q��J0?`;jF�ۋ��� N�^}��n�٢�84Esxdǎ��G8�����sVrw�8�*��]��?����a-����t�Y�>�q��wal���H��܋����(����9���p���/4����>�y�_�X(فi��͛�����g����"A��bۇ�_�7��dV�����hy���G����Yvm��o��*<>�F*A*�����~�-����c�Ϊū�O4+�\kQ��`���&KA�F�Mƪ�}��,`5}���u��s�Z�2A�iL���G(���$	rj��^����y��i{��C�Y 7C�_B=Џ~xsz���U%2�j����]
��흮��6hU떟`4��&p�[�K�">�E|h�e�"0����n*�|�`�Z;5�2��^���m(�wL;28�rN E-2*�El|��~�H�9�x
�9 3�P:�0��f���kk�㵳�yW>Ս���Ue����PXЂt)�|[]x][�䴅����R^Y�w�$Z�2��k���2�Tu�8�̒�3�C/絃�g��q��/Ӭ>�7|J@6��^{]�4A>dyL��5���k�Ba彈V}��H
�fj����αcǠ��t��]��\N�>����'p��>���a����s���f����],���=��jX���^Q�-����=׷.U�����?O#���;���{ث��b��O;��7��[�<�7��&��8�Ǐ�v����zi�u2�4M1�=ׯ?��g�
���ڻ<�_	>�on D��$��_��q��5�����h�%Qc$<��<��|ys��(w�ȱ������6��:�����&����e����
X-""j�3�?���^�Bʾ��&�Gu������vyceset�y�h�9�~^cd�j�h�S�@�B��`ޤ��{��j��V}�P	�z$�b�zԈYu����A!@��غ_�V��wR�M�e��B��h� ㌍�X7��S�_@�B.=9���8����?�]�}H<�W�2Z��'ڛ\]F]
���-��~@5���Gm	��a��O����n�!�B��am���m a�)�޼j�<��9�vBVW�:������,��xڥ�{��h��-)����i�9���jV(����|��}�6�a����b�b��"hں��#G0<<�d�H^�?�ӷ���Wz�C�tj'/Jz���p�^A���L����]?��🥳:8��O��cR`kW��\ߊ$�sw�w�齸I���ڕ�ŧ<��&ޫQ�4k�Ѩ���z]˭�H$�8�"6w��מ��
��jg�f�����V�T:����ԝ�Ge�҇�9[�"�l�,#B *��ڴđl�i��S2�1�1�H#32A�3���=��l;���$�)�՛֥��;���Ɣ�N����I g�4��Щ��?M`j�Z�Dՙ�������^T��Y�~��g���X��Յ�gy	�|�P��S8�I	TH����� �� Wy'�H+�,<������� ɚt$��X�?�V�(������g�R�ku�Dmõ0AZ�z�˫���(���K8H��&�j$�
�)\Յe5���ݧ��!�g?4���'��f��� ��7:�&��zȏ����C�گf>9��� Z +��xH�~sW^z�N�ީ��k�R�Oo]+w
�%���1�o��>��{��ox넊���7L��٦�*͋�w
��-��s��Q�؆u��0v<�ӷ��^����)�����C�X��P`�{P���t��>/�?n䔳��=3`�{#T>���u�x��"ｈ���o#�yF�7w����?��-.��4 �W�@�R!�vl-T�́8��?|�?a G��2)l��[Z�'I ��}��X��y��;i��w^�_�>v�<�#�4�w��Fno]� ڮ��Ǐ����8n�nb�d��F���L�̚�\��6�K�#�	�hR[�Db�j�#�E��	[���c��,P�f`�;��o���7�;�K�,�
�	hy�?Y�n^�d^�:�;L���;@� ��@����&�4pR||gè��c#�3@���|�|��~Z��j��5`+`�x�:ֹ����n����6)Ho]����϶�Px�&$\hИ%�llb��lh_�\-҇��k�Vk@�4o����05�A��=44�6��G�@]>>�'2i۵�� B�v�y��4��o�y��1�u���G�F���_��\�n�&:T�[$�բs�~���/�Ԗ|���U�Xև����7�%��[�+�c���^�M:l1y	zR���������ɓH�R,�Z�~ǔ-Q���GE���+�=���xlu�%��	`�Uz�?\�pr
{�;6��.�ψ��������r�[��s"#ݻ7�o��w`������|�w˝��\�ۀ��������w[%�k`OZ����D�ȿ�����":3���
���M�,mk�HVG�i޺�vI��|�{}�|Ao]|��r��O�G�;���otv7ֱ��j۲�:}��|sk�
v�-��CC.��.���U��8�-�����dM�kJ4NP�d1}��=�<�3S�Ө���J[P;���� ]{�p���_w�^����3��[!��3W�\u�[1�7�D�w��M�] Ϗ�,,�l������qy5m�q�^]Jx�4�g���z4�!O�E�i��I~���Ǹ���?��ﾋ����kU,#L��4SIs�[�֮��w.]F���g��Z��lPP��"�e��&㈆��� `�3�|��i�Mbt~��`hvs{	�4�/no٢���0:	I��A
/u����B/`g��vF3*��K^妷�ҞX_8`}�E�K����z��ֽ�^ȼ��o�������N���grvQ8��;��D�^ϼ�!y�	��<u�s�s1���8ˉ�}l���x��鳝�_��o�ϒ�VQ��Cz�8���~?n&~�N9yt�?B��we�`�"P��dM)R�p�	�f/A�zw�b�D龗�����U�xc��JKV�Y3lO2��[%#{1��=���%l��#4=�r6�}"�Pz�@	�`e>�0R��@���������� �&�hp6�O}��n]�ŝM���Q*��_}�+k��/ �������Sf�ԩ�7�!���Sٙ'�v�֗��|(�E��{'C�LWc�5���m�,��ƪ��AWo��L�+����-����=�V_Kc �d�ˑc��*6HA"����0����~�	\�� F7;6J᤮.��w�L�;�Ժ~-E]�.�Ϥ�(,��f)�����o����j
u��^� ]3�yH'i�J� ���+�no#F�*ɶ
������c�i�e� �G�^������- �m����@xh:iK`e�lm�֬f�|�w�v$A�i�J�!����ˇ஽X<��{X:㷺`{t��f�t�x��Ԣy^�;����}a�թ�|�p���4w�㕺�gʛ�����W����^����򫩏�m�A��J׏�ɝK�a�S���������^
��*�9�|������\N�y�i��\�˫�Dt��ɹ=���"1E:ΚJ���I��4�iĒ��#����d�&ǩG�2!��y�����w�I�g�]��CN��L��!�՚�U�B�a���4�Cd�$M�ŕU�\�@'�D3C�a�w�0B���&�(3>��@��>�*b|�e�:p�Q��֠�`'�f�A�\���&��W��h����<r9�!�|p�Cܸy9��:I����	��|�QK�IK�Ԧd�zW�wPj�Pn�P�����pj	
���uúІ 2�M�*����!t9�V��󞓉.g�.���[ڤ��A�:Hi��^N4.`RZ|�CE�P�⸏�;���^���U��U����)�9Z	{�=���"Qf}��=�"�,WP��D��~��N����h��gpzfS�����Cl��L'��O����&H��K��	-�o�h54i=�Ẓ^-���7�as�?M�m�
���"�J+�ĭ��Qx�_^B@3i�,B��S��	b]y�-e���v�{�M �o���S�9��}�E��9��m���u��Kf��.�M=	kE�)4̖��'QX��Ց���<�Anss�g�ͭ-����Y�0+��3Z��o�<����?���c�����0�ܺ)M}Θ��+�c�[�Ś�pzY�W��MM6@9����M�T�R�A-b��CQ�(\?����	2�4Wcki�+�"C�]�Exn�
��OS�Cԑ_:'R}������%8N�ymjt�hS{@��Es?��v�;�Gy{��=l/��h1�vW�2^�%���9��6��J���E�]�����P�XE�V�_�zRc�ՙ���L��������	�2������0kg����,=g�v�6��hEm�BJ�4h�vП��ڄN�;�����9�
�D�[,�g>�6�j���|h5b�BK��-���bOK�T��Hڹ�N͆Ɍ�S>w�Kּ�����_ʧ����_g�6�}X��4u�K�x�u�U�b�^8�#'N��tVWW���-��F��_������R� ��0�`��l'�<ە�;�Q��tP*atj�ӓFW����z��w��tӶe�Ӳ��lF�C'��y�4��h]�]���ע9�&$oK�J��k/#�%��vkԛ�L���b-����C�M��"o;7��%���� �lΦ�2|��R �չ��3�ϖS:�1Yb�	9����ʬ+��W(5eX�V��r���^�Ǐ/�>�Z��@�o�'w����A����s�>�A18����sw��ܡoH���'t��>��?#G���~���^�."���Ե#���i�(B-=t��%�H��X��j��D;ڒi�Qڅi�:���y���v�d�ZM�^g۷m+TM62<�Mjs��'��'1~��	���M�+U������+�_����+�mo��;��zm�%�����nH����A{�ػy;���-t�9D�t��N{ɐ3�*i��N��0�ui�� +�
�"Ci��S �vW�u3]�V�������|F��$�"�G=�PO�/�S$�����uo����jQx1�&^Տ��+Pk֌՟u�(1�*����u��b���ah�b	$�ǾS�z�a��;{fo��\$�o������&_1<5�}X�k{Y��1�N��A��F�)�0��M�_�2��o�����*�4�%��i�4{�O�S�(4*���z��wP�5fs���E��êV�f���\�` ���2�����������U<��9�:y�@���#�?:��Q;NP�i��m�˫�K[PW�SI��N��k�k[�ͺlJ����0�Y3�h'Ӡ鋁X�D���O�N ����'l��^v�����ϫ(&D�!�0�P����t���~��=d��54f�v�;8~��v8�k�O�={,�����s�>��1|����G�1���*8���_�+.�^���ݚ�~;/�B�ܦ���x]�>]I d �A\}���̩)Wx| )ҩ@�!I��mN���n�1#���&�m_�L_{�����9�I�	��������A��	T�x�긶��^��6��@f�i�3>���k�k�)�����j6I� a:��G�C��MSj�C��,��P
	�m�%�_Z�B�!MV ��v76P&�ϟ>m��bdӾ��T��X��#�_W��&$�2��"��u�����Y-1,��4x�wC'@�z�>w^��N��H��Ǯq���O�亲L�S�i�|H@�şAjd��e�YEr�3mr}ǫ�W	�~�Tg�T�\����m�Y�f�u�����Ν�AT��!UF�t1�v��_�2N�õ+p�qh��"��-�J�c��>3lo��Ӛ$��I:M�z���M�V>z�J�:C|����W��W_}�#�$�&Ʊ�p����9<��s8��}��Wp����7��z�R��I����[�>���-^]q:�6H����0��{��3Cv���!�� ;=k{���Y�A�ϫR��x݀��RY��
Ї#Q�KҺ/�����C�4p���U,Lஙg�G�Mk�^3����ܓ;#w{����ƥ�������Oі��t?{�]���_��$��E�b$��dC�EO�s�ui�Do�O���y��ɉ������]gC��Eu�)�R�d��\���#�k� �)�g�"��i�놩�Gc�'���w����{�z�Y�m�8�N�5�������+��ܺ���&r�$�љj�![��F�oׯ\�Ε��Ϻ����YIähb��ؤײmu	�l�kZ2o�c��n�Z=*s���]GL�Y�P5	"m�	D�{�����U�ʯ@P-��]�c�O4��s��������^��ON�u*}��p�����iU���Lg��jJc"�����Ց��+���?:�w���;��b�]��/���� ֩�B�M����1�����׿��_zj�:�X�������N�0;��5�;˷pt~� �6���M�l��f&'p�Z���0��A���Wz0���q4����$�E��RY�}��LR�w��@):�Kc2AZ��љL���,��t��"vHg,� ����D�0���pf�2�D�fljlb�(���I̞=����"M@OL�`��I���+H��c��q��<M�?CK�$F�#42�"��CS��kM�/��o���'���)�� ]��:�I�
��m�������@���}�����O����?��'u9vu-�����_4�3YE����ݻߎ�y�����BS�OB�lۂV*��"j�@]�QK��)�e�j7��W5ji��ãipT�HL��Z�q�?���i�5d�a�mm���^rc�N�C�U'	?4�;{���i��Tۘg�G /ǰ>j.��|H��(5~���K���&ض�4��u#��P����	�a^4_Z։���d���S�5ԽDFnR+KR�"����,_��jב ���
.ͺ�ba�3iOǪ�0裬i6���������#:\��k���oi�
5um�r���4s\�l�O��*i�b��i����RԲ{�6���4�[B�K��^]x՛������d�(h_��<�<��<m+o����;L���NM4�33c�S��詩�2�,5�.ifth���L�1?;��f��U����ְK�JeR8�p�.^���#"�-���˯~gϞ� ����C�,6̻��:p��k׮��?���z��U,�ܡ����bT��i�!j�x]�{ll�e�Drb
��L��>�4��'h	L��3s��'�� �p�1;)�6Nc��&����ƆG�H�v���#Oee��z<G�<V���IN�z�,L]Uu!i.�������k7Uk?׌�N��>%����c��}�'�v�~z���v��[�yOc����{��Y��9�J"/\wޟw�~^!#�I�j�za��lX��j*�9�xߴ�N��A�Z���i�4u��Q	g���r�~���	�Ӂ����(�n4�}@�f ��@�$�i��j��o��;>��$fM�&���c����}{��ϐ�ni1�Axjc-'W^��󥙿�x��f��P�8@�� [�P$2�a�z�,��� ����ZD��/d�Ng&f�AӬW�Ԥ;( ��ؾ~��2Jw�QX#Phh"�/u{ҡ��%D������������쉅�?�7�3
�)�$�W�;�VW��@ϴ H}��w6{�"���z���DX���ۍ!X�\89�s�7�����[ػ���G���;���g0N`���R���R�6��ִ�j�z��sgN"F�+�ّ�DS��m�}�5�y,--��k���f^�8q�4"�$��7��ǰi��e��G�������hǏ��D�T
$��'�4�e�ƍvv��J!q������x�wq{q�@)bg�TZM��潣��Q��$fO?�)j��G�a��)NL"�x�̓�;�Rc�7]Z*]�u��d'�fuԢ�i1,ZQY�������3�(2q�$��!Xq{�����Vk��:�X(bow_�ʫ,��uw���c������ܑ�;%� /�የ�ɜ��~�PW�\?݇��1ѡ���6�q�U�{��W\.�jF��C^�	�ۅ�
�]����`�F���V06��ڧ�.!ѩ�CN�^(�,���dֻ�xں{߫?O}��΁�f�S�j�:��Z���2�vw�����⍛$~��sG���i�f��)�V�����*���[�(�E氁��,<�b�c�?��Y���\V���YG�Q���Տ�q��F��9�?�%c}�DI�b�-���M_'��Q��S;c�[�����S��]ܾ��?�#����Z=��F09��-B4��23�Һ-��.ab1���m�9�7{���u�����u�?�,�+�<̆l��[6g]ϵ�׾3���1��xUF� ׮�a����vՁ�]�1�%���^��!W�~��x�4����cOhv���^Z������C1��!C��6D ��gݷ���E80`���4�*�_~�;���H��5 ;u���$�l�@-5Ƹ�(n_������qk�L*����c~��Ашf�H��R|��s{i?���7����-lm����Z��6!�@詻%��.9V��Ob��sx�կ��Q�=17�	*��U��=i�S���͐a�i���mY,��{����מ8�N��"ȏ��P��a��uw��^?�pm�۬wi���Z.��g����-�A�oע,�[�s���
�!r�s�� �~�g������,���N%�Ʈq�[b��лR��=�\�D������s}*@���l��[�L�!�I9��S(hv A�ڪ A�QY���ݖƦACi�>;��X> ��4�":Z�����4ş���;�Z��Gʹ��Y4�:�u�@+W8@C{�P$��bvڔ+:2n{�k1``�#�oܺ�v9G�������i M��Y@-��� b��5Lּ�};At��f��r�I��yҦf�}�cl�>��Qؼ6�Q,����*��jo�DM'ԴL�QS5Uod5#�����s�^�yV�+�N�1��"dt��9�))��+ƚ��r��o	@�?���B�h_�X�U߽�v/#���x�<�}m�i��dj>�_}Ӳ���� 0I��>�Kf�y	�;��ٴ�h���o���?<o���;6�qxr�T
��b7��M�V7N�`�=u��G�`������"�@���G����  ��IDAT��)����������Ǘ.�ڍ[(Ut.l�tGE�ͩc�-�ۗ�É׿��������P���R�jҞ3Z�Kw�{{;���8k�Դ+:8��Iv�����S��E��4ōl��R��Ј1���+x��N��2��Q�I����~���.�W^~3Q֧�[Uۋ��P�/�ܟ�9�8� @�܃����=ح`�3R����O��,ew���l4i�di��;�k�N��۲j���9��i I��YBaߥ�"*������Nsz�tT�o��đ>�P� R�R#o4J|��E��'b�L�꣏?���2J5"��M����=�:�۬JR]<����IS�{�9$Ʀ12{��	�l-�釕�b;+KԪs��hJ����5�O`��b:|���+�^}�e�|d���1�5fҠ]D���]����r� �ajX����#��z#Զf�Y�h�� ����.���s�~����;�w�����5�&���V�8I��<
�%���_�pIj�lƦs
@w�xxi�ҵz�6��T~��5mG��-}�;��¦��^v�+`O��a��Ѫ{n�y����1L�������o~�����jG�1푩t4F�K�+�u ��[o"��?�<ub�V�j
��ا&'iAV�M�����<��6����~���0���Q��(�I��.-�z�R�s��c��/��˯ 57�Z8�=2�69�,�.�������_����g���?�ʕk�y{�##�,���T7�O�%��{�ި\��&�������g2XYZ�5�Gjd��H3�4s��ĸ������	�k�'�Ty����K�]�~��?�3����s������ӑ{(������r�<�D��<K[�.MeQ���Zf�4MO�hɴ�M�:��+m�t�y?A?`S�$ݭO��7�����;͟�D| ���r�Y$bxj�M�U'ȴ���­[א�$�H�l��Ǘ.���*�hv����U�!��3R���)�(�m||�
zɱIL
���:�8��}։4be2�rFhU�hR�Ky�����\�ߵg��A`1뢥�'-��3?�ҭB�Y�2��`�&w7�A���zI�}������S�	�4`̋�0'��L��A�A2����k��"C����w�x��w��~9-N��L��{9��Us�5Cb���K+�G�ԴG�c}���$�EJ����3�N#;2Lr	�>X{J�%�2�o��!��՘��'�t���V�r�_��ī���W���Q�:Ij@���q��r[��%�A�PÃc6XߨS8���XGO���/|i���},�`hf�f�D��?�����ѣx��l�ԋ/�h��:~nhh����]�r���M�P�����rZ;�Svr�%�=��{ǿ�
�N=� �4Ǌ�2u1	�{���+������;?n����<�VH�1
� �Y�U��kՙ.դ���Y��G�G�deQ��
L����;��v"�� �l�yG�ſ���f��BѸ��vu=ɋG$<]8����~~^g8��܃��톑�2���w
�8���8勞�3�N����s׏��.��BM� �n��Ҁ�P]�<1�Z��������z<���po|�����Ȳ`�������}��I�����e���s�9���˗�����������j]��W��V����j�qX��)[Ĕ�:���(�$�?
d|�L�i�N�,ؠ���@bp��3c�(#L�%��Z�-푴%o�'�l��ڰ+�JcD��AۓF�@�9�:�M���H(�;�1/-�wG�IC�T�{�F��RCYM�>y���i�߫>����T�}&�ƅ��?�ӭ޷�:��f����OZ��2�ȋN�K�O�bWƉ���w����O$ x1�c�wm��0�8�w1	Q�@�Y�Rʟ��I��P�Ci�:�Ĭ-k;��wGq���>��7/-ci��S_�:~�7�{|����3_���3Z��k���)p�_X@��t#ALL�Ѻ��Ƶk(�J�a����py�fԨ� _��n,.��E��7r���<fG��_���/�׿����"}�$c�v���ljJ�M�º�r����.��E�S0=��H��;+�n/u4���:&�K�`<u�I� 9�h[c;e�q�ā&1���z�5,���G���_�O*�EfpSS�v��C��ԅB�Bei�-�ؤ~��>甛��H�&U�����=�[�C��O�7�{Na	�=���O����E]0a*�Z�H�V��uzz6:AJ"��ʥ����H^N�,`;�\����(�����0]���	�M[�T4�*`iak�\�wi�R�ÃH&�F���T`�H�d|5A��;@�ڵ�Q�m G�ۄ|С�P��� �'P%HWY�:�X3@�b�4('K}��f�����y��1}�!
����Ri�~� �B_Օ O�!�S��}G{۰n5&J�|��o<�b}i����d������eȸ���=剒��vb~c��6Pg;��R%h� j�ၻ���Ѥ���?�,6�YXź%�B���D��ɴ"�����-w�\`�h���Dz�bQl�
׿�ZwO�����x���N	>J2���.�"�l�|�ZB�Ă�������',�U��025���$������n�Ze ���ǎ�:<���U���
.��"l��/��jЏ�k��n�:r�}ܸ~���65R[-hf���.�Z������яߴ���y�cӳ��[�Z}v�
��,��;}�Ͼ�(-��D0��&���u4�LSgH����SI1�֔K����*-\+um�W�����v�8���i����$ݵ�ۭ@��� �x��_ŋ��O8�4��>K#q���0I�����,lMyt;Yl0ճ���j{���KqⒻ�S������.�\gBB�֫NK�����v�����*$�i4�A64_�˄6~�50#f{3_�˙T�K͐�A:�]%��p�B�ڑ!�y��f�@�i�U�f���\�f����bgD�z���l��9�bZ~cjVm
�N0�v0j �d�t���h�� �M@_!�ij�N��?���O�AҜ�2���!FQڶ63�6S�	��tZ4�sG�K��#i��^g��,���e�ŗ��c���N�O�|�i$����8�^4n�	B����6�;�ڑu�y���=c�щ�-1���)e-�H��A�i�d�#�f۩�I�$� 󞤙>@uں��T�]�~�{N�������-
��do`���~x��W���yl_���=�	�Q
����|
�B�[ܩ��ʻ��F�Hb�s��\�U����s�&~����[�_ƻ��t��Ň�<y��複������&�gglk���kW�n5�*�=_n߾���~������yk��@�\A�R�q�۪��&�f0{�Y�ڜ�Nzj�5_k-�D��5���i���La1뇄/�k��� 62L��@U��nn��퉵�=/>֎9�B�JG��>��رSB3ثR�R8&�C�7�:�B@)T##�v��hI�S����ޏE��=Z��3+R��9��7��? ]�P�%�>Up�3O���9�V���\CQ���3�ػ:m�y-��F]",��CT�_�4hjO�Pؕ�e������[�Ͽ4��i��[4*��χ�v�m2��`��4�ї��;(��qp�cDڂ6_�y�7o��52�EB�׊Hm����x~~�ڍ�Yc*�4:��C�v]KG2d��1�`<�O��:N[�K�i�7��H�U�&3.!�y�]���%��Y���@`dc���ї^2��&Ү/��l��Y{P�g�#8��hL����'N��G��;�_{�4�6c�}�8t��-��3z�;ԍn���m̫4��i���R�`���Q�� �+�O�3��ِ�z�	��@]^�].M�柲aj�X3�4nj5�V��y;W������ڵ+���ư�T2oԩR�L$ⶶ!ݫ�YVEm�I�	d���hn����"��UYH����c���j/����+���L:��Gg1�L�;��3���,]m9 ��y�6�=�����o�G�������	
~ C�`��S���!�4ۤ�:�B��Ҏ$X#,-$zR*t�G�̱���5*$He��d��I���*N��"2S�vV�E%d��E��-���ܵ�w'�_LO�H��T2���֗n�U����9L�Y�������Wס"Tu��u�Ri;�r�0F��,��۳���*��g�o�������[���񨸔)���tV�~�'�N�p���+o�:���s�ɫ���, P�I�:�]@/��Nr�GV��L0�����b@~��w��k�^'6���L ���t�ќV����j���Z]��5XZ.�H���H�x����p�#���7Q(X՜$�2ԃ6Y�<{��RG?��4�]��,=Ӹ�Ly�ӆ��յis�Y���A$(Ͳ�&��ɘ�s� ��Ҙ��Grp�1�8����42Բ��=�&A�b^�!��Ɉ�?2�P��,��em^sz�(�?��@���Ijvt-h�7jo֟�]�뵨����b����w�Fq��gm#mt{{m�����h�I�� C����Md��Р͈��.p9|H��+n/Y9a֩�mMQ����!�/]�ҷ�||�Z��Q@���)�%
���B�,:�/Џ�6b��U��R�"�0�>BM�[*�U�۔��fД?�O�G1|d���Y��`�VW��Gmg����K�`���v{K6��>���<Mڢ�k�mϕѱq\�~_�d����4_<���#�����=��Ͼ :K�e���H��CMDP;H)#5@#'�p�Ԋ�v�JNN"<=����*N�%�S)t"TNX�6�_�֞�W�nm�o�)mM!�E^��ڲv���d}n-�D7w����pdzҴ�>B8kI�߹)�T�6�{}'��~l�;F�p�����}q>����!`�="�G���3������<�ˋË�^�{Na�\ଫ�<��@c"��d*�n�/��.Pה2����l��7�+��+�����u���"fS�7�`Xf[l��O�������D@ڃ�Nm�V/��.�k$�6�8ҙn-��;���K�F�ʌ�¾g����6 /�&ha��j���x/pW��]�`�r��)t�fi��2s�ZF����1��.5,E�%h�jIwf�娖z��#F�R�z$�̄�"��,���8g9�8D��M"&\��-#�ŘO�Yf��=��T�V�31k�b��j��-�|ߩ�Yx}�Li�i)_@���;��k��Y'gB��.�d6m�1���<v@�ָ����{�/�H$Q
�	
�c�
W����c;'���(���VGqi	z#G($5��%�Pcd���W?�ۺ���k?��>x�~�}�ܸ��+�ug�����H���Y��nI�Ε���X ���3�2�wְt{��s����������NK����w���e�4\��I��"��)�Q�g�`�� B-�&�N�n��4;E�����U��)�����eU[؉T����-��3�1z�¬�6A]�Qm�+ի_�����@����b��6ͪVU B����(��]�!�xÍ���x��e�N��8X?�S9u��7iY�J�hLʁ���9G��v{�D���4�u��ˌI%���O��_���+��AkX�M�������$�b��8ɀbE�-@u@�@�����J�^���g��S[�qv���Z�8��@�JB�3H�qk���T�?��0Z����k�d�Ğ������I����W-+�:�Y)����V>O3�� ډ4�bˮ�,��)���y�d9��-%3� ���[ױ�t�7���ͫhW
��2�!Q0@F�GΤʢI���n2�f�؊@2��Z��#������&h��(`�d~��o��W����\�VZ�{��p�ι���M��w4j�0:m��}m̪��d&��u�7���O��R�\������u�~h�s�9W~j�� 
ʈ��(,�H�	�W�V��P��VD5����u�:��4�L�jʤ��u��e\{��8x�=�?� �z	�KP|�-l��웵
���(MT��t�G�Q$b������IcZ��-T~Ճ���~�����+�7�l����k4;h��|����/���O��ܵ�6��TU&�J�ߪ[���U(� ?���d��S�>NP'����"B��
�@D�A���x�D/���V5F����v�U���˛d�) GH�I?��!�����@G�/`zn�ƁDkʫ�O��U��Wy͎��a�Y�sמ3w�A��oF�fڬ��|f�֏�u����;����= o?�=����݃܃���z@z��nP�m�������p�*��yu�h_��ii�6���8�Q���Ԙ Num�<�NT*M[�`�X,h���A��8�xu����ű���k׮�Ns��m�?ͧ-�J�����%j��h��"\&fΕM��e��m�D '�P㥦.�h��W��8�iou��h���v7������w�	h�d��X��Ce�Q�|�J$���(z�
#M��؅���S9�e���ĈҺ]�	]���(=_�{>P����A��*�]g �
��=v?L��Q�K�P���r��Zu�F�:P� S_�����6��֬n��a�Kn[	�xa�++�$�.�V׻��a!��Ҵ7o�­�Ǵ;��w�P! �r԰����k_Clj��S5c+!��`;_V����7Q�~:X��_�kPC �$D�n����,B#�v̠��(3���
����ۯ������Vm���i�>u�t+~!�S�m��|��X 芇Z,x�uV!|�5��)$g��&87�nG���D5�H�KRՂ�>�ǲ�XyZ�)���Q�)�Q�Vl�X@��jTJhQ8u�ak�b��@�g��k	V�'-o�	��2N�t��-;����c��5
�:��ӫ"�F��b� �-�b�om!�<�6�v4��{-R�#o��&=HY�!"n@�Y��[9���ߞ{гG:�X?쒰��ݓ��I�����{�ɘ>΁�����"t������T��|'��3	 5��Q�Zd�+F�?��:y�EuU�lOÂ2yJ���#C��p(�ݽ
M��,��2�1�Ny�v�>15J�nPsм�A#إ��Gm���-)�r�r�B"�ف>ue�b6���������xu�8l@��B��@��~m�������+8=I����Ԅ����'��jАq4Y���Y�q��������J �U��k�O�%M�˙G�*��u�Д� ޵V?,�v�����+}��	�V��h>75Ɓ��*�1' �]��`{�;F�@���.7VᄑELg��5�|J�k#N�I�����a�`����5�B�e��72�~�xꕯ��)�ZAl'ъ� lБ�k�o�X[G�B9�4hS55珴@(D�����E�y�0�hR� �X^��G������M�m���T N�8�ٙY��9-��@���:6�w�]g�KdP�Q�I���/":1���Jm��|��O��?�������MS@5S(L�RWU�����q�X��]��V�v�:5�0���ȳBX�N#��lT �[�zJV	��U
���\~�{���ظu����N�c��d����f#|�$OJ���7������u��P���k���p��+���<�o���>�S<���x]��a�i���8K�I\?��~w���a��1��D`�Y�>�5�KF%���d�8S�4�0�_��s�ʢ��j@i012��9��k��u�4�,�e�51��bl��*���u��%" �-����������%�=6�R倄�y�;���m�S%(�"�S�)��}�c>T6�l�ր�����"	lNҌ�5[�Ű���t*�v�����������7��"��=�\��LT�����������L��,א�0a����7��S���emƫ��>Df /�k��X�Dqi���np���r*��g��^�K�"��9����OA�`5���&x��;[�N[����R=���ri���'�7P��{�׵���\�I�H���Y,�ݭMV	H����g<}�|���A�ImӔ�	E?����D����W�]YD�iu��X�F��;�}�Zx]�ff2.-�{���Y_�>���A��֏��o��瞷mJ咳���s{g��DK��D����O�>yڴ�n2E��Ĳi�g�܁�թ=q�렖J��n��8ij��w���G��n�`��e�6����5������#`Yg�:��m��Z���תב�R�g���;���{h�w��}��h�(�7��1H�8�/�*e��<�m�0i�����Ix٦W���qc�+��/�����O�ֽ4���;�DN��%�~����>*և���+C*�*�
~/{w��}������P���ΫcmB�ߎ�Sj�xq��������@3ļa-��Z�6�=c��x��XgX�Ϩ}ˇ2aS[W*y;�M�T�ĢK$bah;ݕ�eKy�"�mFL(���A*bk��׎v�3"Q��U��:B2�?�i���tFM�ҙ������b.�1�̴垿�pi�*�4���^�7_}�W/ჷ��ji�E&���u��,��6��|e����*2���xSG5x��I�$&�I�:b/Jm)�d��V��f�ϛf:ǌ�C�Q3�`��be�+��5����ݫd*���)��$2��]Ҟ)�����n��ǋ�]�+Gq��:�w|j0k]1��-c�&1�ie�u��u.t|��k�1O�|�>Yj����cr
�s��ī�!;��)�Xw5�KZ����Pc<�.�%�h�����x�DH-��X@u�c���W���ѣhR��ɟ }$������3x���w?���fp��I�I7Z'z�̘��u�C�\�ض9��^ ˅2^�2N��*���v$vo�:��L.��4=U5Ĭ��a):'@{��z�]��ɏ���y���%?��O$c��#�z���d{�VW�	��,k�JC���5Y�/عv���@�:�H�J�*��ڞ�KAؠE|��ID�)����6���4}TV�,8��kľ�	)Ҩ3�V�ˉ�ڣ^��5>�� ��a�2�M�O���=C�C���݈�P����}`�r����_�e�b?�ßt�-�'3;��i��t�Z���m{^d�����m����>��*BԴ�껦�H�Ef^����>��}��&�)7L��VZ�fm)B:wt�ff����Y�6�=F-B��|��y;=}� �*5�d*i�*m�6�Rn�.��jђ��n6�i ���tz�f�"xu�w�NS��I[�m�w��ʙ�Љ����!�[&l:�K'��i��)���f�$�4k�(�h��	�d�V ��#Ԥ���4�����w�2|\��et7z��UwJxa~I
���A>lX��s�i�w���jb��G��*�Չ������H����@F,V�Ԍ�f��m�?.[m�y?��$�V��n��lci�I^,�~��_�W9�����la�e+U�s&�N"�8�ff1qlQ�k�
�^�3:mA�0R�i�[:�2� �SG'Vd��I�S� �y��1Hm�?6���<���& E-��b��y�&���;[x�/R��	a~��Y���i�˫k�>(�ܥ���J :q
щ)��OmZ��n+RY�~�ܭ���@�4�e{�QKo�`齷0���a�{�Џ%��+�
@��5�h����oĺ3;�U	]�)@�F�t&�|�������FELjq֓�AP��2C8�쳈�F��G�6��M1���0�S��'�b^x�16�{Ԕ()�Z!.�]��Z�j����=��J�ƭ'q./��.ǟv<����XDu*�~�˩����Gš�λ)w2ɐ�>���|�������% J��y�Ġo�cw'��u4%K�p
AC�f�N3N'H�5^O%�{�Z*F��hD�ƍ��v119LF��*�QP�� �����#�Pb�8	�DA��Zaj$�Ы��-��� �$b��˄��[iꣵ��if� SG����{Ԋ��%��������g1;G��C?�F��b�6ɚ�����Fi�7�{w����{�4��85ʈ��E;�Ӂm
���5o^Bwc	�[��S���ï�ܗl����Y6�dڴR1�Mec�Ҟͱ�3��u������S=���ڱh���[Ю�5�+�hiY��R��^5e�8���տ�=⩃Yw�KG���>�w._����k6��M4�;����hRk�2O=҅Iu��8��:��"��9���|5�'�.�����>��i��'1q�N}�˘x���-�}H1=�|����\W>�c�/�9�����Ƨ����L�)�?��~�o��]�6�&y"84���#6>�*�C@4@��u7��^|��Έ�,��wO���J����q� ������8�����`u��UF�V��'�Π֡�W�Wk*I��ƕ���R�(�Ի�ڭ{K���iӢ!]R:#��s8��ˤوM����4���ݖ)<��J�S��bm.|P��ƶgè{F}�aZ��E<���)�4�6ˮ���ͽ���g����?�Ze�A� ^,��IX&]ٸNc'a�1�]S�B�oڣ�x�\v;a�W���<I&�Eܶ��֕-8�cR�djU~� X�Bj�T67�	m�ۼ�(�!Dd�E�/�[o��qw1:�!@V04�fp��;fLS�O��h�V�K�h����PDr��t��,��Qjd2��)~��d�	�I�=2T�b�Jӓ#̛UjV: x�`%#�+i����򫯢N�^�uƮ��z��~�ͬ;a˺z��8��.Z+W��YFk�"�|��_�׿�EL"�S���>�d�P���6�b	
��S���/Շ{�_lw��~N����8�F�j����$���+���όP����V[��#g3���Ҧ�����%':��4�d��-#!��=sB@�h�N��!>�"2u_�5Ƹ���N�g;�"�$�H㜘$�N�OͿ��Ӧ[U��d:��iƷ}�*¥����8>1���5�E�����e*�ˈ��O�y�N��1�BUS��?K �����c���оDZ%�V�
�ThYF�YŤE1_�KIG4������l��������r+�1@���:�Z^Dq{��o����a�US��76Ц��AZ᪮�h,I�'�V����2���Y����5^��_E4���K�qO��H�b���		Lvֹ�f�I�95�M(�S���z�51����U�zџ�J����]�~�]�ltGZ9�����A�a��R|g��pʀ�V�c:Ϲ�ż�
�/-{o��޺ax�	k ���{�˕�c�F�5��ٷ0?�)��#�,"$�A]Z�b�M��{G����:���B�AP���>��p��ܺu�_a�4}J��4�D����b�Q*_�rZԚ�R�$)]V�K_��F����F4���2Ԓ���_��^n�j�F�:�.���ډ C=��ڣz���,��7o��Ң������/����ydXbt5��}�W�fe4aڥ"zd��ꔹR]��5�^T��.&���7�a��Dz�ª;H&�869��5��ݸ ���V��/���WWv�I`����ы��L+����
#�ݫCO@ʢ��ɜ�i�ѝ���|��j�~���WE��W2�;T4�f���Ob���iS��w�u9E #A޶#S�C�aj�C�T�����J���r9��~�mYd�7Y.`LZUg|����
~��W�³g��]\�v�j#�#6�_�p��3�&S8:7gZK+���C�`����Yה�{�Bueioym����k�g!{�����cA��V,`��%j�T�V��G��y��/"N��^�c,�Ĺ����O�o��/��7?���P3�Ҳ+�S�1�%}��z��Q��|���p��8{���Λ��o�+���&ݪ�KJ]�BTJ�hBڵ)m9�w�Ԧ�}P��?y�*����A����5���%���4l]���Ѥу?����5v9T�=��<�����y�X��(]8U8)��c�5 Jb��R�w�Q������ձ�D��4��L��>@*6�/Ơ�R\�u��SڻV��p�'c�G(��2)��/V�z�������s�0d�CB�٩���ׯ���ߧp�3N��4h& r&��A����Q&:�Ӂ��p�j�`���tL^�\D��LM5��?�eVZ�^)��$�$0���i<�_��bHD���������&ppPD��Xj�:�
��$uBjov ��Si@��ˋװ�����IM���i�W�9��7���h�s�&�&n�ѡFX� l�Q�,���Vy�V;��=�v���_o�2��N�/��������������7��iȩ���uڐ�/�s�1f��?�ӽ�?�$4$��S�ܤ!j�ɔeA]��m�����'ČE蓌v�2�C]݃[[��b��/M�Q���������+���'Q��dYû{Hիx��ij��Q��o�ɷl��~�V&)�R	������k�nYwQ'C�����d�fm�TG̩�>�ߣ`�4�AK[I����_�Lk�G�]G�iU��o^��������{�/��E����G?����?�o3�}*�T/���?��k�ȑ?bã�6)�H��y��Jd1�p��Y��p3TJ�Ϝ�	*&!i�̏��ho$rb�Ӥ��G�5Y�jkUk'��/���Nq��į����ܺ��lSy��*�MZ���q;~��)���G���y����0����[w��pA���"SF��ͣ��|X%ލ_Ͻwʯ��6� �EI:ZK�-���f�8�!�'i��Ԗ Z*���,��F����b>2�}m��l��5��VU�I����ɺn�.�]���{���_8���1
�i��W�`ee��X-��d2�iE�7���2B�����z�p���hfv��i�(-��0C�P�,�F��Va���È�[�����w?��_���t(����:
D��S��.��������Ǻ�:��@a�:�"����(�ۿ�?`�W��v��*��V��
�Bf-SlQ@YwK��r3�������%�'��߈Q�#Y [�P)��k�G!�xծN�f|.K�fJ���\��@��&`7�Z�?���֣]���JO�Y�_$sG�4�8��^�/��O�v��$��`~ST&z���(��|KK�_^B��
����|�u�q�&iD�>��ă,k�䠺�"�naT݋k�ݺ	_�����\<��?ƫ�|'O7z�X�������.*�677�/�QaQ��Bχ������P]D�_�ZY����W�\���X�~�+��TH|T�ȓ����86��K'��YȡD-�&��&��������'��K���]�@K�����	�&&mQWQw�Nq��N��n�Uj��͌�aza����ؑ���5�Z�š�k�f�H���ɪ�^�fmi��'ײr��7�o{�{á�����u'��͆��� ��-u�J��@^�J��.;�,}����?�1����=�}�{�7��)۬@�R,�F�4&�h��6�r�M��I-������2��:T��D��vi�bgi�Z� ���ө=�c%���	��K�V\b ;���~��^�3ϝE4�խ~�ie��W��Tɤ�C�����(H�dS��U
�/@WW���Csj|-"β\�U�KMM�k��{� Oc�Q
� ��HK�G$y�s4�i�/)OE�e���`�����Y;d�͏>Ƈ7���C��r�2���dz��j�Zu4���hj��X���ƹ������{��7޻��@��0����W߫�%��(�Ϗ��Ė�.ֽ�Hx�zQ=��0����jgiOb�2�Z.��l����35��տ��I�c#iRL�g�������
��?k����h�ߨ+%�`����Gc��X$`5�ڔ S�S�����Bi��o��r����(�mӰ�U������x�f���@�Z�e�2��;�D�o�ĵ������/�č��R��k���P��Y�A5�H@�չ����ʵ�(��yzb
ىi{���V͍M��� w��Q�r	�kW@Ɂ�hK2�m����,#���v�oٔ�<MZ�R���=�/��2.3����w�V&�T%	��ǰ���,����V{���H�:��R��N���>+TD�E�/�AU�c�5F��&�G�M�v;�=�ڼ߸w��:���8 �U^�Z�R"5�YX��ጔ8��nJ�Խ���ֿz��ד8�g��2�"=����Y�>Q��p�D�?�9��|��4v�!��9Dm�1_���P�ꦑ�m��u-�g��M���2�Ĥ�GO+@[��6�XU�0N��.	_r����T��+d��+X���olۀ�	2���	�/_Ɲ�;�����Y%�������t�Q=ze�֩��<���Edr2s�Ps��6��+A���ɦ0��̓]Th���'w�̜��
֥2� ��9�����w/_E��Z�4���q^�v�����|�ڙL`dj
�Nk�:�s�.o��X����ze~�y1ae����k�]�ly����!����n���HZ{*�"x�q@`՜g-�R����&��e���T"��H*a�"�Ȑ�S�f�(?�VV�נ���3VK`+�W����w��
�/]���+�^��65�D"�����
A����Uj���E4Hͽ]�>M��֫]yzZL���K��]�����x
-�U��m!B��]�t	�Ԣߥ�Ԥ@���į��_B2N�U�QK��~��T
��J��+�696a��׉C��х�s�Uik���;�����\��P��_A�h;���8�''l�,�"W��}K�ZҔ���-��S��G������{�c�����K�����-4#I$�L��I��6Y�~�k�z��.A͌Q�R��-ƺ���(�G6�v{�Њ������՞�wwjgko��v���v���3�ܽ�L� 7�w�RySJ�κcV��ͅ��E�1�Ro�q�XP�?��7�b(OJx��ןd}A�����g޽��Bz~8�'ɴ���R���=��إ�K[S�^Zv�����
 ��Q�G`'��2�� Ja���̥F�[���w�%-�mG���L١��l�٠!�O���|�w�}G��#�I��$�<���;�6�6�҉0̊��� �K��ϸ�4�)Ӽ�S��H˾���i�$ �Ҵj���ETh�w�욆�ԩ�̳K)�,�M�;j���ؘ�������k��g�=����s��Ҷ_H��#`�#�2Ap���0M������SPdf�{�c�2�"UX��#�`{ȰL����m����� c���
���?_S�$�4xk���h����B��.�9i���5�S��Z��:6󙍩sMc�����]w�aѓ�٥ѯv]m~;�f���'��FL����_�y�Ct���w�2��������(!JEA�Ts�+�F�*{;譮ڊI�z��D2��lC� F�q$�~�5ߛ�ޤ�(��.�[?K���r�L1�+F Y&����j�t�n��Ͽ���ƒ�y����x���_��'�I�,;�\��5�S��<ZMq�3M㌓f/��_0��;�>��$��^��UO>sc��K��7Y���ۋX�u�����y<���ɟ�)~������<ikdb��Y�Y\��C-�@x|M�%��0uè�OkR�C�\��D-ҷ���b��]u�n�{���]����bE�<���s.���{�r�����)h���>�J�ޤ/-^ϴ�]����1��_����9/ħ4���~�V�q������?v�s��4Υ���P|jDi��^Q2"�wa{ð��,��J�Ё�����.0`�y $�^`��������z�I�Z��sNB�Z�agk�vk\\��F���N؞*����8��y<��S��9",G����,��*��P�NF��Z�U{�֯~z5)0g�����K���lf?T߻��[��|acEI��X+�P��il�VM��^!���4u�e��E���R����HM�������
���mFK�5�-������`<���©I��)2%5\��9��� s��Fu��l�?¬�v.�Y�h��z1�id��H�|�� ۴ɲUr���Ǌ���|i�c��c�6��1Z�C�N<�&U0ng�{��j�حΙ>yWw�g-�����������=H�҉ڬ
V)����<�6�- �i�֨ɮ��sg����.�����Jǐ	�=����� @�b�%� $58��֬��BS�4w_Sd��s���ｃ^)o��ѐ!��/>��Ց�Z�����:ݟq�BD2CX�&�4XW��� � I
�@��?�1˦mr�&:`&��|T� ����_Ff~��=
-v����D�R#�q��IӶ�h$�06}��9��FР5x@�����q4�q���WY�m���)ѽ�Hl���Vr�BF���߯YW�D��WR^X�<͒��A�+�����_߉��9��T����u|��|l��<� ͤ�&o@���J�d�k���m��a����z���NO�7����≀]�������?���g��ye��u�Q�O}n.8ڴozW��֍@�g����2km��4q���0�d�ۖ�G$n4�z���wsEl�P��Y��5�h������G�m��<��9j�Q�����<5�?���Pd~՗He#˂� \�u���{��*�{%���
]�y ��ʋ�5M&�)',��
��HPׁ�����65����a����#��k��(�do��4��_,#36��/�(/�*Ң1L�ZP�qGir�$��i�B��A��D�&DЏ3�VF���1J���
�6�+�z'L�cDY�X߫k�@����u��wP'h��4�l�M�(�Cl�^��X��x��t�����e$HT�2�}�ΦѥP�S�Xov��j�_�Ω��^�a�C���IO{���K���2�k�BjA5H�v�QS=z��>���J����S��fHd|��i
�&����E��'�}��V4k`\3�4v��`I*ZaťE�z�'��1!Jp�S�����2\ҀD��
��IL��a��>42n�D	�o�����ݰ��f�7`׾J����n�j�C�T�D-`d�/�����D�,����u#���Tl"H#�b��4���Q��I�H'��YԨ�o��Y�i������R$�fB}�갔��u�93�mc�&H��:��`:�$�x�E)�[X&}�^����^�nM��>ٟ���'�=���ݧ���+���W7Χt���=ڼs+���lP���������9�������4����
$�s�8|���Lx5��������(m��(����K�����p����ʓ�� ��ս���Y揎�3Pg��Լ³<2�UN�W߼Hk ���-�l�LQ%	�e�ɟ}�l/~�DiV7	JZ����ѕ+����� R���L�8EXF�$nu�>>������%��Z��n�UV��U��k���B��M��o�A�,T_IZ.�P,†_(�ty�����R��۷��|��o�����W�s��n\@kc�.�����859�c�C4*d0����,�2r�fz�Zj� �^�v�������x��,�{<�p(!�(�O?���&��M��"�{eO�&�V�z��-K��[��u���0|�<��
�.Ja:��֟�":�F/d�f]]M۝��Yt��	/��s���g�lSlo��#}1!;��v��W11���i�	�*e�F�x��Q���3���Gq����&A� D��Y����O;�Җ��z8L�7I�����f��=W���tQ
�(�z~f��\�[���7�N�Zh�!xf��������-,Q��\���R�N#KP�QG'm��f�k�e<;��W_���^G[���h1�jk
�(�g��@I��*Yf�߿z�?9=�<�u��Wa>��Z�,*&%�c-V�v����&��i�=D�xui�,�� 7�y���!�͍M�C��ƶQ[E�/�JJ��R��A��F�2z���R����S����g�� 'z����)n�ۦ���=c]�tu7Μ1��T�{���'Nc�2�0'B�D��+w7��ˣ�?�����`��?'�4��B���.U��:P(��@�κ`$�Ԡ|.@�i�ڎv����^�X�ӖW����4u}�=*-���ݢ��I��%� ���'Wq����L��SǑ�R�O�h�&�!A���.��!�Yi^j^�����/U"����r�9!Ha��δ��A��՟~�\9텽���Wt,;�}���S�
b�	�֏�/�E¥U��V"�R����/� X�D�����|��i���`ra�h3�)���i^��b���paL�0��RS���`(��H�������"�� Z�F�`=���n���!�G�Y������6��a�y���\e~��l�c6��/������F;��:A*ϴ��ԚId���I'�wY7�fVd'�0~YT�@Guī��yUOK�핦����K�� ���,�d��F���9���l����r�����b��t:��N,���6ЧI3�Vk�+(�
��=�bTH�yg	�Q��S�$�'���]Y�ŷ�D�Lm��j��ͫ/	G��p�駍~��+EH��T�Zg�b�!˔o�V���:�Y�?���8A�a	�� ����=�ę�q�+}�J�(��Ö�E��۟����p�i�'�F#J�'�� �k|�J��F����(�T����� ��S֚V_k9,�&�o�ƕ������������E���3��wH+��^���lR�gۆ�H��{B'�9���C�.���,��8�zt�N��Q3gt(�+7>���=>�0�x\a�������!�z,`��ć������?�.��0/V@V$MW�x�OJ@/ W8�-��I h�M9�����a�;�]���hI���[_�4����r{��:��`i��#�DIČ�?�����_����Y�y��d�?�����P_ ����xj��c4��#ak�J�� �7ѩ���٪&�dV6�W��R�k|�k^uo�D,�s�-�������]��^��T��#���S�5e���&͓�<ZU�y����i�����*�99��$5:�4��X��d����'#82��p����qz>���NL'pb<�S�~����,��tʏD��/?s��R-��D�y�R�O�*i�ٺ�tm/����v_��y�����o"�)��D��:��
NF�P+�fiI2���ז�p�k��I��s��T��;�]�F��f�˦�+S��� �o��W0Imv��i�X�%����s��1=��+ϝ�>��e,�E�Y��v�<h�C:��3�G�q��	��\���w@i`nr��n`{y	]Ҳ��ڬ������a���|�)�3�ӽ���,0���>�~�}\�rM��(���G��^n�[����S�9rٙy�4����S���x[g�?�o��퓣}_"CC�LO�����!>4���2#�}	ٴEu&�.~ʫd���8U"�]������B��?���̵[8��@~o�?��bbj
#㣦d)h2,��IT8^�}��Ğ�^D������<��kZ�f�y3dL�dܮk�ahiy���Ԏ^�����2�]�^�ʭ+��B$m]}�lh��F�H
/K�/ T�in�va����׊�4R�JVw��wh�}����8��wJ�I쵇����JM���k��a��t0a���;���$� N�<�A���ŕ%\�|�4�������@�yI��	���Q�{�f�v�kS#��f#`�s�lʴ�K���#&��4���φ�E5'��ځ�)���;��F�4��Ơ�����[yb넯�m��n�yA��~��@�P�H���m� sՑ�^&[�m�[�5�;�h���ka�mCm���0r���<��h����'x��f�0�?�/�է����Ro�x�(c����:�xn���΍�峣8wr�Cv��U���)��τ���6�N��0R����!��FYX�O��F��E�V���TQDs2�����:_��#B����"���{�L?�,FO�F'�@�q��T�E�M�gj8�����6�F�"��H�/���FGHccx��I���/�9�Y.U����2i)�L�0�_3p��t���6c��\�t�NO�裏��;?�[�n�}�}�]Y�b�ro��}ܸ����w�.��s?q
E�j�ס`�ĩ�c C N�:!`kr�u���de�f�j����DA��r��6]��Z/�l�]�,Z��閶`%��A$�g��$N
Y�1���.\D�{?0+)�o4�7D@�8�z�]��p��/ �:�Ι~�d�B��4+}Ks��q���y�'�1V�y_�s���x	�2��T*�����X��L��?���d�3~����]�S$�^$r��>��N�>I�<�Y���dfTx�V�/7F���8������>���{:&��4`��J��z�����Տ��s:�F�	��b8&����)ac}�4sc�ҩ(&�3����� �=���vvq��u����<�̲b����̦p q[��%�NL EFN�"���1ST��7XFm(����I����>VV�8K�%�Z�����j�w��s}���H�@��E�R�d�n�@�$�Ր$�G�]�w����=TK�>{g� ��^k�̵�Fn� ��8�u�K����@��"��p7�{�^���_��d�����W�d�l��,��T�f�X���t�"�jk��.MTs��w#IZ�M`j0��$0��RH`8�F;���K�L�D��߳-e�,���4æYC�.��Ѐ��rS�t� �h��� �dcԮc�cv��Vt�F���[��{�#�rbz3�v����u,/�d}�q��~�~�Bď����ul����`mm�:����Eh��ś7�,�)�dE������sm˫q�i}ii����=�mk{���wq��M\�|��\ǥ���܁n���piu�$Ө���h|'�V_yCkB�P��P�"+Oܣ������=���$ؒ�8i ���q�V��/`�h��uth��)4���TE"�T4�F�6M�ȯ�a��-FHK�|�Т<�s��K)_D�ә^��h�#�z�:�->�]e�ѹb����r���7���Ir���Z
� ��V=�3<ra��n5k�U�؏C��_���?>�r^D��������Փ�� w7�C��U�:�N��DJ�$&U�����Efce�I<jpv^�~�6�сŪ4m���\� �n�&���ԥE��	\�&�x{��;J����2�f�h7ǬN�g|��?���<��_}�N�/����&W�H�=��YKW���m��D_�$l�+�_��'�G׬�d!2��|���U��U<b�Z*�F,���˱���vx��^o� ]��g�[u)���LV������i��j(�ł�_na(@����������+d�u����`;��n� [�@�B��P�V�ζl�)	�=O���U���m
�e���UM����wL�7P'�ѩ�2�}
�
�-�r��.�Q��Y�0�3L�\A�`��&�ڎ�Ut�1Lf��7i�j���`��M����]쳍7�]��Ջؾq��זQ��@�Zvuw����w�ff�!�%�6��K��TRm� a�b��n�գ1;����@�@����1����n��*����y��_�%�O��������eSPmvQ�6l�N����[[I�"�4@9��z�ַ+��jl��Y4f����rj�+k}G}?Ӈ������`�6v`�!�q@dV�0������ �P��{��CZ�k��=͸�)H>�?�#j?�!Z/�EPo^���?B�B`jf�i�֙�&<()��B������ݥ�@�@�����d<�4�}�+����ʠ�D!J�I�@P%=��r��{���p��o�����9=��9Ҋ�tP��W��pH�����]��U����2!�i͇�?���*�QNqXZ���b��y�wԬE����=��S$�QS��:P�HN��$�F�b���u,..ag�%5�4��Vc��$�ri8:�4�N�)j�x
�h�V��*u|t�*n-��_��P���e��p��5��ԍ�mI5M'/ipKl�$�� S_�A:�FME���:�������E��a��*�]U ��������bpW��x���D�{y9=Ӌؽ�3�n�W�v0��N�?�$F{8�:����6�9;�s�2�c�`�G�C �2l���֭[L���q���j���������\O�/�I�)	Y	&ֽ��b��� �t��6�T���$F~סf٪��T�m��
�7[jm�02�b�.5�t��_��5l��������6�lm��k{m��*��(S�ϭ.ce��T����n���k��6+�`mK�P�c�j{j�1��4%�aی�f(�A2/�lb��l:���I����G?�����=�k붫���	�U����>&�gp��,/-[_�`�."z�'������$)@�i���>�f�w�q�F���,�@ppĺ[�2�C���I�6d����FYIGA���,:�A}�6�L�������'@+Y5��cq
)�(D>�@�u�TB�A���btX�V\O�OR�a��ɸe�Ps�����_�59� ]�WS��}��+�3�f��.y�'��cS�z�xwSu������U�ukk�f�蹺`ԭ�ƷH,��]J�x�����~?���E�:�Yb�ӻ�#���'��Vx/>���r^��4���{�t�#ןI3���j���F`#�[%mnn�٢ZJ-`ג�(T��ׯ���چi-2{&&&�4#i��ʖW�͌ղuٔiB�5�A4���>��s�<�cǎH�@n�����7iN���S�o�ٶ��|���4	R-2��c��4%��:��&��,kd�#N�OЏ#���Ss6`��h�Ma�}���\��S�X����&s�d�zCjI����U�Y�_� P�ךO��`�@�B�O�K_8��)
��>��["�h��1됨K�E��4v�Հ���mn���,g��0s����rtY��8��ǶЌ�
-q7֢}|�.�K��E��F�*߲隚n626�@�픨�Z��Z�l@�}���L)�&�P0)@bQdq��l
� �?�2�2Z� 跷7P����B9���u�Vn�H��NM���J#�V����2�6L�����WI��js�S�K��?��?0�Q;�@�K_|�3�����za*!Zѩ.�8�� o<@]4E��.E�fZ#h��}�&mRy��ҘhF��t������`�B0���Ha@t���M
���������{�m�[�M�#�L$�0=�B+U�)"#���cLo��������ɓa{��i�ؾ��f12��3O��� !���kz���{�{a�p(�@��5v���=������_yc�O��@+
�CZ|(�J���(P��v[1�g/0�tf�c��w��a���u��E��5�L�Rm�:t�.P3��%�q�WX�a���S���m0���W���"v`�7't�?I�`Y��$���}�{�
���i�&QyU�++ʍ~IcPa��LG��͔��p8�D"���!wv���B���2����$ݖv���lE��CR��c�}��uY�ױq�f�~�4� 5+m��,Ab�����e����Ĩ��UB���W1��`��߫SxBF��S����kͣN��k�f/�Uv�Zz/�ԁ��A�0�����ǧ��G��	FP��I�k̮mjp�i����Ф�:b��ik���楺�h�����������Q�h�C`��?�*&��H'�oN�"p�;k0��%"A���w�ֱGn�ڈP' 7z����6�l���ĖYC��+Ha�� :z,��=��V?c�l�Ї-l��z�ֲ�c�5�I��$3�>.>�D�S�k�J�u�<�c1�#1Z)j�,�b*���� f2)LTf2I�fS���R�&����:{�hl���|�uT	썍M�@$	�Y�K�YG��.�]Z����m9p��I:ا�)U����җ0=5K�����07wݩV!ҋ��S�N�# �X�0�@ /�k���ZOc�����4�V
�ffh�X����S8�寠H^��#����>A����j���Y�qW����#�xA�H���p6M����(5���!�ƾ�����ט6���`]����z����g�g#���FmU4�}~���
��y#Keldn�Ǐ#;=�6�D��*b�{�Q�� ���Q�z[T_<`w�W�4�����/��8���;�0P�eQ�+�D��z�_/	a�;x_[�8�w�S��^����U9�9ϊ�3�=?F�%/m������szI#m])�$Xf��4`y���L �3
5J, 5�{Xj?FJ��J+�;��y	��A�`K�u�?�s�[b:!2o<��6�C3g���ŋ��V�V�樭,��6i��5H���X�L�f-�cx0cK��L�Ԡϟס��/�D���_!��q��x��ql,���ͫ�� ��\��
>2�F��Y�j�O�ȯY��H�v&&�]T�Ɍ�����d��E$;l�3S3�LL!3{|V׷��V��G�C����/���HV��_f��'��O�'M���W�^���IR�+zx�Y��7��X��vq{�8żi�S?����^�D�[�4@
�V���J�nR�����@�Z�Ψ��
�Z@��C���-�����b;��Y+PЖ��S4��ϕ�i�@�����`�D��`��8�l��[��[k?*]j��4zlT�tBl;
t_���	)�T�i���5k�Qc���?-�E��?D�f���j��##˧�m���%-C� I�7o�D��y��WpBc1�:�0�Lc}e���͆�&�-���W���m�M'��O`�����[���IM\ڮ@\]95B�VP�����`fi���d"�o�����_`�N�oҶ�������}�.�����޹M����� ��33�:( h-��B�"����c�'�UiO��6?#�C�-���
����^7z��ε
�ѬT
jߌ�ڛ�Y�-�]&�X��̬I2����M�����&F����1)TR��:iܘ�9����sD����O��=0�eJ,������Jڹ�\N�bNؤ� �zq݋��7�i��{�\HK�+�>=FN��\��3�%�u���4��- �[̫����j:fjz�7#CڡU0��� �9�Κ9Y�9�t�x�T9�B!�k�ަ������6�����b�`����d��UW�\6�Vŵ4Áe��*�KZ��&h�X,L�O CMM'��L��������W��������o��Z��N�?��^8G�r o|���ч�3Oq7C�����ͫ`#��Rk=��'���gu6l��hs,M�k�^d�Y�P�$�h/�뒲���eb���<���d���;註A;���Q��[�5��L��4�H�Py��;��BAmYg�h5�H2@�"@>���~�uܸ��)�[TiI�P)簿�κ����e�6��1 �Մ��4u�E
b˖g��)�m���I���� ��@eWכ�w 3���~�i�v"F��ֿ�EmU���^��H#�	<}��^۩6�;B!C�sP�[��� ��cu�5H����G���N�@%�ƊƆXW1}O�����J�]�&���<D�}6���'�b$5�����%��'��m�q\Y��*h��)Z�Yܾy��_G� �&�RCZ�����k4b���M�%0F�~�0�Q�c��-?�2�f��"����P�6�%1�-��Y�,/^E��O�\A����o��z�W����3���c�(,7����d�j�ag�q9o����Q��7��{��W�C==h��az6&�D*��－�ﾣ=:h:o�DD��i�;�cg��⌰N�洚ZR.��_���uOg�=�������PK�=���l��	��\���6-^uު�H��vC?�
s�!�{R��;�3@�EݹZ �x�6-�U�G�):VM��9�<N�5�h�	��/�9�?vϼ֋�A[}bd�ȩ������>��`�z&��釚%" �;��V������������}�at�d�$�[`z�kv�-,b�ǩ��>���9��mP!��~�:��L�[f�f���|qmC�C���ə��`�݈8Tn1Mt��`�͓'�j�*����HǺi*��؈5����J>_��|�����Ԝ��?�G{�����oH���?���� S:p��փ,��B�h���\/�j8��$Z�L˳[�O�� `g��֜�"V݁����M�]۬�	�Y��P+�a�v�A��_"��`�B��n�L�.5΁5�v1	5FjqQ�	������-�1k�S�������`����{�~��u;x$Jʦ	l�^�25�l�ך>2m5�N�PF��t�Z���ے�`�n�����.����p�S[u�9��(ȵ·Mk5"�G����K������sO��	��MR���M�4V�>�|�����+x�����Q؄P����j��% �X5�
ʐv4>��sUj��P�J˅ub��%Ia0Fp{��8=:�.ˠ}fO�J���i�k�Q��_"���>�T�JɶW�BH�îU�X%��)�t(�,Vmz�`��/��[��E!�Ҡ'�Gm0�ڂmm��@v���P�n^���k��n��%?���K���w��m섆0}��8����[_Ceo�Z��~��Q�ֱ� N�G���]|��������(*juY<̋���a#�I���;ĉ<�p)Z��Gs�{v_8J!��J��U�%Y�*�t�pb6�A���DN���5�t�S�X��y
�a�h�eմUђ��4'@W<8m��#�� �=`�2?R��nRhw�;����O�&}#`W7�����V�0����ݺb������9�ꗓ P�{�A�f�uYh��An�.p�WkUlԙ��Se�ڵkXZ\"3o�s���S�;��S��֞�i��|��6����L���f�33��RA��I �4�	T��@m�������1��ج��q�kfv8~|gu<5��ǎ���5���$�3)�}�5놵b�����ܺ����i%Q���u����<�_��+�JF3����v�ԖI��F{7kf��Z]*;Lͱ`]1>>'�H�Y	[�R���+��T���\����P��u q���15��&ci��a*3���Y���&�h�w��NMꐑ�߯����t�~���Q#lR̌���W��`*��/�����oޤ /bq�J �b��;1u:f�(�7���
.\Yǝ�66��X�k�`��0�����UG ���.>�����6n.j[�K]��!�u�F%o�
��Q�z|�L,�O��ah8�aj�#����D��G�@&�4�WZ�f�T�k=l�W���@��%L��(DM��p'Z��Z�T' ��Y���d�}ey�_9�������)��#��8���K�C�V��Q��MG��,�@�S���Ӵ��r�:�yT;j��� �K�ѓ�$.}�Mњ� ���R�j�Q�����Ә>� m!�'�Ti�h�i�i�<�"�k%�_~wv���ז�K����'E�`T�3��ۣϼ�X߷h%ߡu*����1V��
C���I�����
�;%�Z,�Ƈl~�Y�)N$XS��$�s}�������kg�X�B������'ڙT�na}C1n��c���P��� ^���� ٚMw��h��j,_��2~�@��o��x�;�˫�x9�����ob?v9ﷺTԵR�F�������, �q��_'xi����7p����A�&�B]/����m a���JC`�k���'��D:�Q�?�B�7:��w���B�T^3U"4�TYV�T5�JG�e3������'�@�"P�D~v��	�9�g����'�G�ij� +������i��ŮN�aY�oO�#ԱHs���1yl�X
԰�*u����vE
ß���������F�40<2<���)Z"���?51�F�@F��n�"��:�12oۦS���z�z	�Z����LP�	��%S�Nj�(>�ɨ��C M�~bԎ�0B�5N&O�M�ƻ�d[ȶ���nţ���W#����u��W�!�E��������m�xG`�Ñg1<6G�$0�G�s�������P���Ɠ��<u�Sd>ƱAM�jۭ�S�ɀ$6�-�23'�\}�"c/$֓�i�2nd�d2i��dIc�u��Q���Ҭ#���FQ�@(������o0���X���D�2ъSې�۶铲v�-u�Цa\Ҷ,NG�%�?� ���?�EŨEZ�����5�r�h]_�X;*:�Q�UU����"\��Ƴ,/Ӊ�fB�U���M�(�� ���m81M ��_�	��(A	k
'�L��I81��'Nc �D�㷽d�����/��C%l@�|���TN>�����KKX��ב ����Q8��D��F!�� �1O5�]e�j��k
E_K�0��N7 ��z���3����j}ϫ�%��ϒ��vIz;�����������s]>��Jo�,�q�F����T�l�:y\����ڄq�˦6*/\��L�[]������M�Y>���M��늱n�E�Xu[��E@����Ⱥ���t�j�;k�4�^ِ��wwvM���� i��^�ب�u�!��������=�bc��)��έ�{j��>::�X&I7Uv��k30w�����S3S���%hO`ll��t���z����sj��*5ow���7..��-�������ϕ��q��%���Oޡp����%��t�Ƿ�%����7��X��h6mf��z���.�52�̑y͜��z�Ѽ�#�~��_éSg��ɺ��C0& P[,�;5GW{�k�?��޸v9Z��Wq�����+�V��}��[`��~X����\��\7sV����:�I]���
׹�_@`d�X�d��IT��n-����j�]TrM��򋧑�S�'��rZm �	-	
:?"�yT: ���7W�ޅk�xc�y�M`�f�lCx��p��Sfy�\\1��3�T��e�4��d� K���l;NC�7�q�ҭ����v�:�`�E�"s'	�aҀI��d������:��1�W
���'����:3��>����']�vR�@��O#:�Y�aR��������tXK���<�w��6[+�.��2�P��^hP��|�h�UY�}��� ����N�2}�V��+�Dz�%��R1H�������ȘmDWR�%�Q'G���Ŝ)r=Ҫ~�6G�f1:3�6f��A�����#ә���IK�ɞ�Bz�?���Z!
E�U����yW��g�ܪwu/�b������n[�=�^�iM��ƭ@P:�v���Y�뷁?��ں�"�	�M�me��ҫ;Va����ݬ{����W|�gK��^�ڕ�~.oq��坿E�̐�[)�RF���=#�\�Pho�T���
yѫ����~ޕU�o��o��.��i�,��V���9Z�,���w�v]'|���_`f���5UPsd�qšD�8U1��]�;o�f؇yU`�=�����}"ǩ�'1<8dV:V�|'�A��i�m�Y�@V�DA��ۋ�6�Y?�ݸy� ~W��KW/�ڍk���V�.-R�-c�BM�O/�Y�*����+H1��&��?���p������~�4E%�F�)�9y��/�볙>��_x�<���o�測�0�k_�9���:�෴�g�Mje�?�~j�:,XW��EP�r�@�&��*�cjH�mX7C�'֠��^Y1�8��ZLD4v�P��U�/0/ڿF�J�\�&���2��}��z� @����5���8O�Tf�`�M��B����'=P�4 &���]^]���.�׶p��-ܸ���i��	��٥i�LDq��<2Ԧ�<,�Y�Э�T�"_��D�����Fj�|��Aq�H¨ݰ�
A �!6ͺ(�������M
�:5�2�����G��ꯧ�E�Ը��B� ���`�ACʇ��Karݗ ��x!�E)$�'#H~�tP�)PQV�t^��m�L�c|�]j��Y��l�}*G�ύjy>�Q˓&����g��_��cuo�eU3M��C��Œi�Xo]Zk��(x��ż�z�⠙]rZt��Z�-��4M41!�D}��W'��n���i�E����n�]��z����O�-��-S�e6vf^�ʯ�u<�ٜ���
?��\�K���_���Q��y��z�Ca�<�.\��kv��0�<	��lF#ܲ�X�����fv�{�Y�S!=7oa���g�31V��ISW�nO��m�!����������V�k%咻��%% ����{j�����>��C||�"�LmSZ�Vj�źK<�2Q<�*��̙~� ^a�	���DL��!/g�+ދ���It����� �[�n]0,�����h�r������ｋ�?x����-j�Wp�`~�����-�*O���ڴ��\n�4x	3��@ꊑ�(� G L�p��'����W�;����¹/���P��azt#�q�����I���Y�o|��(ʒa��È�/_����}�2��KS�T=�r�[��̫&�Z>5D���I� ��L����Rl�Y��T���W�M|&��mX�a��Mͥ��h"�4�W"�E,3������|���z$ș� ���q
؛����M
Nj��Y��p�D�����=��oa�*q�E�c|Mm�3���'���Ըu�ݼ����������[j봪$��MX\�qEBd\ǜbRQ��:�R�jc~۬��ި�sH'�1Zw=2�F��Ý�*./尕g�k��7+ƳYG=��#P�~͕냺-��*L�fV1a����j;/�����Iq��jeڠ�������*�"O�p@P�1um�Z�Q�����_�f)�~���5�:�!h{�[��_�9���!j�It�V�%0Ӟu_'=5�E��d�4a�δ&f�ن=O��:
h�Es�)�ID� I�^g�FI+Z)���u�R�i�kg�S�[����7A�7�zf�aY�gR��T�6�Aq{N߱���C���]}KFiT�+�(�-{M�e�o(,�8�Nʋ獦�!������w����~ʰ�N�.ӡ���$_vf3��!��`�����#�C9���)����)����[���];kR���������ַ����������h�0jheP�d�tѦ�������������;5���	��1�=�����z�ϴ*K�4Q��s�3K24���`2�U�b�h����67�u!�^Z�m]E{�2Y!E���^]E���H���
��N�&x����v��nb���OSS�c�Cc��~�F2����b�����.M۠i�A!Vw��V���ʹp�c,�X�����i���.����z�#���Cm����i;���7����Щ)��5j�Z�4 Fd��_��+H�$���N�/��/��̌ԕ������LO� ��`��4��ш����>�#��5�.h��va\`�f�Q�����.�]*�2+�
�ŧ"������U��Y<�?�ׯ_��Ǐ�����q�n����O��c&qIgk�������ŴT�5uӇ:�W��n�T�]4x)�C�kCC���WCh�qz2�~�lTc5z;�㕗N�Ԕd��J�ޖy��4t��T�y�*��:�$/CP�~�He�);�k����)i֧f'=��.K��r]�.�k���}��"���C�V}7ؖ��#١3�<�]6(�b���^���5�!H;uj:Ξ=���8veCʋ��K�q����S�ͷ�� �a�d�������\Qc�W9��-�q��@�����}b8�G�ژ� RT�EoC���x(L`�����eG4�)D���ɤi�����o���D���?��d�@<R8hR\fHo�4�)5�S�_��N�� �~]�V�n��K��g�C��s^���>sTi�U4�4�U��5�݌̻۫�NE��5�?ݺ��3.@R);Yc��Ƙ�����\#|��`e6�P?��_��0�����hP���cR}��̜UށJ��:w��xwF��V4;�"Rąt���`2��c�Z��a���!�L���,[g� ���)wΖ,���J�A#��y�`����?��O�p[��_��E�GG�th�,}�p�<n�T�F��IPk�M���r������T@��k�7�Sx<�W�6�sc��W��&�.p�L @��{�#�K�^K�l��v%f���P��o{p3�q 0Ķ�ܤ�5���:)y0$�M�U� ��9�J��,�@�iE;�_}�M��'��4Ջ�����,��Uum�������[�ɝ�q�֝��6�z/�5SqG���C��^0�,����>����"��2`0a�N�hj/M���D'�pd��A#:�1T鈑����<71��1�ލ���j��@{'��[q�������[�g�Ǟ`S5E��'��ܩ8#��Rc����2jD_�@Zq�@��_��G���H��CU��A�^S�aO�n�Ɇm�_qs�4�J���u�O�]:?��qR��Yڕ*��:��^�M�G��Z~U,�	=C=/]����12<b�'��1��̡�?YP����#��A���el�M�ƚC/��[�S�Td7\$(>���<&edbf&*�R�.+<���2�k�:$?I��s�.VTȊO�M�v�)�uY]jMC�zE��K���FX�T�l�o
�Ђ�+��tѸ��ءZ�[a���Ø�����P���ӃڐRTU�+���z.L:Ȫ<�Gl�䲻��ӖJ[�)��  j���L �4jI���~aJ\�s��+v�aNZ?S��ں��n�ޢC�9��,Cz�{4����m��X�{,��Qm�+4�_r��2EdÇ�+�v�cW�R��qqjr2�Fǂ�M��C�kU���T��J�%s�,'7:�j��|c:�J����̻�o���W���sR���Sq��l�9�J,˲@\��$�4>:jˇ>�C����*N���$%�wl9~x#4rU.�-DzV�[x�k��
��Q��Xc���U�`0��'�]oI�fM��ȐҮ���h���@}H]�@ b��iZ��1<^UL<����0?4?��)�P�
�� �Ńi"[{���x)���Ʈ
O�+�������������T�1>:.2���d#��8u�R���oĹ��ԭ���{�bC�к����U	�I��yu���1_���]��܉C���G�yo����{G�Ҭ/=�I��֞�����)0-�E�+�1%5r�rc=��j�bB�G��c��+&h��ףO@�)%��M#�g�v�gkt�}o�3Μ��|������lo���݋�ȷ���7���,-����J,�/�����D���n�a��\���5 ׯ*�ݪO��g����qO�h�D%�O��l��t���D�|~�$4O?�� ����<��y��MhO�Ȧ2&�ў����_�h� 	�cK �����՚j,�j��M|�ޔ�e5��}o��u]qظ���dpG��ڊ^\�K�N��h�A��s��i����'�cKyc�&|n KYi�=��n�4'F��W�|��{^0����4�^)�֮DQ��	������3 @�;]�������Wuo�K����{��Tj�X�Li��3���i��$�G9���eP��XI,��Q�4�M��@|�Ȋ!���r�����	���O�c�rN2@0�;���[W=d�6_���:�`"8ɘ9�<��4j�v�����3�;�,��i��k����]�bz��w�����<����?�k�O�:�xl���@���~VZȩS�lϞ=�dq�3
7����ymXD�IOY�EQ�@
�>�H��9�����,_��W�_2�he9ː�60�/���
hgw�k�`�u�(T�.%����u�",�NrkSA]`��2#�]}%y�{ͨ�L���{� ���c�\��rM�v+6
�p��bH�Ƿ1��u��b(�5Ͻ�r��x%:{b�yWcM@���;=��j4Yf�-�3�A!�J3c��U,E���U��10/�Sg/I댍�%eb7fǆ�P��ee|��f|��s����m��g�^$K��51��U5�l*��`�� c�qTZ+q������z���P\�8������v6���u9��_�7�w�p��v.M�IX�5�M(�`O�y�w!����z�ý19��������-���I�}�)%�V_��m�N �+���ڂ�}j���Gct����LUj�P-���.�R��+������j�f_5�@c�����U��ճa�"�S%V�z�9*��2��J�H"O��_8��3�4%�L�҈�%�%���pœ`/y������2�A*(�
.�����K�/���;��^֏�64 ��J� ���}���T���d(��'�s>j��RjZ�ʂy���@_�
��Iya�����9���!�����+j\z��yg��%kKn��*�28+�%kCyz��?�L���Y]���ȍ0��'L�W���Ix�O1U%{,����9���W��eV�(��l4g�PR�
k��
c�jV�]�~�������dC�a���0N>==�^#˪���a�6�_<�x!�p�5�˅�j(���h��_��ﲆ�=Qn߾�H�Ii�,5����
vhx(������������ʕ+������^���O�9i���� ���Z�&�~u��f�5"�2�i����*�Ǥ\Z,4��>i�z6wf.�*`��a�:O#��*����m��ɇT{��4Z�,qF� �f�d�'s%Xfa�ݒ#x�I�0�׿����=���Cum�<�\t�"-o�[��s��h�H��P��Wa���u�}�129s�_P����x����h;��z��4+3&��te��Uzc@=������3�s�w��8����-�=	K���֗ń�hl-���_�����_Ā�XYX��Q�M�J����Uē^մ>�ˁ�Lb3��ױ�wco�N�<��V��W��\���%^vv���n|v�����Ψ�鏥�m�m�6X�E@�։6΍��ӳ���������Q��<y(m_�K����Xo��ܩ�<7�#�qz�0�ǻbf���rbr�?�Fk�׳1O2걱����`��pQ�>��D�'����P�ֲzs��q|��-�� 
:�0t���{���;/`���xi+� PB�()�:�4$[h�l�'05�K�HpW&����_��-��Ge�_��W��1l�-{��ڕ���w�,>~$PVYz�����k��K��n�5C��=nؔ�[־z��+�N	&�fegF��[��#yo
�+�K�S��n-���٠��Rgr4��s¬�R�x���麴�������_��B`��M@O�\?��)��T��W
!������+%����U��	����ߊ��{O����lgC☔0׹-2��THI��D�P�/,Ba8�'`�����?��$(��|��apOŷB*�]�x�<���U�o�,a�?�Ս�G�P� p����/��'XO��SS,#���&�5 l�]ap�׮�AxN����x<o{��U�˗�SCq!._���	>b�]�Y5_z�5ӵ�����^=����I�MP��kS_��	�.�AG�ȡ O �]δ�
��b�:��dE�z��¾��Wc�y�W��^�	��
��dP�+��p`��[��������]�|kj��WgZ�`l����f]ھ44-{��	��z��\��7 ��� ]H*R]���t��p%f.?o;4=;��XZl�$�T��R������߈��O���/���R,��[�����B�x�)��X;�0Ք�稯����b���^f�{�שaiٍ��pV�=�R���I�Ţ�]+�X̗�6��K���26�������^U�p*k1<2��0�{ �ӳc�?�z|��Kq�¬�z���*��O�M!��qF�<=5�a1�`���fM���td|R�R��fĝ'�����c���C3�M��4S�B�?~]�Ni�l*�w
t����Yԫ{$c���ڑK4*6�c�;'"�m�u�1�&��aD���V��{S�.��Z�]>iث��%�*n�8����G�r���GQZ�QU U�eD���-�� ]m�E�:`nE=�}5X���(5=h�R�h�� v�O���s�>T��P*��9�Z�&��zt\��~dd�;`h,�ي
c�	C�Q^�\y ���h	g?˘ϲ���aii���ܱWu�gg+jjк�	����\���q( ��K�#�����00��J9�Ed���{Q���0�cY��yE�eB�
��?�#�@2�A]�r6Ds�% ?ʗL�O�!�&��S1�W�����t�iQ�`B��$��	�a�"B	øg��(2i@1ap�=9�J,C�h�j�Ϫ7���t#>��eD�F�!M�CY��8��C@4�#u͗�6τ��
�8�/3��l��H#�{U�䰻}"%��5��F�[>�L���D&�졉�bXj�)!�D���ڛ_��VG�z�$^���cY<[��~�=�f���b� ����|t3v�|1@o6�cE�/	��� �[�>{K�nPg�Q`�rA��`_��-��hɯ.!n4��1۠�<4�h�[�
�jx����@��o~=�^8��ݸu���`�i+����@�ҥr�f��{�Ge)^0159$�_���rL�ē�=��P=�I��G=�W�Ul���u�@h���7�%E�Gp]ɔ6���]j�g���1����x���+W����k[�i�k|��$�4ﱱ������>ё�%=<j
a�[��T�8w�z�����Y.X�39=���a-V��~|�A����X��PCݥ
+[=�5�!��`(FZ���_�td��-��=��NU��^I#��2�Ճ�3�C�_����Td�UqE��?W�mW�g���`��1z�`c4>�g�#�`�%_�����D��Ҋ��p�������F܋�R]f"�͜^���R/���|J~�����D*Cl����K��ˏsNY-աk;�J���� y̑w�������W<�@]���4ܼG�l4��C8x|�~C���ć�sY%��eFΙ�� ��l���]�̭�p7�y�m�$+�9��K/���$�c犛����,����嚣	u����[��	�P �S�J�Fc�4�������v��Enx^b��]�]�����.]n��M%���#��K>Hb�<ƛ�޽'����B�_��']�2����ʊ�	Oc��2�3��:M��a���Z]���t_�3��w���]ZA_j2!KA1�&vZ=�Q1����]��K�_�	��$-�]�h�Dg9!�<�6�����3��3�/ƅ+��'��E�4�a�D�U��*x�{��'q��ig�CU����P���*��p��Fb�@V�bSPS�u_u�^<~'Zi8��p��Pa<D���(��Q)���`@z����������s�Q�\���N���1����R��.x�269�f�||�����Ҷ�e�S��X���N�@_W���Ic���Q5�} i��t��Mc���z<�)�R֭�� \LN#��������8�z�.��,b�FJG�x���)\�'OO[=�~i�#J���Xy#��g�Ҁ�h9\PW�LN�ǥ�.Ŝ�}lb��'�Փ<sN��������`!>�y?��o�I��a�F�@���ޖ�]� (��]��Ŭp`��H�2f�]����J��%zOޢYe���4u]Qy���S��>w�v������8��D`,�b��Q5�4�>[@u�� ��4	0�3���͍u)3jH��ѩ��@��#%A�ʺEe�[�l�Vm0/�!wH�i�h��=��HP�k�����O���*�����YvmLKy)������[��D.��^�|X;Udx���d��0�B�/��L�on���AR�v���b������[�Z������^YO���#�rn�e��3�VX�:P��Rh�ǂM���pAQ&,���hLMOK��ahVe!^��Q֬`��0�l�Gg��(c��y>��!$|�"�t�r��o~�;�e2�e�hi���;w>�]���quey�|�!m��'����Jo�L���( �Ű7��W�\����ؖ��͛>T����Ǎ�L��;i\�����"BO�Jc�&�g� �$��%R��`C&�?��)��
$�����1@��ab� ��QE�B,Lb{��i'����9}*��s����q�c]�o���)(�����,��_�3��U�Y�Щ�����M T;s)*Sg�����K�
"e\�q��x�i����R�8��k�r���Z��Tn|eJ���������Hܻ�Q���ů������{wԻXY�ٙI�����d����׾j��rcW�	���=���g��!�Ew��9��P� ��y�_���N,�ѕ�"=]Y�Y��ut&��֖U���3*��+�#�����q���h~E�! Ra���d�l��1���j���{W�J�p�KV�%ヵ�V�C�TΔk��|�7��p|x�N|z�Q|vw��z[�#������!�X�N���ܑ)�\�I�"m��"���^��w
�8�1�~�g�h�[�U��$5�m�z`U����Q�'�y�Ft��V����z5�L����X�B�4�&e�{m���܋\���HP�@��u� %=Y��oF��{8y�����]�]����H����$d�u�x)�.d�:����wt�Sj�L�d��\GY�����No[��{��ءֵEN�~ 9Y[`��b,�?�M�d���!���?�7SRH���������� o!!~� �� g.0r��5Q8��T��AUa�������������e��F����L���o�4Uk����]
?��ne0)z^祋�SQ���"�՝f��..`��6�&�>!%h����b�^V�<���HL����@��?����X9�oЗe�:-{�0.�d,t1��8?�:�l��pj?�&���X6ӡK샮�v��! =K$S��c��3�n`��U!0 `����8�htj6�^~.��]�1w��x�P�
�Żb���P/�@^��zC�Q��U��;|~=:���\t���n'���֢��"da2D�)��pg=���UU���3��fx�,�`-2��6�Bob��z,_�o���s�q��Lt�4��qW���W�;�?�u�wZe) �p����W��U#s��G*g�EOW{'��7��W���������V��@t�+v���O�	`�	vx�]>�BH�@�[њb��2�S�;T��"��/��e�����$�,�œyzv�ivĔ�E:{�B���O�Qog���,%����$e��a�]囯~:�C����z,�m����qà�8�ܟ�F�S=?z��4r�� v�\�z``W�#G(��3'mkz�5 ��Mc˖5���S�����J{��*oE�zm񯡸YqB�e8����9􅡘�hx����;y���4,	��v�@���c�@�U��U�C^�4�33��k�電j ����
�Ӊ����c`��Y�R/i0�u�J~PLC���u>��ݺ�1���R�綰ggm3���?�u'�����Ǳ*wE��'e���M��|m���RDFzU��k�2���d�b���z� �U,�4���K��L&�Y�ǁ�-��.�D�<��(z���I7�9����\)_/	E١����]����؂A�������Q�6c�B�+'C��Y��0]�r�3�djT�����ٻ|�.�sj�L0�!�Ap1��Hi�88�5�Ͽ�B\�z�g�^y�x�IV��u���JӘ�d���ӏ�
�AZP�
p���m��寏�V�.Z�	p$�d
���%�a�� �VTjCq���8}�R<\Z�vO_�J�6T�u�U�a^���5d+~O6֢K]<V8<VC�Z�W^��ٹh�FbO�c��b+u�^���S�x��/�MDW}3�ތa�&����b����H�):��bB��5�Y�c���MH����G���;���/~˼o���pI��;�tY�����>�o,��bH����VhW����L6����|2�^؃��Tyt��NKqo@�a+����ҍ��u�����{c���뷶Y+�K�[���T��>�[�������}5 �j<�&"�$o������ |5$3�l�������W�reK��mi�z&�G�i@M��K[�E�e���h�L�!/��$Q9�hmokˠfeA��Uh�ݪ�ҫU�!`�F.p���Y�ԋ�^�W�P�J`@+�E�R�S2ŇB����G>GG �ܬ�X[[��z]F�9�CW�8 ��G F��5nj��
�l��/ek@�iG�;��ipV��#�$��$.� \���l��D�,�Ⱦ�[Q�v*Q�K��l[�I}s;��q�q���X�o>x��x���6T��>؃��G�VϪ�,_jW$�S��q)"�h�|�,-Ƨ�|j��Qdm k t�}���w�������ʚ<����� �=���=��W��o	������GH���G��(��}�;���IPǸ �� ���P1�[��<{��^���,�D���;�0hج�a�cc����Yqjr�{��u>;�k��9��ɫW�5:��{�쌗N��-%�@��h|j���0�90�1vz�Ί&/2�3G �`�5xX��-�\��F��}Cc��A^ݑ��U�-�J]q�����A�wK�=�X{p?6��*!�r�ʋ�=<M���P�.�����������b{�A�޿����7b���h��ľ4�)���PqӥwAF�[^�7(aKg��!i�?:4 !�F"��v!����O��g>��g�<���3����'wnƓ��9.a����{���T���S�B,��`~z�����k(�6��97i�DE+D�C.y��r��X�4���U��%���a��~O�/n(N*]56�v�3ܔ��hm~aA�|q5�7��mO���X���X��u@qWJˊ��/ƣ�%�����clr6�z�}��Fb~���E��\X3���(�L�1�J�/G\� Эx����Gs�34���[[��0LE�=*CN�b�^>��#? ��_�2Ď��Sʗ��_���G�֐UUz�b�úd�4[�M�!4N����sQ%�+?���^����t������&bC��}@�UZ�o��b������>P����lYM�Z�$�F���ș�RX���6W�b]��Ǳ�P .wK�j_@o�"-��x+m �F���9A�Q=9�R�bH�~z|(NM��-������C&��kz*�ے�'�s��_�%�!�[�#���{l�&E#1���s0�{d|k��x�i�=��e��8�.O�Q��\�m`�3�
�&Щ�-ﳪa`�5���r�.� ���u9�r�ꕸv���>�;^��eD,m��� �w��h�=N؝�{�@�X�_dԹm ]$ƴ�-��ox�c�и��� 4~�`6�]# N>���`��Į�(� �t4�owm0����!,�n�ęs��Д��=�[��[���aLj�{�\���3�6y*��mL(�	H�*K���HZ��%k�[��?�i���V�-��FU�8.�碪��������Pn�*��4k����RT��A�%��Q��ߏ[�n�U�{�zGEʚ����͏?�{�|}s&Gi,��堵�I�鉑h��D����d�n��6cy�.�)/a]����h��/�SC~9^z��`V�lLό�+_}5^z����q���j�k��!�H[4Oضԫ88T�U�أgݕ!K���c�p~�m�I���g/����@������k��׾���Gߌ����z��<h� с���T�F��P�x]�����= �Lx+v���;Z'���_eV��q��Z���P�����k�n�aYV�aC`�R��P|{*�m�)���TZ��]�!���Lј��������$��`�W4�ȿ��� ��P7���5�)���Čz�a���ĔW�q&,t�����޺@�{c-�Ϫ6?�mv�7���!f���u���-��n��zZM��C5Z���Ɍ�C��"bX
�?�UVZ*D ��QZ�_�V]J�dv+�ԃ���u��q2 ��ύ�iF3=\����U����z�n��ah �*��J��=�@N���&�9�P
&I��)�1G�rit�r�"�X6*�x��������J�g^:i���3IP6h��Q~��f7,qd��%�'D�����"�%S��ɟ��|��0ݠ\E��w���PKb�4,�ϲ#�B2���?sTN�����K(Q��U�Jq��3�.Ǵ����{���X��Ⱦ0Ğ�|a��y"�z���DL]��/ǀ �ol*�K�ڪ���I3�0�!2�΁ �_>g����?cgu)F�����/\�׾���l�b�-�a�U��H�哖誫�-��s�n�U�#�	r-&�&ܓ�?���x���w��(���j����޾��܊��n����V����'�F�J��Ҫ�m����uUP��Fw��C��95_�ڛ����x�����g�C2�&���NZ�*_���A�@0���$���I�������
&0��Uũ�zz#RDFF��^�U���W��ŅW�W^W�rƻH~��gqO7s4 �1t� |*)W��{$�=ʪ��||��v��Q��o$G̉ D��Wx	Z9{� kԢ�Tn������[�(0�R�RWݨ�8�b��;�-�%�0�QY䐲��I�*�i	���>����Ǡ0����g�z��g�t�[9��Tw�K�M��JO%g˄&��7� �Y��>�l���^�@{E
�"�2�*[�[@/�T�7h�o�
�4�	�_YF(69�͵�\��BHV�U���3��3��^��Ώ�|��
��А� Wn��s,�z�7o|b �!bU��Pf��Lے�e�o�{�\�0��S����(W�<�q3��t�÷�؉��9�u�ei�B��JbiQH�L������|D(B(I��0�+�;�Q��r2���]�G���R.,,Z3��Z��qv��f�uOt�u#��<���n��)�hw�����3�����4=��ݓFȊ����S�FzD� R���]�[Ձ\��HȿI�2M�Rw�R6ŭ�ގ�jl�?�� L��4n���Ď�lqk/�w����ǏI��H|�XdOR���V�.R��� ��7$��a�J�W����k1sf.��C��}��DpW'c��@��׫z��i�� "�M}��X�����@}&��q�Y�1T�X���$6�c�����XR���J�,�ɂ蕭�_ڒ��8�^w��C�����2C���T�T5�cxt�.�QU�T�G�ӧ�#��j jq���x띟����!2��-y��Q�(_7���G<P%�7��Z4*�c�����},[��a	j��e���P�d���l+�2�P*|��-wC��Z�m��iX���ahI%���>І!��_�O�N�SE��4  K�����Lu�\*�(l�'���v�N�̝����Xݭ�F�%�'���+�T&ݲ]�++T���$+��0�!�Wt/g�ʞ����/@\��!<6"���`��P�����K��*�ܘ:]�N�b���fdv2��p%ΞS���jw쬯���݌\H�V�y�������`T�e�����䡛�m�i����R�c(��'m)H�Hz��2[<ǔ�Y����f"ˉ(?$�
c��O��%�	�"�.�[�����HN&�[��~_dJ������<+�4tA�J�!y��	
+$�C3iQ�,e�+sV���+O�c�Iډ�X����[wnKH[^[
��n�26���ֻh�uU��Qiw�����x���MU$IM[�[Uƚ2i9O��x(: �a8�s��Wh�ٚSq�@UT�[L����7⧿�[�<�H3^`O|ic��J�^|5�_�i�[]��W�s(���b����P���zC����v�����at�����T��q��W Hf-����|`-��;W{/���Ҷԅ�Z�0�Ό�'<�9)Z���\���<��nt��V]�]����c����rw�	p&��/��ۉ���`2d��M���)U�ab� �F�~S<�9K�4?)K&�i��Xk�}4��{�����O�Q �>���n�ؗ��Q&sy�۹*�QJk�g5��cx�=R��$��Jȡ�lX,/�َ.�uH��*s�;r.����C:�8��n ���N-(���������[�@�+.�_�tQ�׌��Z�z��u��oX���$�S�����8%H�+Ý{J�U��Wߌ���k�93�j�Z�CQ?`�K<ٗ7<�����Ij��-<,�KK��_����+���W�+�\]aD�{�Ρ#D�r棹���WC>��D7�����ywǀ�w��;������c<z���*4��W�*����/})����K�a{szI|4�ٝ19��㌊�^�z��w����>�,���9#�1�C��E){L�}%�bp��b"֍��C>������с��6��ui�p�����E�=/	�>CR�|F��0�U 4q�;�����*Vsx�U�>=c�����ӛ7�9����X�BP��R�.&���ķ�׈����7b+zc��|�|��m�!�?).��< ��瑶��Y���7��~C�,j{�q�����G-��z,�ܖ��5<�31r�Z�^y��,m���ؤ�6:;�����lD}y>���؎a���vL��E=�f;���c?6���U���9Ң��ᾷ�ý�Ú�P<���F�j]1>1 M��7΋Ue���PES��qP���A<����!-}���{�-�McL��A#-.���Q/�*Y��b?�|��������AGp�������|19�iP�=%��(*(�Ѱ�^�M���r�l�����.4ʘrUa)�Tf؄��:�w<�HYK�XI�aχ�zt(�}�����s��Or�Vޭd(zh�@�Dn��c�E���`ȥ���q�K��8rrzʽ!V��gxO�g(BQ�	�Q4P��1s
 ��D#H�u����1<w9^�[/��{>���m��O�N�A4w^n�����X�)2����\*6J7�d��aiK#����x߫�\y�w�XvM����7�B�����ӛ.u�����Q��F�s��n�������;?�i՛�֞����q�����W�K��a��reu�<��fv�����r�d�2�6,��q�����7~�s��O�a�,QƸș/�s_1�$�0"��"�2 -e|���!��E��,���	㖕�h��<��5��/	�U.R#ׄ���![	"�d�AdB�10�`�3cι�xߠ���  �O�tU�B�}e�Ү�x�^;T@�W�b��s1y�x"P_ku�VK�S�TI���t��3�4iT��7c�Иy�Y�;���!��U]WYs��~,��,���P�������Ћ�^��Sgb�!!iJmن�,d��*��a�q<��Q�'p2rXUpO�>W��=Ҷvģu��%�������h�ѽh.<�7��xj����qjt(&���论��c{kUEӊ��Q��8䦀Š*���m�nǦԽ]�tZ��,QD�.e�JB��òd^�c��I�֚�g�ZU��/���݆d@�Ј3T�p�p��]gi�D�ϫ+qVmP!؂wkkS[(����}Ƅ�Ð:�-��d2{Z�̑N��4�wb���.�!j�Ќ�	����T@��zfzdv� q�Jϵ\��نԸs����J-�&�akV��5{!ǀ�(��fxE�D�W�wy�&uIV?�F=O5J�%z9�:[T����f�M�ŗ��ߏ��W��nM9�P㽱ӈ-)h롲q�Ky��SVȰ��A�I��B����!+l'^�%����G��r�8�gY1dm��� �٠ >�ߥѥq��)�u�����4_�6v�{���G��wb�]���u�aA}ϋD��?�?Ǜ_���b��q�ʐ�������������gj�(Vlc1_�ʗ�_�zp xFy�Yy-�^�LY/����.�J`gH�4I�R/w�Ǒ-"Iv;�7�V&�E�D��8�/6O�q������י����[ ���E)TN�a�m��窪 �v��8{n�]4V����� ��d�������^���pe+���p��]�<ʚ���̂5-�(&X����4Eݕ!��}�
8���Q�v^�6r�b�\���������C4nF�Ek�^^D%��^���~��G{��l
�p#���U=CL���E]i5�c��'�w�����:�������z1C�bƇcH��	.��={>._�����O?����Z<|,mx�.��j��h`�(�s�*�F5�|,D�Ǔ�XeD0#0�F�6��z��eۀ]&�vꊷ�sU��f�@�mnɏt7cae#ַ8{Ҋ+��#u_�:C9��Q>KPS� m����K�KJ�UO쒘C2��WP�%��0Ѫ�&���_�*�E �3�������a�{厍�8��5`�2Bܖd�1x&.I����裸Y^�p�ϝ��q5��]v����ce�����ϓ�<(iM^U"��ʧ����T��ӧ��t��+qw~)nܹ�I[>R�I�W�tHKq9bY�ݳm1Mo*��=�Vx��c�cx��md��O���%�[i����ӧT7�6:�g�@���aHV)��`��%n�52^+-d�V���x���x|��蒖~XWot�i^1w��9<
+���K��Q����\+�({�L�?($��>Óg������ŔČ|�tKS�cK�Xχ�����w���K��k3`�|�$���p�Ia3����q���ω��ʏg�:�MA��O2�t�'T�]4��,�"��>��Ę���P免�?�������nRh;��]}q��ע�6�Ux��9Ai�NZ���`�
?~�v ��E9����C�Bo�;���9���Sg�otҟs�+_���;p�(�fy� #!\WW���C�Z�[K�1]c�a[`����(�pƪ?�Qo��!=l{ë8��Z��<$�U�.�-��&]����8�X\ZWu>*��DKV#[T��*�Җ՝g��C" �6�X��G��s�9e�a��̶E?S���a��{�\8'u��RECC�n��W��"ZX�" gE��{lR�ǒ�N��i��ǜ��|%,f�i���5��d�����]@C��<y� �}�i+,|y�/��PK�vt�p�W�G�aEA�v�?{p�ߊ�&��J��&�c��tN�r�_�Ml�1{$Vy�L(�Nk���1�
6���	�H���,eL`'��i��ާ��~�&A����������52=s�S�1.�|@�������*��z~=��%��ޣI��}����VR-�+�XR���i�� ��Vnފ��k=���#�֎o��/�sW�X�Cy����e��j�N�7?��|%u��;7?�̍1�� kf7q��"��υ�����Y`?�C9v}���wI��E�J�x��	/�˔gN^kBu_��D�Ϗ�N>�F!_�p�����
/ˡ�hK�&�T���BEsg�1B>���a	�7�*X���#Գ�3&�bb�AC-�4x��ֆ� u}����^��ΪI�?�]v�c�e�6����{YA����v�[��Pk�����RP�\7�s��/�OE|~_b�qݿ�q����cH�;UY.��ŋ�&����iz,���Ĉ|F�a�%��(j�2gy)��-Vc��-��M;�<���Oo���k��{h|bZ�0 {���J�N>��^<�O%w>D!/�G9l �rg=�.�������U<4
����uU��P�<Cc�16}&��V^we�Pت�!~]��w�h],�������Wà,0i���ȚW9�׈jyy���L��K7�����u�&�Db���M�*�[A��d4?(dh�5Թ�e�i�c����E��dC  �=�KJh͢�"->@bU"|^V=�'���9��)~��d�ɰ�t��Q�9���+E�m9;j�RVFctf:��N��ܙ��O�[�V�թ�b�yn������?�СӮ��K}��U���s��� ;�vz���.,Ƈ�'�q�S�D]
�N\{�j����e�3�P�K0/�= @��¹�v�e��0LtR?��7՛�1�*�K/9�E�E�\���I����f6�L�s_>Ô�v}�;����^ĝ�9�xڈ��L$��	~�q��	w����qp���L�w����S����D8�f�{k*��Ukduiz{{�r�e�ޞ>��R/�/Ξ���[S:ݱ��+mP��d���$M�\A����=6
!aJ{Lc�ą��;�UUA�U|Ya�m�t����|���<�v�5�[�>�t_�z"�O�;4lM��
31}�J���ɧ�����n���kEwǾ�anm,Z��R�ڃ��?|<�<�;��K��3��W⅗^���#oG������I僠{�"�v�`��0���x�L;��S�����G��fKY�r[�[o�p�LFmh,FƧ������j��Ug7C� >��Jm�P�I�7���2>��ޫ8X��~4��_~mɘ6�K(r[p3{h�����2O���,��Jk�0��!BEl�u�b������ -�`�W��Gꝙ�eJp�r����״���SiЈ�����I�?�y;{�ǁ!4���M�/�TT��K�PI ��K<���P�NM���c��:}*f��ʞ�����w)/��r�*l���89$�.x�И~���t�u����Y����␅"�@�x뭷bg3����q�KR~._����T�U�?=��F�/�9S�3KK��� ���(,{Y1d��+/�k|�{=�Nް2�Å-���s���^�������^1�)=~�)�P'"|�P鋫/S�Q��y��ió,�2]g�?	�����)�
@͚����4w�V�"t����u;�bR�3�CC�������x��$���Ě@}ueO�Is�wJb�2M��H@3���Tɲ.}�މ������d�ä�_�I�(o
���7K~p'<p(M��V>���� ��`o�mG��+�.�ٗ_���u�{��"P���9�_���,�?�7�I��!I<�}�~,-/����3��կ)^y�J\�zA]��x��D������������xH)��wZ=:zvt��Kٲ��p 3�|r��}��{L���\���<���l��~�n`ge�
zK�B�Y�¸
�=�(�W�'�Fi��>�00��"�O��[�d�v�ii2�=��GV�P��U0�/��"�elm�u���{|�->{����q���rS��^S	��M/JRm`ЍyC�����x����~4���B�=��K �����X��;��d�:7�ϝ��T�����qz��?X&�e,b<�(�1�{L�h��عuT>��5|�L���	,_���`��.v#k�qjb@J]op`�z�"��_	�a��1l��7�S�Z��ݰ�dݔ|���!���1���_�u���=�@Nr�=y�!���O�)	$�2n���Ҕ~'�e����e�:�.ː����N�B����r,����oKx�rǎZ�-��q_O�P�{b��;����7��>Y�퍺z��,�Spu�JM�n�=S���1h��6���H,��S���o �~&��+-C%'J~���5В���l���
����R�b�����ވ��	k�= ����j��@�W�;�U9(� 4�R3*"k�g8�\]��gN�&�ԵfWL�-�z�z��l�a��&7)d�P|:.G�F��/�X��G �4��3T��=<�����E3�Y�ΞB�f�R�vc'vՋiJ8T�\�����{z@3hC�~�Ջ �uϳ� !�I�?@Q�hfY��۲��aa�;�~�d���ܲ��p��4�7$��� W08y��L�24cmO�rb:�S�&L�:�;q�bK#��O���N�L<�M�DWm86�+�f�5���C1,0���:{&&�ӧg�1����i��F<���4��p����KJ�:�_�k#��h�W�,���.�YL�я���)k�W�WU,C���z��wn��ڼצ�����S���� �2�4b����k����jl��"2?������1�\�� .˓m�6V����92C��]�:�'1�4�Ɂ��ʄ�Ȝ|v��c�s��f5ʻ2��
ß!��
��::��5]_��n*k@�!�����w��Ȁ�H*����֤�+�}PE�=?X�����b���)p ��b�����ҥ�\D�С�����a�	
+?�����Ea�'�Y�%
6ؘC��4�V�����Fmt<jӳ��\���s�[��#���HSߋ���x���8��l�	{����}*N�� $[F�^whd$�y�G֨��1=k[�XX�ǧ������m©�'2��Rc']4:����H�82�7S�eYj��W9��N0q B���;��s�����z���]�'�7wm��a�x���u:"$+���K�Rr���+{�vT��e��X�)�����y�a!M.)��re� eϐ�AuVo`��[	�VP8�Bq37@�()��o��5��JɎ�R���{����͜����=u*�gN���x�FWo� �+^%���
@���\�Qp9����C)��`�I���%^��p���WX^���s>Ku���	�P�X���W�8"�n�?��Ϯ��@O|��W���4�_�䉺�]��7ӃG2%_��?7]9��e�+�^[���M��&��~\�Ӣd�.�)[�d�r*�ˏ)�d�mO��2ხ�|��]�N?�хIAO�yN��Չg�9�W^qx�aWϼ#�0�eKq��Ү\�ХuoQ6S����P���ַ��U�������_UW]�B�����aD�+ǎ�q֨�T�bTZ=�$GkGv78���29���t���<(�?B�i�"�����8�p)<~��̉BK�t�����RB���蠺���8쩈�ѭ
ի���	�7bLJnGc+�6�s�K�F�`��{ v��MI(�ٕ��d~�ix�M���݈�wzo��޿��Ǳ��*� �3����� fc��e\1 u¸T��?�+�I��J��ĺF�e�f�����@�5�����no���+�@ؒ�wI*�4%zNY�s;����=�"7�ϊ].3*��cHp?2�����=;���26`(M���h�b*����C�u�v^-��^D�8ӥ�����rP�ȓ�&W�cG�u������K�����;2��z�����U^z?'<C;W�Y�[;�_�%�eu]ʬ�(?���Ks�"�I[�Ϲ��.����މ^�[�:!'�,|��':�/�?y7|���|z<^{�j�1a�(�{ʈ�u��� y�Q�4޾}G�a�aXF[<R�$/�5>�c]v�e)%���^A�D�-�N�pZ*��t�Ƀ�o��o�&`�e �����/�ka�[�Bs���N�����Is�R/+��L�0~�?%�D�e�����_��1�v�I��ojj����+����e}��]~�4塀oX��ܥ�qan&^}�851��1������V]��Á���5"�|+On@��!!�bY����nʺ�3��L1��Fɉ�W>r����P<�A�x��_Hѽ��E�g�4�^�{f�/�%�竼�����AO���jo_����{���(�c�+���
�ID>�q�N|z�ܻ�di%V7�cs�����>U%�jƄ)_z��*3eo9_uY��M;y�$ �.s@��m,K� �Y#Zۀ����+��L�mYaW�����u�[Z�q��O�aW6+��
�,]�"��(?�	��d����O7��ܷ���ܲ<#B+"y�>`��»���z��M� o�ɳ�W�>&y
���/�΍�X	���ZtVj�Q��3�=0�ڸ Yo�7�W[@֎���#&�x� ̱��&��!�\�9eϽ,e_Z�e����]e�Y���*ը�?l��)!B�)?�5�U/nX=��c�����3qvfR2��8�	�W�2��)y�eǭ.��������e��E�S>h0Y}����������I��pO + :�.�N:�W%����6�%�a��o���=��)Ý���0s2���)5�����0�2�}[���;[z�(��Gz�������)5�������W���.�wI��#: ;^���7��]��с�pf:.��0L���
؟��.~�L�{�6ٞPڽ@���:���w�!C�z$��g��3��|���VE�
Zo�����2d�
�w�%���O376��!����z�M�����GObS]��'�..x�_���d��O����Jl��Ʋ����*��"`����F&�=):�l��$z* _9~�ʫ�c�*��S�Ѧ�ō?�I�(L~�@�ķ� ��
[t��+�Ԋ�=Y7�%N����4\��� �e���[�о#@���*MO@P�)�(|��(\F��.�|{QW��R�@i����!�!l��X+��W��JA���*��/�����W�����k��kh,�,}Գ��d�@/�ݵN������e����=*��O4XQ���\+�;�M;w�+���bP=�^x��{K�q �mJ.�ջ���Ⳬ�֮�XS��P��W/�h�2��͌����EL�#ҧ,凼p�������	��A�^�_R�+o^x�y�=0�>���5�=���p1�<å�ʹ�����r(
�_�wd|�x�Hq�#�X��t�?N�4'���&��!d'_��86}�p)hg���|����VK�{k��������T`ʱsh�@��H�(oE@TLr�t;�1�W��S�Bd��V��%�������ĩ��W�P�oŠ�Ni�����TAm�F�mD�@�{��#z���2��˚�*,�,pd��M�X������S ����YQ�KH��GT&��Qu6�b�ލx�ɇ����\[��M=���>�?�>;;E4m�0V���f�-�<a���MzEҰe�QUr�����MnH�C%r�EN��7���`H������f���?���Aq�ו���b06�����w_�~�bN>s%�Ge�[�"����X
WD�+�f�|�ȿ�ʲJs���!o�D#Ŗ��OLf�%[e�h�L�Z�^S�F��Y���D��h��TM���Ĥ�S��N�����s�º�x��G)�y0��Z�,�Q��2	�z�HH�� ȳ�3Y��oZ���FH�r�:�Gx��y�ވ���ē����q���~�gq��K�Q�U�ة�J�U]<3�'�'&Ńp�Xkw�%}��a��dH�G|S�>��#�)a�#���#�g��g83��c�?�l����{�'��yiH������ �˟=��_��@R�=���5���'/M�Y,�OƑ��&����9A��
O\����yE��Ni�4�+h��Ҫ�t��Rbi�<�z�n<,��'ǉ���GX�2NNe�ح.4|�?R���@_L�zc�k?�z;b�Kzc;�F���s����HI[f|�͹�t�K�]���1�02L����gX&K.�dޓ">��Y��+�B�Iѐ����뷯�ڣ��4?kk�.�^Y]�]�f[+�����3E�:6՝d�:��Y�\/��u�	j�}g�
_n�/�dC%=^B��?��g�WY(\< Oe͚/"�)`�����<�6&�,S/'���h���TZ�������\��M�I����Ɗ��*($@��#ԏ�˰O%��#o��q��BO�H��� \����<@���Bxh�a�(�����\�����ٹ�n5R*������ߑlp.+ �\ ȔgC�x����>Y,ŝ�A�*I�x���"�K�fZ�� #�Y�ۥ���Kʓ���~����{wnGܻ+{'���'ў���s��P�cB�2���{�J��"� y�|M��'o�I���A^�fH��������#<�p4��8afz����\�r��-�1G���x��R��؟�@)CA�ڣt�#��bH43M���-�)��u�y�d��F$|�g�5��R�U�JqO�.�� #Y���{�:�b���yJ�+=���J6=0V!�O�%Ka"����������zԽ�sS�q~| NT╳3���qef,��ř��Sbjh(��D��0K����m|� ���q�_�˶ȕA=?Im�GT(�Ֆ��Y����§�ޓ�ѱ��,��ܶ������C*���)��}�1�*= �/V��5)�/��.+Y�ZU[�A��|��ƕ
�SX��އ7J3�=
7<�W�{l��҅�\#c��i"=Y\�-&��ȡ�~���f.)�䅸���{���C�]��6Ed)�ܜ0�� �t����;T�����L����x<�� 4g�����h�S��W��7�����]e
��m�������H,omD����es⏺�8���[ɚ�l�䛱o�$�
�-�#{GU��Q��_��Ĩ�y�V�wtJ����\U/�V,}�O">|/B�L�LMFF�lG{�tpJW�ޝ����R_�<���wġ#~�l]q!&�0�A��aE�ǭ۷caa�e�p2���.��akeN�+��3[�{�5x�	���ae)d�_	���@bR��.Q�~��}^~�)	�@d
d�q2��VϠG�<�Y*�J�
��-�#ThI0��T�=7�W�.ǲ�f����C�eu¶�����{# I�c�KfN���������Kӯ�t�Xo��Y��h�)���	͎�ǩ�����\-���)�����<�g�����4[h���<2b�o�΀�������'����Bs7+�������%��7�u�!CQ�
�h��P�F8˲q�cm�q4�����j��6��O$<P�H�JL<���2I����P�a2]��o
?����,A�]�".�xZF���=JV���(����:�<Xvt]�\]Pn�������#�ꅟ���_�y�4��+\��4��&sS�ʍ�&Xn�x��)c��6�vb�ь����U�ڗc�k+ޔ����n�n����l�r6A����ӵz�r�Rz��pd����^��n�AloI�؎��wb��be)�*=Qc�
��kxΪ����?��[7%T��M��uJq�<
|'�x#N_�h�ʭG��h4���P�B�B\�f����O�ćh>�C�('V�ݿ?n޼��c�E'�s��+���
Oφ�<?�}�5�n��p��Sr��}Zc/Ҳ-=6'*�bP�_�@@i���<��=%�Ĝ��e�Rq�m)��	�p���c�����~�҅X__5ȡQ�n�zĨ��r���8f�;+gkH�<F�wiUUU��8�ś�>J��	��
�C��U)����]����b��_�zA�J������nu��C���ֵ�W��)�Ҭ�IQ%R4T�n��}��%��b������H�}[�B]f�IyPT8�� kX����X��}�c�)V�ŧa-�`0��� �$]�����[���j PA!�G�a����O4|�	v�ʳ���.���GN7�|��B/1%�E@��[�!��uq�X]����O9�[�U4"/	{��\Ex�~VX�"�`�g���.mʂ�,?�%Y��\��s���}�_º�V��{�;�L�C9�v�I�ؖ��$Lr�3G/��mn�{��GҌ��1���&F����m��Rby��{��7Ύ�DU�Z8���Đ�z�V���N�޾�?�i,��V�ݿ�[���T=����g�!�Pꇭqc���%�VVrC(��!��_��/�?�w�vԦ&bkw3���90�V�S�R�JqH$l\�G|*�I�KyP��> ���X~�������I��[��r��k�RO�w���0.�uDօB�9�b�P�e`/M�(�/6�Td �I�ֿ���z�e*S�0Gπ,��(���]�Kt�����٩h�nE]-?�+JP<����z�P�͡u��Q�j}���P���UT(� 
�cc"˙��ҕk��窏(g�eYz�$�*c�]r9�a|�?����Z���G���H�'�������5�!A�J�<XK'����Oy >��fic��ni�O>�$�7�K�7�rÚ�A6�"*@�]�K���$K`����/BGyύl�8X�km^9�q��)mu>�^��/�ł��[��Ӏ�����K`�Ra�LqZ��|U��/���e��ò]�L�P-�ЁKp�8��}���yq])��Pq�gx&?C�QPGHD�ަ��g΍ӡ���p|��A��=n	⩭g�����2�x��4��,e��B>��}i���r������F�U����k�b�έxp��x����p�F�����>��������Z����b���l=y��E'�te>��>x������E�3ߋ^1�`k5܎��Z�M�) +�������*7��	^�*Ei�t̼�r\��_������g���ގ�+�bg3Ԑ�$� ;�D��F�������3�&~��~B<z뭷R�s�|����1�G�!�-��#K8ʁ{d�:��AKwy�LR~M�G|�J��Pĥ��&6MvK�Ms��Sa��O�Q>?.	����2�eP=+]\�R�^���ܯ��g�zJ�.�g��3^�|.ݻ���z�4ޣ��We>�_��N�2��뱱au�����Bc���8�_a�A�	󩿀�����U]S�/+9�]U�
����ec����K`.�{�-xnP�{����h����n�`�uW�����Z��)>9��L����4����7���x��E��q�CUE���	 T4��l� ��}uW�P0�`KAG�	�@{�Vw')&s�P
^1�j���n$o�y���a��ϲ��"'�	=��;���ojs�����%9�p�q�d =��Vr���)?@�[��1����^'��^�H��z"�EXH���r�`��M�J������L]��H�x(�
Z(��<�<p.�\ev�J`�e�!_�sK4�|�S��%o��rH�=(3�A��C�9��ђ��a�c�U��ׯH���8=w6���'�î�5&Ƅ�{�#�4�V�]&�G���ږ4�o~3^�[�Y�L���QHn� H�B��U�| ����� ��bxb*:k��xs#6$�z5���1��(.-�Ǵ�;@��2o�_�(Zy�s�%9ᰖ���N�����O���o�-ꭃ���}/���_����+.��J#�)�7���dy�g0;�w}�7�m�4��l2�YC�z� �*���q�Gѓ��+My��`��%u��V,�l�g����N,nlyp}m%j��|�Z������ ��hQl�kYi ���\�3f7 8w��UI����N��$�pm�0�ךr�����l~}�\�=��Hh�^����.&��1:�����7��F|��������=͸��O���c�^�����1~���g�N ���T�{��8�ͽX�;��}e� �����6�� ��^���G�@9��4���(wD��$9�����Y%9���2D����E��OS��I�p�
�rP�	�I�C:<q�q���CG��	�RcʼCC�Gi�V�,iL�ld��<��D�.M���Z��5��z��?�#�Ѯ�q]�5pە�%�Ua�sS�٪�$�~n��8�Ս�2<ϴ�����7��?+�.^�g�NG�o2$[��7ꬒ
��K.�?*���6�<(<ױ-��ي���\���Ui�+z��p���|O+�Da��ǃ�W���6�bC�.�,���j�
���걩�G J�8��U�OOϨ1�A���3X����ξQ��ݨ��0Y�� R ��L�P8Y@����L���Ļ�\��WCr����`��GVP;|���S�1<<쥨	؈2�u�4� I�i�D�S�w��o��w�nLOa�#:6Ǆ�;\��_���7O�������2�3|��ɕ�����m��/ǽ�����b�[ݍ�K�$�Y]|��(o�|%N�Ă�y��X�����(��v>Ғ� �122 p������Cx�8�J��tI��l�C�\��'N2�F��*�_)H�)���!pg��.-�;f&b|�*�ދ��z�p�R����������ߊ������?����D_w�����2�.�p�T�/��BtT;bPo*�uW����IaE�A��=�|J^���ç|�La�P��	�^��E�J���Py���3��$�lLJ9�5����"b���5�I(�y�S����k@�~�ܐ9�#��.�H'��#�}�*������G�e�x�{�I��/e��r�����e� ��*�r�Po耍ѤAc�KZơ��ā@��Y5Unv�aj9���x��â�{8��~*����s��WZ;�LLNz�zo�A�
�n�lBXe>���K=k�L���#�C�$�nZ�-�c�f˂䘳h�ؘ�,7�j�c��X�_����X�v^_���҃�����ͭ�P����D���]u ��81��%�MoY��Xd!�v���Bv�u�%�:T�E�X^^�AJ�P
dx`����ފ��)��JO��laS�B��-�bz��eZ�woLn�o������Й���2bL�aJ�����8,N�̳�:��ǘ裗Җ���"iY1Mq�K��^+n?����+��݌-��MI>{�t����`O�����폕'�N	`/�� �@���L������Cڊd�ۻ�* 	��3i�^2��*X�X�`Gs'�N�<F��뒠�P�{-n�
`��i�cg{-j�	a�A�llĀO�"���Ƽ4�mK<;V6�]mp�4(@�Ô9h�-�o����O?R�hW<gX�<@-|�*A���E^�_��#��i��Ï��:k����*�[ ����]4u�ᴑ�	�O����,���<��%�BN�Wy�I�SآRb����.��p�|Ƹ)QCo�2�0�3��C?"C\䵤I6�U�Å⁯�S1˃h<�W^�f [Y=�O���¡�w�@����ו��!_�C܅[�c�D�"���xΉ�5[�7hW��h���+@�ݕF.Y�����/����14>��*N��3���̛a�Fig�P��
"�c8�VO�zz
�0��c�{kq)KK�����o����><cuu9�oߊ��?��7>���������`3��z
U5GC������у,d�r��e��(���J���
�m5J|����/�+x�s�+��x饗���)�:mxV�?�/�61K�y�.�������!̉p���o�0� 5��)	?����ʂ}�5T_x!	е�]����,�݇�>۲�Q	u���BC�9��T�#�t�lLWc��}	�E񔩕)�'�I��_ Ʃ��[md0*�=��Ǌ �dX������-�Y��a�W�"=�>t⣧J_\�f77�f�&i+k�����Uw@�fCB��nitǧ�܈O�%��q�Muu��z,<~�N;��t�AhooDsc-�o݈X[r�q���9��PN9�,KŃ�B�D{��xIw��sk겹J�I6d�x��
�VMU5�Z
���*�RF��_�_F�2F�u9eA��L���q�!�rɽb�Z���t�cY�/���r-[<��R����1��(�V|��)�T��3�V��.�W\`%/�0C%�yj�<��p�!ؑMg�6l��`Ox���W�
-����=�ߡ�\��]_]5]��������8Ӏ�O�c�칸��W�Ե��(*�ñ��[�9�|KХ�T� :�8<=�	�luͽ8ŌIK���h�Dc.��$���6�jt${���������b��Q��|ԗ�������G�=�0�7�쬫���L_o���{�H��xv!�.�4	�JW~)_�皲���={Ǽ��;�.E��P {��hQ�1<2������C��v��Q�S� p���Ezԕ�ߔ��%��D?g2�Mqy��i���8O�e�'M�Fn��d�Gﻤ�9��B����n<^\1�oIs�������I��z�t��ا��b��	��J��m���H�5�<hֽT0�s,G����R�DUگWr��|
��,�"��.�+�nU"
֛[)��Qn���㍆(_�1��.�$������U���V�z�mOq��@E�F�?�~=�<~N ���K#�ڈ=����n쭭���hI�UdT	��I�h��»r�9��P�pY�d����y���t�Et�m>կ�1	�ֺ�$N�'(��=�&c!8|I�㗶��;Gɘ`�t��e���Py��Q�S����?Y�r����@^��%ʌ����y�iq]=�C9�!��:�[���+ w9��Yr�r��lm]V�k�]����,.� ���kW�&���[�,zbm����:o�V����F�̹P��{��l��G^iJOi�pi�Rc=�:���c�Ko���l��;��3ѥ8��9g�n�h�W��h梡�_��z��/�g�Ryi4�2�`����JqgX���;�q��v�z�q��ƃ�1$��l�Ā\�b�2�E9���W_s�=�WC��ؘ��C�QM�#q*�K�(�a�7��McG�e݀a�{}�c�
����r��#�=_2���<��)�).O�<m��1A�7%!�y*�g�-��-���
3^\ٌ��=o!ڒp���^�UZ��s15R�'b.�%��T�>��c�Nkʴڌ{d�,¯w��� |HAA��(q��*���*P*-��P�r�:I�:�P�I�~(�N5Vq�--�[�Ó6�j�`�O�u�#��ޏ�돔X�+�[ ۡ�T�X����%�c��m��+��\�#0��Ҥ�͈�n��@�4x�L�:�����!���g��	_s�IQ*5��1�C����&�˗��$�'Z�q�ɰ����ɓ��W65+�9�c���.���ܴȕ�Q�V����t�*�'��_��}I�rx��Ӟ��J�l�.�YRj���Y����a��{������$KY���_���[�ވ!)(6Snؚ �g��qv�CQ�J�nN����d�NƮ�߹u'B
����qfg".��8w!^��/�ȵ�P`>zj.j�1<;��.���31z�B��m���)���)�����k`���9e�g�b��@\�c��{��=���2_���搕6 ��	Ս���X�}'���&���숉�R~)�YN�<��W�]Y���u@O��������N���F�7��v�i��2�+���rڙ&�8-=G��*�,@�[���i
�1��	���g��d��{����<.����Mz��Ca��N���n	�X�Ѷ��Wl-ٽ����ի���h�,-I�S �#��,�Q0F� �z�z�S�1,a�d�\�[��� ½ݺ'���Ǘ'$���^c�6�P�W];^rB��M�ƴ�4h���Ǧ��v[�--��JW�z���P�lm�u	�������������I���XY%mh#�� �TI�#;m��y���p%��~�R^�O�������ᡸH���<vy5���%o9��"��a���������k�	���Ʃ*Mܲ��g���2��}=�O�tf�V�b��
E�
_��{<+��Y��ݮ�� `�[~z���qr�J� u��)���8<���Ḋ0�'���@���T5����y��g�~5�A	����1o��m��KҨfOGm��������8���J�ON��W_��W^���s�73��5�BVZP�Ϝ�3�.G���0�ȝ:3�����}��X�jJ�kccQR�#9�~�`���Gy��l�Ze"y�K���W�s���Tx����bwsӇ��ՠ����(B@���\�YNy��r�k�/��l�um-~��O��#uP ��a�"G�}�_?�'M!�����0G=X�qTg�g`G���o��'L�5���9q��IR��?'�(ޢ!�xB����P=d��q������XZY��f[E���@Up����~#��ŗ^z>�����c5[)�����qz�R�9�X��q�#��7���`_�EoG���E��Z���������-b�˪�xd�\�"2��l��nY�-�ӕUc��+>]0f��di9>�uW��%�hi���U��� 3std���m�F
- aM�92�L��`4�x�O{�]�� �9�&�p�ǖa��|S���g �c;4mx�H�C���4gѹ�]��~��칦�+=3����c��u��am	g�l����_��+�yHD�1h��Bް*�������<l$�	ԅ%,������0�/Y�R��ݤ{ EA��������/�+���Oߗ��<��
ς x�IZ�~�ъ�R�z�.���kR4�M��9s�\�	�9���嘒6�7>Ց�8쑶/-��D��� L�2��Fb}��bf��Ǩ�ye$�'��������\�>>��`�轶��Q]d��a�a��^$K�I�J�ץ�P�G�|Kqc��>���=zK�V憆}Z���w��oKF-?�'��&Uů:������	?�-��?�G9�<��(2)׉iN��TJk��k���Ͽ���{e���܉ϱǕ���o��0e��y����c�L�׎�p�G�R�w��X۔ƾW�x�!Z�����݊�^~!^z�Z�뻱�����7����x�Nm�Z�w%��&�&rݤ��T%t=to+�J�g�j����I��w%��R�"/9� �#\<�_�U��r㕶�����y���8�<^����XYP[�9ҏxѯy�eC�3GG.F1�%����2o�+������z����Y�p*����ʘ����3=�Jҿ��2���l�@���˒ޓFXX*����7m�qtoj��J��K���M��IX�IY�%:X�y�J!��8, �����Z�i��)sě�@\2yD&e=1j��lt-y `��n 2�'@ܙ�/��9��CVQq��7����p�����>I
0l�@��;��'M���Jl���Й�q�S��l�G_}���F����{�!���zćC.cdU��އ��z|�hSu�K��rƵ�%�Z>,{J�8{�R���|�LMǊ���5g�!汐Y�o�>xU(<h��f�{��*[�'���+�@�(d���2-��=0ݛ�\���_�>Xy[�׫Qg��C;���@��|��s����X|�ei2��+.�⾴]�����yBz`A��&��4�'-٣���3����8v�+HzʘN���-33�"��cmk��q0}���!�_�������h̜�����cRDI��*zp'��/7��p��5�-AlJCYY^��'+��p!�v[��������I��Ӗ�N+��:�S��6k���l�)9��&<��hJ�	l>sI�۫�AU�N0�y�jࡵ��*)�8V��������z{�@%��e�h>q�
Ӑ�C�� �x]cJy8v3ޓ��ҚG�x���l0oA�"��E�V����q:Y��4 <A_���
C��1\G�8����q�����*� �"I�׿��-[)�O�$.��nJ	�<�C#���ӟwT�ỉ�J/��Z�yF�T1A��&�2�hp�ݲ�'?l�c��_�͘�(�z�]k�.S(!N����p̞>�ﶶw�4���P
��F��W�3
	��3ҧ���'�;?��XU��w�Fs��%[�3��à����i�HPo�~w���y�����b�у���u�rV=��K��|<zj�$f9��_�R̝���Q��:cttԽ�<]�5dʋ��-�"�}��/��}�����hփ��Ҫ{�C�O�}�{Q�"��"eX�mm����7T53��@�);³�7������R�F�ؔ���5��}�+v��_  �}IDATC�b�~�7~�D�I�Y�gSzDpa��5T@��wN�;��J�-^�9�_����
A@c�R��n���az$!ڕ�����/���DC�\2K�`)E�g�����Ua���&���ed
��}��P���)�r:��_J��m&q�r!�$��iD�	�b�WFq��kmM�L&���;�c[�C8~�**Ҧ�grɃ�� ��/-�@08����^���*I9Hj3�Ls�4��:���G��v�F��J�r��'9sd��� $@ۿ���0��XgVJ����pq9|A���ûJg���7`�#��<ӲVU�`�S\�.�ߤ�w�0ģp�W��(c���� � �szn�g�s���I��g��=���5 �z���b��N��.ě_z->��������׼��bH��^M 7={*zz��kމ��zl�>H���>c#�����ѭ��@�է��8�n݈���8d�ֶ4뽽hnl�g���r?"�G�E��܇�~w����黡�Ƨ"�����R<�ݍ��Y��T�Ѯ�EoO����ȧ��c���}ޠ�[&H��YIoH���g�^4��X_�Q�>d�-09��ߨ`�7S��xE��)KJs^�}ܓ�P�̩�}��_�N�m�A9m��IS*
D��Ế����N�/;�_h�M�����'��)��,�w7�(��/M��_�f�A��V�b[-���O�[��o����8w��Z�^	��5O:�z2��TA�.��
�U�C
/mG{����c�LnP����~��6iu3?L��Ʈ_��
�bRplx���ئ��eYd���a,�{v��w�~/�7Uyt��7�
AP^�'�.����O�����Sxrͬ���@=�]~��ƙ�����K�,(8���_6`�l��wv���el��&l,a��X��q׎z$
]�!���r�gĥ�{�8q�����	��l�����+h��C|�'�c��$[�'8�$O�w��#�| ���
�w�2�"?��4E�5,��_;La�A�~�rc?`!�?�R�����;o�'7��8C>:3?�pjã1w�RT��?Y\��ͽؑ�361�C#1*��xx?>{�Ǳy�vl߹�*qn�7jM�
:�Wu�%Ŭ�'��.��|Ȱ�Fss5���4��"t�A(�Q4����^5�R9q�j��+�<����`�3�O+�]���u��g�L�W���e��N]�W��V*�ׁ��zl�AZZZ���i�[^���_�2�\fOKr���`q��C)���u��F%��(�������rC��aJ�2�Y޸v٦�������rIL�/��/2%��4N���q�dL�].�p'�1�Y���%�t�{4��,��\�㏘�*X>���^����*�l �Dڌ����O�{��3
VV�N�X�P~z���OhG�DS�x���(o�2��ØK�t	�
֭6c��PI��J���`�N��5��4�G�p��gy�$
���2�'��2��A��4��@��r`n�]���׊����|8��qX�/hp�_l��B��W��T
z�qY^�/�"�|7�������
 '(��s�x��	S�����\"�%.���#!xo�M�0_)�,h:
C���E�G�.��F�pɓ�FaL'��b�O�-5zVȤ?�IϏ攊�ar�{�����J�g���o�����L|�{�S�{��=�y���U��{R�<Y���G���-��K/�g?y/��(��+/�ű��������klGos'�Z1V�FG��z�ʥ�q���h@�h&�=��oF��(��6T��)Pq�r|��~9f�>K�sM�rahis}=>��#�iG\8w1^|��wK˞;sF�Q���Qw�yQ�2�b�U�=䰐I��7�1: ��}���>�]�����������x�I�������Bae9c����JL���r)d�Yc����������&�U��"�g���8~�8��;.������ɔ�s� �BX
��2<�K�/���sg�iRH	�2*|�����U�����_Z�����Z�H~ƭ��&Y��`Y ����d`�-�<ZK�UH�;�s���b����/�y����}�l���&��%���G��?�A�ƒ�=��F���R,cP'A������s�O��K�73���I6M�F���̛"���#�$���З��"��h���ǂ�?Ip78��� Un'�ߐ+��~�lD�W�f�&��H��>]�`�x�4C�iQ:�QaSK1ʶ�O)��}h0��M�.'d��y_2ҫ����������������O��g��#�/�I:�PW��>�ō���i��Z����+��}��_z��8S�D��r���G��zTۍ�鈁ޮ��3���ƞj���A!��WJ����^첮W���3���W���ވ��X��At��Z�U,�QU�h�bme#FF'��7ߌ+�_S�rƽ7�D5\�H���rF�\��e�d��gɈ�Lo��|2�9�|PYN"���G==����da���/uU.�CY6!��iJ�N�2���=kJ�(e;�*J�\ё;�
J	�L�fx���'ͳq��Z�|)r]�;��s����*(��Tf�Y���t���/�r�LNy?T+�$��F�4�S+���E�qM\���Wo�C^���|F�3��`e�%i�ApxG�� s�zJP'ZB%��ae�w��=�'��K<�?��#	ђ$\�e����z˿|���tʷkغG`�ؿ&��5`���9 �"����kx���=i�1�x�3Ơ��h�+@e������g�_a��g�O���N�������q��P���$HBSOa�=�=E�H�������꾴�{�:Û~�����wמk�G4��}�p�D���1�E���S���F�ǀ�+[UC^�vyzr2���+11:��7o��a��+�����)��)��y�u�񎎎���Pl--���h\���3�C���ӱ��(�ܔ����c4.�?��o<L�x�,.��n=&fbW�n�g�j�1q�L����H^{!:�^���_��_��M�lwUn;���Zx@��wWb|`8z���KK�����Obi�a,-<��woǶ���ǔ_6�B����J�I��Ǽ67�C^�&|��p�0v��;�#���lv�����B<��7��ǽ���=��W_�S�G�8!�Җ��wR���]��ۿ�k�Q��J�{��t�G��4�ur\5Ô��+A��Q�#��K�T#`����FF��O�g����܏�եX�e���!ob�R��$�qf�z�`�E�8�"��cKB��|���<�c2\�%+�1u�$+R���Ƒ)5e�`����j�`<z�o���X\Y�f�Y�r9�����% ڪr��Q�1	�w4��(䆻r���T]a�R�&�|��p�I��	��Gzn�8�#��s��P���ȗ�t����fi���~6��M|9N�e�d�+&	(��P���$��&=O`V��_���5��K���잴G`�5��闵�*�C���Ѧq��@��\c�g��,��|.�9) �3{��װ����D���11>��7nވ�~�<��z/w��U)�̟�����J�<�������p����NL����{q�Χ
��?I �r����1�§�݊u)'}�������j�I��U79�oht<����ًWb����;�cS�Vρ0laq(��C �1{�Њ���jh��z�ɣ�y���ཷbcy!V��w=��V�p��Gdmks+���/�w�G�@]��yQPˎI0��z��>�cG̞JE�����gue%�޾{;����|[�)%t������q�A��\OyvҔ�[+��]�������Ϛ��f�b�/�s�-�
*�³t�����)3~��k��S9��+紖�^�Ԑp��zY�w{ܙ����ע��I%ӕ�*���$}�$?Ӆδ2�WV����#_�Ȉ�I��Et���0Л�N����x����L�ƫG��GL˫��Oޏť���zA��_it�-
��Q��C�\��.�$E��1�&�V����9��)�;���3&���<p����6��3����%�J��e����ޢ�D�TLzN�=ʇ;@S��a)4����cOޙ��Z��f���?�+�r<M��<?J�G ��� �#�;�K��o6�re�'��_Y�/zO�np7[_`�|�WU���f|�k_��v#��gߏO�_��v�S�A	 [�ڠ�j���OO�t���c#�qzvJi䊛�wn��c`�?�ͯǕ���wߎ'Ң'gfcpl"Zݽ�&���;R��D׾�Au�(5�J{���H�a�J�W�8�=�d�َ���X�w����$ ��}3��!M����� ����1�Sz擊{|l���mo�K�N`�U˔d%y���])�_�6Ը���Ng)���	Ǒ�kR�n����Im]�DCl�ة�Sq��E�]�Ͳ\Q��"4��Oq��Ly���"qO�$�/oJP'�2���2�c��h�-�똆�ׄ?��|߿���t�?��d曱�1����	�HZ�`�5�����z�#&����7����G}�� L�`�4��t$*�0'�u���$����g�)A�k|�q�[�����9ne��$�ȒWV-0�������۱����`����L�W���&+Ab(�c��%�|�t�p {y��Q�q�� .
����a�~��1%��.�@�|�ϲ���W��-�K��&��i6h�y8�P�f^�|V��'^��;`�Ҕ��k�FX��
�Y�tJ{�O/@��]�v���w���В��uUǠ�w�]��څ��FK`?�ɛ�����!�w��~�+_�k�/���|�����=y�*-z��Pe,�qv���؈ǌ��7�#�9����Ҥ&���I��;������'�~���O?�H�����w���x��ؓ��Tz�!Z8�����ҭ���풬��Fkg3�kK�%�~��G���~��� 6�}���؝{��Q���殷`�j4=v���NNL�K/���4�͵��UO��ޙ�)ۮ�r���ى͍�cx$9��_s���_]^��v�
��_Q$r/\��]~�@M}��<;���O0���`����KC�g�x�<牠T�����Y�K���P�>zJ���%�93K���p��U��@-&��cjzF ��u�|]��g��)옄��&V[�X�M��a�����l�DK�?9����`�?B�c��`�+���"a\�$ �gA*�	�/�%�y	�����w~���(4 �P~�&�#)+�qL�O����:{���Go��6��=æ��mЀek��=�Χ,��Iy�����HN��#������-B9J {l�vIs6o��<�=/�e/��G�^�� {��@ڼ��=��_��ڲS\V���g��Rf�����0=��2��3�{<�^hq~uO!]|.�g��4�/��瀖��)���3:�~������K���J�@���R��#m��=��(>���+|��l�.�-Ǟ��o@��`�_�.,/�~����[o{����l̜��6wcIq���V�nLj�� =��=i�icWvoi�g�����x��������{���0��Gl�E�U�.��Ź�j`ʯL��]�e��9�n�y�~�,λ'@�z��t���,-1Go��X&~Y)Ø;=;�}rr� Τl�^���j (	�-WE� �Ο�K�.9-�[��z֢��廘����y6��|>�$������{:|ym���ډ�����٪�(�L�T��B�s�=]	�Є^�ƭ[���ߋ�����:���)��:�#�VVZ�ڼy�?'�U^��,��0�3�'��49<�5\�Ni�4��A+�ޭ����G�i�F �Pr�)[��\I	BY.ZNR�ޙIf���(~%�g�TҜ���`%�㗽�|N~
�L�)h��J�8�6�i�/+��3�=�Џ��z�+x�FINZyszM����ں�G�HՕ��z~���
4ȥ||-k`��9a��r(FS�V����B��V�(�d8����4A���F�
�����rl`E9�O���?�(�V$�F��*?N�K�Z-��7bL ��oǻ?}7���T.7�ڢ:/�z0:�H����&���g<������ƣ�'�?���I������9�ӳ�V]|��]���wrl5%;[;ѥ�g���-���n܈��b��g�~�fl=���oE�ޭ�'"V���շ�r�^���WvK�po�-*Y�����U�_e�!C�}��Gccc�ˮW|��3��;/{��7��k˷��[ַ3�N�ֹ�ԫ&�����b)�x�4UȀ����z
h�46(#O���V�r(&�M�?)������zF�u{<>�ߧ���c���D0_���8`��"����Ai��ۭ�뷲��C#^����ދ啥�����r�#�nţJ��$��tg�$�'	��slJ�#���ǽ~
������eaP(�����Ŀ����x���6E*�b�J���q�?�m�CJ`o����!�ǹ-t�>�r>�@�iR��/BOF�2�N��I����G�Ja�w���ѭxN����.2����7a�<p*k���T� �=�V�X{ )�-�p8x��:�BOi��l��s`��j���P��[�Q��W�+�,7���m���{���i?(�za4B�O���@(�r;N���o|-.̝���?�?��?��>�n�Q1|Ի��A'�x)�E.���Ī�_gN�Lƅ�磻Z��cG��ڗ�W_�������K#gE�qp|�[	 ��խ��?������͛�~�N�?�6�$�P��rrN��FDsG�؏�J��On?���F�)�(!4`9Ħfh��ǧ�9���>�G�g�-�k���//1��QXҸ�^��j�V���3�BE:Y�o����v���2*e��UZ����}
؟5e����R����D@˴������CV��ۧ��D+��_=O_4���'��=��ui3���ة��v[�%��w~�w�$Z���{7����Ƹ�O������y,���9;v��o��)��ϏM��y?ݐ��q�Fy���
WR �����FL�6������?�ݦ�m:�ʳ�H���#�{ҏ8ӗ�z����4�.��@�3*	ę���K���� ��ı1P	|��?�� )��b��2�i��l=�x'�����(�F��Iv�)��$��պF�$�������Uio��Z���c�\�}N(���������"���2�%�,5"�!?k����s����r���?\�\t�'�h$d�aH]+N�9��zN�y��zޗKq�����W�����ͯ-j�=����^,�,�\����Ucg(~�`���KF�`N���ӳѐ�l�p��"<�5sa,�ewV��W�>Z����c�����𓈅�8\Y�X��\�!��ڋ��ztq^�aK������99M�ʽkly./�iB�e�aV���{���)�Ǫ�	i��3���0���y:�X-�i!kf��/�*�x����;l���a��OFڗ����	�.Gb��ۿ|����u\�E.���Ni='S�c���ϊ�4<�8e�$�pU�W����*�q������,8�0��Kx�QM%�Tc�ތյo����}wY�6	<��������1:>S���0��*̖��nfCi�I�c��d8h��c?ZӨ��b"~�8�鶦�J	�-4L��z�� gdt4����/�����ţ�e�*�E�EP�<���otO~�t�k�V%MaU��?���Ե)/�*F�v��Ж�EJ�ZEa=�.<s\�!aݥ��)pK<N�Kh���8e�g[�c�7�k�R�xF\h����d�8���_<>ص�IJ�mx_<��)�|�P�7J��[��2@se��Y��#?��q]N� ,�m�$��	:4e&	�O���'��~ɛݼ��[�;o�@Z`^�3_��eȓ�'^��`?h�z��oJc?h7�G?�^,//y�J�9J���Ɗ|�i�CO�*�~�h���sg�����P������n��O?���^������Ř��8V����Jl�/IWoC)�Ҧ�=l8��@@�0 .͜c�\��O��豄���|�>yWJ���s3��[<O�/s@c��1%���亢�ܧ����onlZ�B������=��/L������Oٗ�N�F&����-Hÿz����1�|yMZ'l����2l�+��J�I7�?�ʛ����9���ɸr<��x�4��Q�EX3V��������,��<W�W�۷�׽-��N#����㳻������[���Ͽ��A��VZI�<��3�J#���%���t�������/+��p�����B����@h��E��a���_���xi5Z,����a#��_��Ll�P�D����E���l��*���d����9M�KY����(YF���X�c+ޡe׷x�ʖ�
�8�"^�[\'����(9��5R��򧪻�4�r�C����/j#c�S�����Z8�qd��U��_�����P�MM=�4ui��	�ZK���Z�"��o"Z[G�iܻYnk� �l���;��<'��_���F��u�-�4�������ZSW޹ד+�<�7v�c��ꍿ�߾���GjЛ��F�������ш�).V�0C���h��;�奥Xx�$�jĶvc�mw�`ܭ+�=�ٓkW ��f���Q��(��'�mlGǁ��KdK�˪�#.��h�X�[d��G��d%]�R��8�0�y��F/y�P���hLM3��t\,Űbn�V��W>"*e;e֤�l=��6 c��};��w��û�8}�L\�vմ���:�x��Y{R6
�3��O^�,�?k���Mq�B80%}�����'����22_*5]g_*5�un޹#�n`n��.S���	�9shg~9V���dqE�]�M���ZL
�)Qvxp�]�W)��	^�G��c*�e<'��y���*ʃ�W�b^ǿ���3�?ZX���a����VXµ� {	�^6g{�>����ɽ��r����J~4Ee�vԂe���'��OYi�T���[ <�oR8�w����+b����%���~τ)-�y�D����m��o����'bhbғw���F������h5�KӴv*z�Cs'.��{@<A]�� 慟�u]+����^��-���C\@�]��� ���?ܴ�k�y�O�D5Ps��6������lK+��ވ��qi���ߋG�z�h��g ˏ����S�'�> c�T�����d�u���z�?xh���M�����
'Ab�U��.�P��P
�┬Q{YeRi���C�c�GyL#Da�u[0#���L�����;��X��\D��ˑ���wz��Z�x(.�Kxohx�ߎlmm{%r�x�P �����i,��裏��g���t����k�_3�;�+��H����$�c1������!�|��й6|�72����-��-�9�(�`�1Y��=N���--l,��(Y�A'�%���V�aM����1���Vv�2~@��+�Ǧ�����:�Ï������ǟ������ʯ�lBN:a�JRȖ�����H�B pO?���4��I���%�[���~��}�ъ>�����g���'�P�5t&�8��:B#I`_t0d�TOXi�`��-,<�%k�&[��=C�X��t� Ґ�̏/ |�a�@�2�Ol�2W�=lr�9���?���)?ݥ�(V�Fh�7dE =45�S��Tw�20�Z�g���/����֭<�Cj��w �1�C��<�@�$�Ȯ�� r��I{�ʑY�G@ݚ���=�},W�'��r;��/��N�t�t��{NJ^�z&��l
l���-�2k�K��"eAZ<C1$�,�e�E�1��B�NɊ���m:-�Ex�oV^j:�]z��P\|�VC==�%[m��QI��P8���`nUE���;��%8�
H.��%�L�g|����R��_���	����>6�	T�asj���mK� �ML�g����+��2��4667bue����q���E/(iJ�S�r�\y.�<wY���GEY+X��}q�d�{����1%����y�:#�H1e�V�_!,q~���9nҔaO���?k�=~Bh
��`���4�O��+�ٝ�����0�4øԸX�֯����?���?�J�au��g�ܤ;լ�"Z�p�
̓�&7��8�ҷƦt�������CӢ�+/�����?��߈�n܊�����.U�������J?2k��m��l�,Z*@εߑ��*G����ށ!��1s<�)�Q(�aV�X .Ue�\��c������J[��^vU�����5�'m��*N8�P4�Q��t��G���/@���E��<�����@��su�ާAU�rK-�
����T��*f����e,�� ��k�ј���s�B�I&d���ʼ).L�z�eL��Fa���.|/,�揞�%�F�������I�%��.���F����d˨S"O��KPC�]�$* 8�,��t%˩G�[\qN	�?�C.�YR�)����Un��r)l���/�!�k ��x�_l+mvF��[偉]��E����Dwvv�G�)�l��>�S��!����i/��X=峼��Ӗ���i�w���`���w&m�\ܽ{/�,�&r"�\�fK�+W��������@��\ʷ�g2?s���2��yM�eB�X^C��等,×��&ox^j�G��y_���s���be;θ�G�T0��=�������D]B�L��b��=EQ�,��͏�U T���XR���ߋOoފ'�q��y��r4Y�0��
T
d�dQ8�G��X(�	��N��n3��������o�ο�?��[���k��>�#	�r�e�F&�_����o�{f�E�_��/a��;�#�7:,�J��y�qd�]�G�4�
ڭh��#i6x���*A�Oy��:58�k�I�@.QiN� l6���Q�-'?��<S��[�\��k�� v�l�������G=1z����W�x uO��%?~ �s����PP���Io9w�yнE�|G���x�Vu�cҺ&��+)|RX��)�C�S��Hr�����P�.����˖��>%��>5�Cn�
T�����u{c=����3r��tH�4�>����a�l���<\']�'Z����;eq]G j��:��◗�]�������lDiJ���'v`�B5���8����=�v�� ��?��b����֛�MI#�?�������tc�?�/�d>�~=�W7U/��)�C;��F������T�#�����x��r����N���W�|�h�n�h,��+{��쳟���9���ѽ�(�g�x6�q������ rEZ'�'�d_�Ӂ �M�m*���C�MJ�ތ��u�X-t���PQI<$c�`���D���K@�S7��yk'�̬�x�B(6�_��*	K�(ĤY�S\#`��Ig��#�՟����a�)�����I|�Go�?�����o���<�~�#i�kҜ�ct�T���b\��bl�5�]WlG�{`$�k�у�;���,{n`{��Wx���I<�9커�rj|ml2'+}�Q�h�mQ��)~x��F���-�I^vlj����w��Z|��ؼ�����k��BK:X@@|��ON{����F������hh
��C�>A�AQq V�ec����`n���ui3��EXn,�_P< g$Yw���yx%S�:�E#��G��ڶ��g��_�a �x ��W�!H1�#<懆E��L�p�P~���޴o�wN;��.p��0UEN*���~1w�܂�Q=�çN��
pw��	\�k{�?"Y5� /�4DX�<ҋv/Giv���QY3���aYjG�h�Y�����9���C��=7"�!�c���'�E�hF���8�@�KW�=!{�yu�5_��| YN��S �Ϟ=��g/�@��;w.�����=ˆ�rO��"�D��q[\w|��w���BhaO�=k��/����Y�sl�iR�|>n�+.e�˕ᬱ�^a�eJ��|
����{P�Yoy��nu}�ZR-b�y���?��
�ۇ�>�� �,xf��Q_�����㗾��1��^l�=�Sӣ����h5��8wj2~���cvt8 >hFǾ
Db	u��8�x2c���5����Z1,�������;��4j5U	;R�VWmsk;��6E�vT����/G�4#�B"9TeR���L0C�d؁�\i���J@����Н_��J�=6z(��6�����Z����h쨡lʯ�'�i�� f���\�*/`Y���h����p����ʔ(e�i�ȈO6��2aȼA��!T�ā����m=K �4褕�h�A=J_��
k�-��c�:w�r~�I�"�ă����Kw��d�ܰ$����heh��i)�)7��x�K+���AdQ�$L^q�����"r,���/�I��g�`t;��w��F��Y�h�Z^���M1���j��$��d��������<���h �=
B:�$��oo�����N�x���C>3�βS�RVq�dY�@�C���#~>b��Fx]������e�Y��N�V��HO~ux�z��)́JwI�co�矻/?�2���
��%�N~�F�±{m���Gō>�ڐ%�U�˳:�_��ߌ��z�/����d������o�����W��ˣ1 a��/JM�O�/d���_����-D��I���/�1����H狞=e�8�⺸82J1�?��qK�^�� ɣ�V���!I�@�o�=�'��[���������k����]�;;'P_�0�cfj"��$��3gf���^�k�]��h!E�\��%��C0#D����MA������.������٭���Qll��QY��	�;{�=���K��J3���hu�G�#�R��������B�F��/���Va�+i��͉غ�[ݖ@�)�jH����K�)MB�
k�aeFѤ�HN�8	e~�SU�=ZA�����qc�����zO��*�s�(�ja�����f�
�{?е��'CK�����E�,�J=����X��F������TюE� Cڻ@F��)]g����Q�K�����6��z�ґ���h,\u\/$���m)9����
ڿ�IIW>[Gk%+DF����q ���u�ȩ#6�"ýj(�ʸ���\� 
�� �h�|���&���zz��53�,`�� ��y)���@(>�i��$�.��tA�ę���r7˒o�:��9�����cpB�1�s��D�IY�29:}�a2��'[�����٘�t9��]���SQ�플�$�����[���)����+U�@<�M9@%2/��/a8��vzRl��X�Nn��E���YM�GG�A�mll���u�y䁯NY�X?��M�JS�4%��Zny��ɗ�5�߳a1�.��|.�g#������� ���L� �}�	���8�ƍLL���H��_V�z�>�jmm��z��"t��mq� �*w��Kȇ�j��4��J�����^���i؁�̧���@ ؂*�#G�O���<�9ݿ��?�{���4vU����4I�H��R;XXi�]�QW%���=�:Z�]*ַw{�!��m����ϲ�úxlK��Һ m \��C(SRp��$��5K���'���K��(����"[��	lmkC^]ӧ���<Tk,9=��%�C�+�}͊��۫������܉w`�q�2��+��a�W��ɐ�]+J� ~�|��#K��S`���HM*ZN@Kc�s�@�T~=�{�50H /��<k��r=���9���S�H*9��iW$K��i+��|OF����z�O�����)�U���u�P��]��b�$�٫�G�S/ht�d�!>�����$��S�� 0�r�	�P����A��9�� �F͑�`�}_�`�i�J)`�ʻ22C3gbd�LT�&b�̙��pQ�}*j3	���18uJ�NG��fO���sѫ��o|5ν��O>w5�.\�n�{�eXV�L�����X��h�Ih���t�L�F�V~�@�����vw<D�{�1��·Jo��F����\�����M[���1�$.^�W�\���t��,?�+�e\��mu�3��N�����p�����$�X�+a2\
�����oFኡ?m?��?�fW��d��i��c}s3�����'ާ�gT�gc}#����W�����F��	H���*��è���>�K159�]:Ν������	-b�6] yD���х��v�<ߺ{?~�w�� ���^��`c��Y�M@*�eb�1t���*��� K� w���)�>�{��m���m��@��k��L�h��(�GdB����pќ \��olx�'�|�34<�#jTG�&���i�M� ��a�������<�OOE�`�\6nc,����Za�p��vU�92!
O������|����Cl4T�Wnʋ�^�r��I�N��Ǥ�"mȨӰ��qo�-��y�g0V%/+$r�FC#a]����Di1Y\��W�?��9=��U�
�0���y�2��p:���d�ٚ���[����������0�Jw�Qf�`G���-�Q ;�}���ۧ�z�h���и(q��}��oKcߑ2�T�bn�~<��#�\t�L)/ ��y�i�۪|�箾W_{3&�^��ə��HC�6ޡz2��N���K�f;�ۣ�S�f_���f���dN����1{�R̞cO��xp�����@�_G��ڥ��`��G�2�f~~��1_���mE�L�0�A��E+o/xI�]}�W�kkk��w��e/y�9����S��L�4G�p��iUL��Kbym���M�
�D��]�#-,>��y\��E����㊦?�1
�Pf�	�T ]9NZ�Oo܈��}�?�$��������`9WcwK��o6��|��P!��6���}��\���"��K��4�>\���h�1���̯"�_9��doܼ����ح7=޾�!z��hH���������>6%;������[J�84	 >Wf('3�W�5͕R��E+MN*,��,�z8=W�k�!�sqB��F��R8xO#����\l�ea��b�J��#섛=��Z�3�Y����+�h��ӫ({����!��F��������2�0Y�<@��1*��5��Z��5dK���76���Ô�vn)�#6�Ǖ^�`��-�S�*
��9@Z(=�G�|�L#- !�"�
��:B^�J���<�Ki���n�_w�$_����G� ��ue@�V��P	�
�]�����E�4;�gG���{��`Wy������mU%�+]W�ڱ����u�l��a�vȄgͫ� ���qi�}�R����6�aH�T_TȔ�n�@ݽ�Y���Xk^�RWU���ۡ��n)ջm�צї�@�PCyN�z��ה׊���S�5 �h0�d��rO��M^F4u7�T$��>t��3�u�ndD=I��������X�_�Ǐ{GQYF^~�e� ��c����2��M��Fj���$c��~Ϛ�*~�sw� �2*b����w���5n	X[��O0(��ۻ�
�r%��7�0&r�HE._���},��ǝ�7b�#���ң��4��T�;�ާ��c?��Cծ�떖!���ߑ nH�،����\�����hG̝9��t�f��N�Ce��KW$Y�ܮ"V�]ռ���چ$V�$�Pi�J� G�����+@K-"�y�b����ƥ�����eݩ�_�ǁ@��`[O���V�Æ�,���4�w���O4z&j��n>��W��ӵ�d�_�-�Z���ai!c��8l}���o� �T/ w�����D���}�9�{���������܉K�K@W%V�r	BF��%1&�����;a�+�a��c�T#A�-���=�]�H�E.��8T
֤�эlS
G]�~ǕS�34��&I��ch�XL�m�rC��_Se�'�.�dWB+1h�/���hF�Ik	��ߧ��}��C=�ʷ���ֺ�^.J/���v~��Sc����&��醨��ʈoK,�c�U*��M�� {1.��F�������h�W����vW촑����؋��_�O��I���������/ے3�{s��;�u�B�Ta`7����$hͤDQ�A��E������^�����Z��E���&��&� �\w�;9���9�����;�ٙ7o��Ŷ�8�fĎ�o<�F�ر��݋��>�,
ϡ��ݾ����;��u�q�뻽1{��x��W���?q!6��c��/Dq �1Yw*��,�IX� @῟�ӥpjN3��^x���?>m����������Ř�`x��Z<�/���:j�*��'��`���O��S��M
!��X���}U
�K&��CNl����n�񪿿H�Qb���d^,ؐ�.--��Z�R,�,�;� ?R�����qO#"G���eM�RSߌ����W�ƎF��ٸ4tN��ooĶ���*�k5��ؖ��祥������阛)��U��Hvq���zQ{�j���.		5����7ߊ���W��k�}�W���RB�b5œ�>}�psZ�(�X�u�C)��4���d�����T	e���\���.��5{jU�{����=�� ��ǇR��^Y?J\ڷdM�9̉"�c[������-�#�s�0��`��Ql�F�ê�� �dI ����r���Ĺ���c�=��b�D�<�1��$�t2O՝+�J��Ԇ�2I��'��D��x��ys[�Ê�}�y��y Py=�+S��Q��5~@Qe�Ҡp��Me�;r�ь2�<�ЀK}Hʤ8
����[lud�D2�rM,��L�r�O����UY��־����gS���i�m�օ9�(�����Y(Olv��K��[R�N���W>C�NHc?�Cc�s[+�ݩ��+�^)+w�Ń��4��G�G���A��n�Ŭ�qi�|�G��M�|Э����b)|K���~��_��6�v����Ad�;kTc��wng��q�<��/~�soyD�̓���Ϝ;+p�u�\�x1~��_ă��{`ë����{�铮��UvYs7QdM� �� �݇����PML�����k����hX����
\Y]邷���.���<ey��q�?~�(��c3�E�=z�1�a}�|��������:̶�!��2�k����������c�qbv����5	$B�Pxi<[뱦�6U^�~��W���\���B
~�	�il�C�;���U}O�%L��n���K+��?�~�譻�����[�` �H��?����l��ߒ��N4Q	-}����H �$O���1�
c뚎X���
��*�s�ᬱ�W���-p=��O���ܻ�#)n�u^!n�5X�M�\�@WeVI�<�h����+D izUH�2,�t-�f�G~�9s��;9q�v�<�PH�%���i��;��܉ӉG�8��>Y]�2b�ۤ� ���nnZ��M�=������t���֩���$�b�-�m)Q��V[�&,�.�p�A+8���G.�%W�O������F�0�kR�.(��;z���K�=��������q�liַ"P_R�*ۀ)$Kkjw�ePs��G�f��4z�dL��#'x�y.�f���n0SU\�o?{Q�]�L�߼{׮�bU�%!�35'���@���ǈ�}p��(��	^��-˞;ro�ſ�1%1;�=j�()ɕt���nrf2y��Q���X��ʊ��m�,������x�;�
��\�.�~�-c"a_z�%��{���O�[3	됍<����?���G�����QƝ�Q9�%��%
b�z~ޚ���nO%t����5O�9��y*.���ӎ� �6Ȁ��ԅe ��S���?>��Ek%���{��>������b]���چ���id~��g���s1!���F,���,Aڿ�|qiY�vSy+/��?����x��3͛1�@����j}j~�3}ԭ4��,3��"@��;����w�g��u��j�BN�m�>TN	�ɋWb��314}R�>f�(/���f�t.�����<Ӯ�e�l��w^� ���F>BiX��y�C�-u��nJRi�����r.mK(�"%�,�=���x����1ĩ���XW!���~OR������#˓��!�HՑg�G�1�+C�J���tX�͕�5b�� 
���D������^�I�R0������(_����%�Uj~��wT6o���1�b�8�O�M��°���̘�U+%tf<��\��wcki1�F#� xՅ�yp��+r�?8��/����k<66�m.K[����GR��@mZ�����.�e2xƻ�3�����>s�r4�ƥ�O�{�m�q���5�Qg4�=���Wߏ��~��HS)N�8s1F�</��W�_�\Q>����[k�5
�V�`
���D�wL}���G1��V�h�����k��4�:�I�� ����XJ$Z;+�?���[�EG��	�W������}t�x�����u�:uRi�ݪ~����G��L7߮�������/��q�:�Dy��"<��{�W5����v߸q#n~���FۛҺ�ܽ�5%�wOӪ���r��k��3,�}EZ�� �/�����:�����F{��ei'�A��}?,�b9Gip�{���xFS�Q^B�,	���X�Lb{C�Fj�A�V�ӿ���s1ڿ����"՛�,2�ε�@��jV1��?�o�R �������(��z� IZ�ԉ�125{���A`-��s�El���Ӏ�L'�@��������u��*7�o���`�x���s�����������m��'�{ ��A:��T�n-�"Qn��VЮ��Vav��놲y�B�r�+7|���Ȏ�_u};�2ʷ��&
�]���G?r:2e�qB�)�����������o�k�D	2P�W�@���ui��
�v����.�{99�YJ��wzUJ[�=�Ӿjsoc���Рʡ{<�#I^ē���i/m+`�p������?�2�z=`���l��7@:(d̎x��K|n���PxX�˒��>�9�)zt���>)_�k��<����Mj|�l�Ϟ���hlKCo 묍SZ�ה:�8���������5:,-]i]y..HS?���1xL�ڠ����������m��ޡ�a͚�u�_u��9��;�Ⱦģ��rp�ԩX~ܓr�}�r�����e/���뚱���re�����u�������(*W�{jYd�N��-�Q����C����Y:�؟ؔ���Z\\�:������;�n�a9eeu��;���� �wLK8.�}�$�樆P#�#��*ʘZ���� ���	�y�5?���k�-�s)] �:17Ϝ?k��ubi(#Ҟneq^�� �U���������P �L�4���f�KI��d�O��M�Cã�1��o����;׼=@��u�^M��I&&�o���|��$퍇���#�����*/��<�����}����Gtr
�v�}/��䃮�]�4�]���<`��{�ul� �=/ǈ�K�^�/ըmP`�!�����m�~�n���z �z3T�����jv&ǥ�;��Y��,��gRZ�|�"dCzIyrZ�	�x؅0�!/�-iqG���PNy��n��oJ��ĳ>i�����k�~�E�;0��ڔ�*w���X���yߊ�E_߬t���}�N����C��G,�DU�>��e�9���;q��q�V��c���^��?�g�O
�gԯF��@z$?�XXa4X���b �QQQZ���Z̞����D�����CK^�l��<?�~�N=Nܑ202�B��f�'��L\�ϝ����7��ܚ�m�x���Κ9���u��3$,c�|����j7>��Jr��~��d�#S�ϠQe��[�gΞ�%�_��׌��$c���fto��y�u����!�)w��,�L�^1`�����~��'pT&���4����ү^���7��۬щ�;�~ּ�4Jy�F��S]�w f)�Ni�P~ݲ�{���ǯ�\1@�5n�u
p r���g��=����܌:U_l���m�}�S���%J�Wq��������4;Q�e��(�>�eMN��OLL���j��o��}w!��F%bꚃ���'��e�W//ٌ
���c�O�-�K��<�|Ά����&�粎��:ë��L���zr ����u��V�;7J>
p�u�|/�ؿ,��D� �d޻̩] � ��\.�m��W�?l�sO�nՙ{rgl���G��v��VX:'�E�����,?���"~q+/��-C{����<h����|b F�rW{���o4����!�tg���!��<���|�Hy�U�A���JZ�:�ۭOm;JlC����֖��Tc�i�壤��%YP��r��E���n9lx���{��11�����Вk�(:�������36����d�Pl�ͮ*º����EY�Щ�A�׀�+���-NN��ʴ)�����4�u0t+�rS��`Hm��0/zۢ��G�ɏ���!�i����x��X��P�����{�N�k��֠�' �4�`�ơ�/��R���_ǥ˗�zq���x(e�U����ߵXqE�H��O����������w4v:�Q��Ŕ�����d&�3"�\r�������w��5У�{�R���M�v@n(�@0�dg�)�D�Q�����W/{�`�@�'X�2�t�m���:��Sإ{ 4	bo޸�����ywH!Q|��7�o��3��rEڑFt%�)r~�O��u�|��Z:�~H#������x��oǽ���`�=��|[sO��G�O�:/%��t�� �«n	�t�bg}�C)�n�ذ͵���r[�Fr;�P	�	>
찤�S�h�Qn��@%O�9�6y��"7�
S�x*�O^�C�Z{9~��q؎�o�:��&�gd�i;�Ξ�Q�.;�P�I���>�t�i��~��A1���	?�t��.��`�?���С�*-�C�O�bԏDi�.���	��Bs��W{�X׬��,@��ཹ}��`>3$eC¼��N,ܻ#*�Z@|zr"&�xlnlz9>3S�� ��o���v^�����4���%)N�JC�wS���s��T\~�����[10s:ޓ����[��?���JP�K �z�43+�cP�pv5�YA�����V�/-���B,=~���T޶��y=}�&�P��9�zwu)�?����c���ؾ7����Σ����(���cX��1
S�ӳ�!?�ԡ�3F[n+<�d�H�K�u�G}�C���7�!,��i�|r��8|���p��W��sp�%L�M�E�H��0����������q<��i&;e�L�� ����۩5���GD$Mi&��(�;�9��^p������4�|���X�̒�ʀ�Lɋ]�1����b$�Π����A�]:ۛ(�:Ϥ��vLkj���>��_��ě���0�W�'��AY����n�����$�������o٩~{  �\8cpB���G�_P"m�WQ]6��UeU�F #��Ft����c�����b���6`m`���]��3ӫk��Xt
�ˤ�ķ�k��}�Yсr�B���8"Z��6)�r����K<L������t]V�N����W:	~�Û��w��5i�NgǸ�Gh��*�VD��%�#I��	� D.G���;,[Jaّ���]��Ɨ��wH�R�Q6֖cC3���e�j�����ʱ�ǦF�>�ٸx���hǛ��J%��0���*��,�ܞ��L�}��@06:#ý���bfb8�6Wb����{��S��R\����ވ�Ͷ���P2�E,�*�Ae�2[� L{UֽwT���˷oŪ��m�?��%�Q7bcE�f��l��cJ���kwnźh�������-E��gu1z�û⓮g�{bN��o��ϒ*�e�P�SNe���xM�MNL?6���̥g4`��<|Pk�)��d<R�w�[���d&glN��J��ם�A����{H"�E�TPd���7���w"�O(SA}-7��[Y|�OT���h��k�"�a��KЗ��ArJ�V�RLj��	9���M���̦�����j� ,���K0��D9�FF��0;wv�(�]�͋7���0�M�,�#�&Z��.*��)lC�V���w�������:oI�{*'SH�;S[��U'@S�������?kҕ���h��6�v�K)�� s嗚vR�Q\���$���L������F��&,e���%�jP@��:g�a� 8u��$��S�a�\\���v�?-����Ȥ�M��~�¦!�=�ٹx$���P�H3�U�T����[��j2�뢤0��� q_��ov�h+1����N}�>�x*��G��H3֗��--|w}=v�p�C>�<&��t��)��wt�m������a��>�)Jg�-:r�ܿ��� ���ߎyʹ�]�n`��a³'0��P'׸�#����o�ڇ�ᎍ��S��~I{ܸ���Ђ�&�mx<�^z>�\z!�<Z�����Ku�A.���b��Ѐ��%#!y�̣G ;�.5�ڊ��*�n߈ޭ�ؿ�AHU�f���,���܈�[�cx�7�?}"��c���"��cD3�Ii��=혓f>�ۖ���=j��E�ql�7Fy���َ��gL�|�f�`޶�2�7���z���f��d���7�T�l���������`6��٢m�V(H3�A0�SGc��i�X3�5�B�CUP���Q>`g�C�V���f��>�+ ���� �1x���8~�xLh�W�899�-@���� ���Zy}�rr6~�C|�p�mf  B�4�2 ��3# >��˷X].�����ഴ��`�5�[��<�׌C���@��%�Y��L�_��@��$�����+��x������ڦ"��k�*Ϟ�pn�.���Ǧ�/#����Cx;�#�]>	:�耱�`��޾.@�{��E�����.�a�5qW�L��`'�D�F�U�����w��Ф���[��"۾VrX�$q/�3��Ɖ;�;\-LG~7����A����%�Ku�0�}�->v�&����̦FN_#Kal�U����U��8���;���i�>'}M�ŬJ�~�!p�U�#ʃe	��/I�W�x��R�H�y��U��# ���'^y�eϰ�~��h�v���(�?π)gU���[W�ق`	g����g�����W���wbE@��{o{�1lKD�=�\�;��+�v�U�Mi����ݛ�qG$w�4n�g���6�2�_���X�}=����~xG����Y�� *�dx%����s�QkS<�����I+_�Wϟ��^<�F����n��ǌ�'5ø|�D<{�T����a����ր�ґ����1 +����F����n��cn�e��W��Uc�;g���������j���Ӈ���܇���b:v :�|G�]		�ܛ޲HEXGb���K����ޟ9!�F#8���K�T٩�)k�<�Xv��H� a��O �'���x
����ۅ4��-�zهBypx_ G[�YT��|p�֦��'�ªߛ��E,�/�Gu��W�O ?*mekA�6��}�y��	�)MgB3���b��w����?����G��}Dњ:"�O40��2>sL�̘:StftF��Ѱsm���m����� ��D%�? `G���V�nЭ ߄L`w�4�~E� @
�VF �C�
�2.�Gɑ�ͮU���:�p`�UzY�ȋ��yM�Y�AE���^�s�_j����U��GǫHq���n���u�|�4B��� uZ^m"�SC#e"@9$=
�n7�ϰ���@kC7���4�M!K.�T6���3/�y�N��}��K��1;V��� �{��Aܼ}�{�����C�/��R.����`i����+/�?�{�Y�Rz����މ��5�g�<W�}A�6�n܌�Wߋu��p{=Fۛ1�\���mi�;��7��֬z��R_�l`O�^~p'�_{/Z�o*�fJ�TO��{,i�������]C[`ޔf<�؊�~��x���x��LL)��k�x953�?��������p�,>��^$�O����N+Ss�'�n����?��O�4^��kƥ�ׯ���{w������ލ�Kk?�� �����w0�Cy��س�?���+��" E�>MF!4q���'3oid*x#P�#����j���҄��MT��ʦ6͒�ˌ��$@�1X��:�;vlN��~����#�� ��c�3��>����JP~�1 ;����Sf:/;��A����M	��7b�ƭm�cDeg�	�x{iY���4�f���������7��_BRe��"��p :��og�h
6:�8w��������^��־��	(��\/�%��m�)�2�⣑�f=�k�����T�G� ���i�o��t�J�"d��nw�#	�6&��E~�J�Zp��_����Hit#�"ηx�_� О���f��A3␧y�=�eB�[����E<�˥3�Q}`� @w���$��ڈy۞����8k���C�|��[��|�e#>���Y�d�ҐK�^��V��보����^�N�*K*7?��Vԝz�|]"��;�����8)�kD
֣�o�����=>���+����Ǥ0�o-Gk#�Fzc����q||8zw���}lr,fQ��ce�QܽqՀ/h�ۋ���m����&��+<�������9:�O��	�571���eܿy-���⫿������
���ZlJI���]��JJFE���R��1�~kX�իW���Tw�_J$/@��A\�y;������5<)!�,�#iQ�
yV��;�~ؔBah0�S71�r)@���ζ@}nnNڹ�W��a�삡t����>�{9�HZi�,�a`*���$��^^6P���|�Pǟ�*���1&������y�cS�X����T�t9kP/���F��766u-MR?��;��፶�'M}��B����Z]��'�<ܽkw���1#-}K�O���������͛���dGi���5�;�Λ���g�F'��>?�϶���|Re��2�·h	渱�S��K�pS��/� �^��|U��`8�� ����M���h\[ �k]��L?l���kk��T"]��Ґ���^��{��=���[���kWc7t:�L-�z�����5:3>��,�j?G����+`�#�q�e���@,���Y_��a	HY�t)S)/�gF ��i������֖�r��y����1CB	�(��h\�������Oڪ華ť�������۟6��DY:u���@��e���2iƎ&��+/{���ØW�㝍m%3a���^���ڗ�_z{k)��xkCJώf��C}{156�R��9��>���?�����Z�����B�(�J��#����a�̙�9u"T���Q���;ų�/�����v?~2����w���XP�_��x[��N�S��5�ڐ0V�P1v+�"����em٘u���4������fXK'�yx<k<&�SI�0𹓾����W��J�	�$�kF��]�T.9�� 4]k��ҧgg�������'�Y� ;[:��<A�S��������I��� ⴪��ƝO�T���t��m�EO�"L	��F-��m��Z<Z��6? <Ѱ�w�T�����S^g��0p���ݸq���x����������wގ{����gK,U��ҋ����K�mc<4�#�=�/.���)��j��F��1�k�O���|���\c/�(�>ԣrwl:��ԋ���/9�����l�<Jq�V�����h����9�0ܳ��m�aqk`ŭ�K[�T��] �?��k�U폝�U�Ly�g4�����e�H���{��=���[�B � I�U�ސ���hFH�yF������!"������F�(�0�kcq>��@���Ν"�a��G4�(��I���(N��N�۞����^�/�������+�e��T������v<Ҭ��2�8y��r�._(�R�x�B\�x6.���K�OH���K��F�J��p攀���p��T���6b�ѣX���VN���a&���Ƭ��9��H�S�q����_�zh8�����^����b2���{�ʫ������O���J���;�C���V�q}Ɇ<J/0;�I�`�����o���Cp�
�����~��*d�I�A`J���	�W=}�iGe!Ç��^P�E些I�&8��ۣ�� �S��^�ίǨ�H���̜.G<CGw�RzR���3�v�����,"���ٳg����/�4x�#�S��*���w��y~����7�p��<ɟnL�#/+�T6������*����e�q��n���v���xGS�^i[ҿ?ZY���Oo_��r���y@Pz�zGiw@]���T�>Z�31}�t�M�)����~�UB���h�h�<8e��
�{h� 4�Ծs!r@��F�*�%U��r�K8���X�C˴mw��]yH` �}��4@��2leC�^�ƶ�
�g^���!��a�5��\���r���Y���(�ĳ:����/�Y�^�㷟Q�8��%�٣��y(=+%r�c��D�v�N����{����8Fxp�S��艒�]�mU&��<�&ΪȀdCwqSL����J�)�m)��iJ��/2���*Ͼz��R36$?~,���u/]��g.]T�v,/>�L��-ፕ%XǤ����߉�������Ĺ�[z��\��,��a)j}5v���D)b_`�~����(�ELL���+�/������_���x�YX��n܊mu���/�����w��/�S'�ĉKWbwb*�C#�0�ܔ�y��J@+F���[�#�����9ؐn��ߺu��6���<?+�T]x���n���O�r�T`�zd�Q�)�h� +@
�Ra�^ؚ�S�ʮ���"^��}�� �0l�a����-�-`�H����N�>/���w��M�B��Õ^��k|,˰]k���.z&�B��n��Y��uy�ruo�A� �hA,Ѡ@UOk�I����^��$p[�mEZ�����źz���[U.N���B>�N<�PHxY����㚅�8CcS�֥��^�ω�戶�ڡ m.�\�a`�KK�K� $�l,)IX�q�e�qG-aX�OW
S�Z:B�zX��ۯ�랁Bq���!� PN#�c?���]� ���ć8�{vw����ΰ��!��f�ZrQ�3 '���y߁N�,�Ά���<�!�9Q�*x�t���p�� ��滄��|nxj[����L`���5lrzm�g�H�(/��i���S��g���Ay]�Rf.V��g��$dC��L�q�ŀ�m�𠕗��w�dȁ|�����A�H��,��49�c[��8%���oY�Ôf�Sִ����N;� v�O�_7Tv	���=�]α��t>Ē�L��L<��߉Ko|!�Jw]ᚚoi���^*������+���ً1s�b;����;6�~�2h#VcC��?˗l�G��|)W��������|w|B�oX�H|S	ߘ� W礴��� �k&���Y�`�!�6���r�ӽ��I��y�2 �ƺI��Gt
�dP.76��jl������h���{����1�t Q"���^}�5�(ĞO4{��u�Dg`�̣�1�A���t
�=��'O��ii��D0�77�P�N$�.�:���a@C�		���uA�~���T��:[S~�R9�����8- ��crSk�)t[��2����N���i�����]|fP��؅�]��-~쬉�-�,�`��1��f��p����t�m.�h )�J� ��v�9A�h���5p����J�p�Ja�]ܵ�	��M`�Ӷb��]�Jx�Ӑ�+�7r�ڻ��|� h��Z���3ño8?fa%@r�t�/�凣�~uH��ǜ`j��<��*����|a�����p
/��-Y�ړB�+-��XF��ب2�.j�s�x+>/���0�'�
C=���gLU{#+(0~�D+��"���,������(x�KaQ��r ��0���|�O���|�l�L(��_��='��2$��,�/�g�|&�����������������?�����T�����>�6�����gbOm��[�M)}ñא�O��s/ž4��׿���5����Ď@}���c��75��/���ɋϿ��K_���p\6����-�����]���B��ܼ��;|���e��i3{|��A���13=m�bcG���L;���n9"�>��w�q�y1�O�������{�R�y��i�$5�j�Z��pE�xc��BUs�pF�M�t C8߅��Y{b���R��B�U.�aXO��W|f1[#5>��#�"�gp`������҇8푎�`�9�l���3/B���h�ԉ
��V6-�j�S z7�bx��Ӫ�婙xF���Ͷ�y�o���P:;�/ �aX��S� �;�0l�/���6豓�bb�&�\ϫ��W���� X@��"w~�k:3�`%h�S��K�U����[�p���e���0p�Yvl��X;��������� ��l+��v+y�v�闃@�a<��Β�,�=6wj���~t���:�v�@j��u�t2��/oE�g��Nҙ%��a4�����q-2i���+�����'�ޡ��Dke)Z���p�&ڕ5d>z2�<��]�J�h�x�4�=ҳ�3nwf�~�H�zї��0��IP���?�;}ݣ �a�Cq�`�
�iQגt�zN��C@;E ���I[?u>�'���;�&�ge�Rb��v�Wo�?~���΍[�8������I�j�E[�#�i�|�zP����gc�c��/�q��W^����_�S/���Q͜b�g 6Y��L���k��q��{��㎨�?a����o.%��Ί�Ů_
��i�~�n�@�"���/�K��t��3��˗.Y%n�|A���bͼ�0��q9�����w�/�}Bc>�I���f&kE�Lև�C(X������U�ux*��5�1��4S�����0e��3�fձ�8B>���3��\҃Ih���F�x9�W_3�3l)ڦXy�$�Y\Z���qsb�:ͨ�l���bNezFa_Qz��kZ�D������K~���
 ڼ̄��1j: /?�3e)���Kq��^�ђ6(P���a_u^D�]lu�t^����sA��m�ϟ.)*8^��ή�%$�*�nf��*�@��w.9�a'�z��xU��K���D���!"O�5�X* L�08	��3�<T��ֆ<;�s	E6�
�8J/A:�H�N�f�(MU^ʨ{�!�&��l�`;�	�D��G�I�+��`q�e3?'aK����>�-��#�S���L�Z��1z@r�{ȃRF��p5�(�� �d��_��7�)I�e)��T~�g�ξ���e?Y����^��U���������$[���1u�bΞ�ei�l��n��Ա3qB
͇7n��{����g�����@vK����hl�Ş܃3�c�ԙ��|%N��b�x鵸 P?���b��s1~�O�������h��iF�ͽ��fv%�c��LgTŎ��7���}��38"EK���y	���C�Fؓ1T���9�u�l�@����~�Y���s<��(����gU�'|k���v�]&����n��u�u؋IM=�H�ObH�7M9>��� j���%%�Tnݾ׮_�=�K��u^��@M�P�؆�W�S`ъ؛����N9�TX�Zb��,>^�3(`3�ˇ`�+����\��r룏��Ӹh;J��(���L�9q2�ONŸ�1�;���/��j��?�+��W�Ǟ>N��ߺ?��>�݋uu梭��!J�4���Q��AM���G	�E	���q������,�- `�B����Y[��ֹ�n�A���A�g�9�p�2�'�J�MHf	��ԥB:6i,١���T���a�[�0�U��� @�Zw��m� ޝk�y>+�?�r��f��A���S�T��u�/<(����p�����3U�����Ty�@a37'j� ���D�L38�=��:_�'�n��n��� �);u��*}���VP�[>#�k�����o��������w߉���F�7JR��ˏXT��K�g0$��6�;��M�
�B�|��2I�nhh�v�����1~�\�Ks���o6c|l*.\|6fO�����U�[ o����dl�Ҿ{F�b`(��'blf:zf,>ni�)�j��FS�]��}y���SECI����R�Ӯ�_[\���혗�[�|��7����M��~F5sr&)QUj�ߵ��ڸ��B�q�_�����؞^��
��	0�P�h3���<K�RQK^�ޅ�1���O
�^�a�A�9���y�}��V��A|@�1#�*�דXW�C�T���B�C�s���t(��f���cل7Pn44p���:�PGy�����J�|E�#N�:�Ab�u!-�8��ǆ��`�:�F�x�����ߏ���F��".=��+׮��GbA������P�%	|x0+�р4(!��r��i뚯��k��F�]x&�ǧ��'-ß�c*�2L�u��F�j������6ﶧAYZ8�����Q!,�f^[3txM�k�,��A�mJУ��vW ��� *Jp�0���ݺ*��8��ok� � �́%�A%�I���\~U������TUW_�?9;�ȳ+.T���a���7d�c�Q�S�f���Tv��?��n|Ђv�W*p��ν#��5�e���f(��*�; �/<�gfJ�+c��{�q���}����o�B��%�T�}�%C_ �9~�../���3*}>�?���]��*�M4
�J���������ˢK��/EM �.��M)`�ޜ�@o*����e3��V�p��!�
�dg@y��	?)�������Ǣy��V�k0�Z�{�ϴ�K�_Z��V3�b�ֽ�]\����XQܫ?�e�l6�Թ�1���F��լjD���^�v�3ˏ�%+k[�����r�
/h����~~���杷���.U�w�@�u������ivM���LJާ0��b D�/��H��w�ލ۷n���� ��'�kF%�p�!�y�E1C 2�c��܄M� �.�vu"��Z<��v���������M��nH3��3�XZZ6���?�iܙ��T�~w��*�?�ǃ�	�Fu��>� �&�瞽,��L�jnD��GL���Y@BqR`=�i�k�7�&����rr�3p�5"Oń��٘����c13w\@0��J��V�w�;Z;���$:���'�Є�I��M	E9�
(��M @&� ��?	��ҫk�����@e����!Y���2���P�n�A���	�,��6.Pwz��v�8m�H?�$�T�ʒG)� ��`�/u�]������Kz�����0�G�3���;�;Q�ɼF�������aH�k����yC�ϙ�@]�wQ���|�7��r|p�d��q��^����{���6�92��f��7������/<c�7�2}mҿ����p���X���w,Z�����xx���ǐ���x��W�cQ���o�M���X��+�/׺��FKu�Hkτ�nߍ���Ǎ��q�;�������~+������^�2E8�A?�0��
,��������{�������ƍ�ߏ�?���j��ޫ�ƕe`�U�+ܩ���g�0��w^H*6�w{X�`I�8������2���u�����j��[i� Z7��fH�h��h�|�a\��5v@e���!G�x��ѫ4z)Du�'s]+��2���
��F*��j� �'�[WVV�  䉼�Q*,���E����HE�fM�[��3����5?��4G�x��Y���6�	�e?1k�c3�q�����R��`hD�~�q�񼿂�?,mK@ދ=$�aiCr��*(%�,��`��t��you�Ux>��RO�ǝUvO����a^J����Zov�Fe������\��6�a��,�rY;�|�S�D*���]���a��6�������0 r���A"��pJ����J�����LN�-����r���v��Ԗ��l+�vxl��0NӜ�x'�b�M��8*CB
�A�$���[+��<Y�d�f<�ߗ-TĠ/xxڣ��YȥɅ9���Q�h�> V{���#*��O���ַ��>�~Da*��\����`��Ɩ�� @꿲cϮѥ�J�q�c\�L��?\�����k[k��>��fʛ>C��"|a�����HZ��b��T�J1ړR���H�1�ù�|����ߝ�(���P��ׯ�v�'_x.�f���ٮ�~�3SV������}�h,�Ǧf��#Μ����;��6��#{�4H���k��{�Y�
t�EUw����xo����y�\y֛B�f�bI�|��_����'^KO�8�%-��H%���L�.�][���o4D,	z�'&���~�#)��K�"D�W? ��M)6���?�8��4�˦�S^^bf��э�� ��a̥S��ձ�����m��h�����9ծ�J�~vذ�~]�l�o��V��ݍǜ�,p����=������_��'�#M��Ɛ�����Xƞ�~���r�$�S��R���5*ᝐ����ΐ���F��#���tr1�����k�Lk���wǦ�q\ �
�Qnkƪ{?k�t�
�Zu�2�J�I����ş4�a���u�����r6P�Q���u��>��s����G�7xs]�t}�>o�%ȗ��ͼ bj��}��Wd�W,�yג�L �Z ^vx�[�%���,p$���vS�}�]e���)������Jo��s�Q��@���G���,�=�����{�G�(�����f��-�K�0�w�t��V���_ղb�֬�o�����]r���^2���$ �T읙��'�-��d�vGFx�{ky1��nĵ�̺Xf·O�\�S�&��&c[�aW�2 y��V��N��L.1���Kq���ų��[R�Z9{fs%F�#r��U/��ש���`����l4��~�]x�#�N�����-6z��ER�ҟ�f�O�mS��G�i��!ow$�R�b:�=d�?�v2F3�m*B��tr��:q빐Fa���M������Wex�A����A���@�N�D�i�l�m��K����lI3_��7�5�g-���e���K��Y�AI˼馚,n�Ǜ���ߍ?�ַ�k7bG��H�)�4��[�X�j��v36|Õ��;�0}n(L���𡎩�S>B@*~�	�v���It��n�`tCe�A3I�a��襀���G Y���;x��T�*��W�K�����ኍv�u3uMpL���؀�ݴm��'��,S}j�	�p��||�e#,��a�K���S�Q�y�|)q�fցNՙ C�����N ;�D�R#PQ<�5-a��� ;��#�2������l�K��cː���.��qd/�h�òG�2#f}�ʓd[J�"��,� ]���&��:��h�ȋy�2{ƮH(J�h�J��
���G~��q$})/����u͎��Dk� �����_�+�[���������'N�.�Z�2m���!;��(ഖN�G��������|5�4 �J�j*61�\fb�/�����3b�ʥ9.���q���c]�Z��������mn��ގ�p ��Uɥ���v��������������+v�x^�;�mY%>�2��is�ڲ��;7�m�g=�'l��&�IN�E{G� El��_lv'.T^�� '=v��q���D�j�fS?/�9u*�\�/>�B�>u�_Y�xQ?�V�h譊|Z��])����{�Hn�c�'�"�k�-��:�T��d	�_""m�-u��ʾ�[Wn��m忨8�$T���X�mE���AMi�ŷ�AZ�CW�IR���>"opX�>��igxiML|N���]Ɂm�'apÛ�6!r�9���X��hi�"@�N��3 ���\�y!�!ybE��-�~	k0U؎�LY�gҪ�$� W�^#ҳ��8 %K��\w�]��-sW�ʠ��u~�� �?��A�~�<*wu�E���*O�My<�F�o��;K�<6����_I�<p���$�JI��K^*�P����>d�:�[�cyV�k�+��9CMV�0��cr-�A@!���T����F6�w��*ۖ� kXr�����e<��^,��(�֗c��L�����럋׿��8~����b0a&Zn�ĉx�˿#���Ҵ'��߈W��ߊ/��?�g����� �T.JK�j��>��]Jc1s�|�~�x�����3�9��F<�W��KJ��=��
�]x���)㣇��s�g�|^�pQ��R���!��5cf1���%-�`)�<��8S��{� �<-�	N�2z����/~@*pԔ&���)#~
Ϗ��`"�,w�t�Â��f�C��>y6���y�g��i^��s��gݗ��}J�e��r�5]�͗�h��g  hM��(105���Y�ѽ��Sgy��4��n�*���m��6�X��	�7�ǡA�b@Scg�mVr��R:mI�eR�gKI�Sg������O��2MC�}Y��r3}W>^�A�Y�O�_�y�ь��� �p!�#5a:�)f\� ���k �@|��2�z�ΫR������( q��%�& ��m�������p+|�]�,y��W�}�F�9�n �=ʉ�zFT%��(��y�Z��;��GY)����`g��L� (BƑ���������RV�[@y���h��jy��U�1k�P֫��J{��,�TwS٢��zW���Ҷ|����K���ѼӢ���*1���G�L�$��"�eҥ|�)>)�uoOj���U��ѱ�:}&��IK���[���[��6�?�9�TfQ�663'�\�s���^~��'��P>-)2(N�Y4ي��d�%C����M��N"΃��>����K1��lb��LS"�)G����˝�^��G?�3�[�]��1����*��W���R�Vs�'�Λ��K�U1=3cwɏLJ�]?� ���τ4N��$^7�0?��ͨ���7o��k�DMoC���J�E	RW7�5�*}��/����������n��`�A �mu�{����f�/.h@�� �l,���LO����PʒZ�;R)�Cn�갈�b7&�*b+��5��B����B]OZ���}@�¬�FQ�.���e&Ы������T�����)U~G�l���Ɩ_|��YS�K3m��������!yX ��ÔA��|?�����}�yn{�`[���mo�Qx�T?�<�c����j�Q'�KZ�]�˸�s90����h&�9׼i���ZҐ�+���\�����F����F�Q^@�5v�f��pB�[[큶�q�O����f�-+6L�yo~Ҳ��	�Gf��� �ල�ǦWb_���nY�*UA>�Pxo����R�.�=�<���'�s��}MN�,���7pH�~���5p�-�M���JLH����n�V�����Uj��~�#^�'�UXq��FM�7�>�c��e?A�Y�d�O��\��[_��s����l̝���	ψ�����iڏ�~ꀂ����rW�	�G�5@�l������R��恮Tf�O�������x�QL�/���M��2'�hn�H����nl����������oZ~X�f���t(�j ���?�q��g?w�JZlN�]i��}�s��K/yy�3�y?	��Sk�GM�M�t
�V.\�E�Ν��}괴l4�ӧM,�p͑ �U9Դ�O��V(o����affV���]�ON���Jܼu+�3岉Fv�h���M��NhA��6���Q[u�O�m|O�* �XX�P:�(����-z#�%����� (����
�r����4'N��Ai�h���%[۹&o@R�͇mTeKz�f�y�#�,�m:9u.׺ϖ��^n��g��N��t2\��u�uH��D��DI?�r���YU����ܫ����}wX��$(�.�<N��4n�|�2l������"ǹl�ınM��[a� _-.
oȟ�[�yl��Q�����Y��G��"?�c�Q���`�/���jk����۱+M��tw5`�
���Y�;*��-L4��hi�������>�E�`}�s�d��y8|�����׃��|���x�xA
���!�L�4�,T���`�6Ő!���ȥ�P>�>)9�:}.�_~.z����Ǧ���R�$�~SY�]Ջ.���W�4��
��z�jvj����Q�T	��\:HY�J[��������Z��/�p�=�f
��8�k�ޣ���G?���7�=�7s���x��w���+�l������x�]'��r#�[�F^�́n���-���!S"�#���k-�=�.\�Ͽ����������<s1.]��'�Х����	?�9� p���������g�7_Y�%�<x�o~�e�ֵ�6b���u���Q�hWj v���������O���3��]�sM��0um� �6���J��������nP��ʫ<؉������u�vGux�B���'f �Հ�w��l��h��Mvvw|��y3�@�c��U/�|�~v��<,�Չv�J<L._d��d�L�N��=���-7�IC{6�ICa:y$U5��?͔r@���*ud?xU��a�ia(�AP~�o�Q�R���e��N_q��+��p�>C�����-o���e���fls4�����r4�����zQ[�����4U�� % �M}r�<ͥ(2���Jw6)���h�ǎ�/}�K�����r��.�3��A��{�wQ��O",����f�U$N��k�~+�T�ёa�lc�C���O�-2�\�~��~����6���Vp��ʃ>���.���rl6D���*�S	��e��Q������n~�Q���s^���< l�K�(��a{�Ϙ���Q4�9�j��e�0@�P)_�-M���S#���N��q���x�3���N��� �Z9�g����m�O������Lh6J˻L�#B1uk��c]Z�z��yR�VC��,I�[jP�ׂ���]���v���#Az���À� ������v�����fz�c�cdt:�Ggbl@Q�X����H�p�� ���I8������ԯ�i�������y4�zi@��H���@�:=͔�)n�;`����k���.�tZ��t^�N��x ���^��ŏ]NT���K>�Q����)怰��H�T�-{Ca ?���>ow2�(y����=Y��lLw��z�M����n�+�Cz��:n�p��&�yB),�t�h�U+������s)Dr!7~Y�j0����$����v�sXRQ�|�e{s+n}t;����xbD�S1;�(�Í<�g�+��/E�#2�2��5k��*)���9S�[��Ǜ�'��|7�$?>6B�|���������GT./렔� ��ɓ�^��t�d�	�(�|T>ꁱҢ|hOv�4R�e\"%�\������W^�3Hp�嗃�|��� �j�+�������L��9ʝ��08Le���/n: ���WB�#Sh�3�J��fQ\U��N*����8��X�֬H��KB!B#�����ZSSfi�M5=� y���s�9�s�?A��$zd��5���]�_��S�7:�#��?<��]Dӱ;<���������h�����x���+?��U�U~��{Ԩb����b�}H �♂���̓]�������ݓ-��h�4�:�T��L]�u���c��dX:m�Q�q�T��vY:1)_�~�S����pj�YĚ�@\�Nw����́z�M�a�,���"�l�T�w����
?�2 �J�FiJ\F�Ay	�x��20�~~��wU65������yÕ����a���xs��A¸";Ȋ���e���ܗ�lq�������?�fܹ}�3f��h���U�3�|F��K��l��;����5�"߹ޝ ����R������?��~���z�0w�1�{���N�=u ����Л�W	ԙ��#Tb��%5�m�Mw�C[�+��|ĳ!p�!H����
�M{��^p#�S�!�r�K�^��1�1����Lue��wG�;�@e����o��U�Z��	���
p �m!w��\L����*l
��8�Q��|�����e�JlrL����CJi�;��`Җw�{X(�P��8	��A��זE�{��OD�@�w|&z�g�g�X�͞����b��Y�OGL�������4k`*�&bMi�*�5�������m�vU����3+d���%f��Oĕ�_� 3-�b���>VAug)�|��JH�}H����s��10��aý�!�WT��+���l��1��u��n�u�q�T��:n�%��Z�b��+���<ܫաt��|�2�&]@���[����� *�x�`� #�@�C�� �<W CZ�5�������[��Pԋnw>��E�l�)<*e��t�(Oj�]���X�8���_��o߉A�%��e�� ���lx`�,���ZK�mOMLy;3�!�LL� 緰f.�vb�@{ �H>ot�lʹ{��*V?|7ƚ�1��@=����Y��Epf0��W���@a�$)�3si3g�]R<�Ҳ�D�}�p�wJ.����ɵ�?U
 ���z�ʕxp��W1���s�xvH��
f49`b�2S���`U�Ue���us���t�"��Q�Ŕk��P)�����G���43�#i{����x���k[��g�F�!P�e<'"�Z�#Ң�w�����>i���m�V��F/�` ��!���> }�T�L����c����謩1:����7'N����ؐ���L�M
�ǣ��8߂?h�����[/7��N�Iu��ھxU�]b|���7L��[{�x��v�����G�2��N��Df��|��#��Z�/k�i ��5��6{� Cp"�5�P���w��=a��;id������L� (W�8��e0ڀ-�K�#��r�:��r'��?��dP��iw�SI �]e��ljl�'K��ˊoeG��7��Yw�-�,���:-��kS����(��j��ձgP�[,���4S[�k�z��$HA#�i�Y�����m�/�-MNŤ yߑ_~��3S���vC�c[��f����W?�7��Gњc����OPfxS�	꠴���i��i��<*��9\��Μ��g��j��iҁ�2�)g�*wjx�ུ�hM�e(=İ�����sh"��V?���M�d��rvY�9���!�m՚)��L�{�k-��Z;���t)�!� "3N�_v�Ս��}՟�B[oI3氠]i�{Ҕ�d�M沈��}i�=�S�6�.�Op#5 ��������=�X��{w�x�E{�'cW@���ϝ����������y6��3ќȏ��'�"��H5xn�D[χ��y�3
�2����׻|$ ^rQ�D���56:g���2�a B�m�������7��h
M7�~��G����:m{ ��*?ޕɇy�%o��D�AH��E�J�0�ǽ��T�42�nX\�[�&-4 ��ţ�	���%�$�c���Nr[��m4<���h۔�0���eD�}	�
CYq/ɻ�z�������9W�N���E�u]�Q~�-�{#���Q-��>���2oO��\L�B�\2�,��Lz)U�R'%!�g��e+3��@�ް�܊��5U�)m�,�?(���Op4�آ�W�x��?�� {s-������غ�^�\?�ߋ��F��/v�;�Qw�IJC�܏�c�xa�q=+���+��o^�Cm��}�G �qɒ��!���Y_�9#��Wl	g�c�#G�3���ϋ����^�}��%���_����T~U�z]�*@!�l��{�IP�8ђA-���C�YԮ��]�c:��A,� 4Y�ߐ6�Q�����We�e���D��l�M�E�Ա��=4u<����
��deG�:א�}�&�}O��M*�l��ƏE�h[�{��I/��<C�.D��s1p�|��}'��𙋺w.�#S�f��x �]�R/��	���!Z�{�Rc/۲��.�JAD��N���^ ?����8Òo;�a�c0�ƝPv��vǓ]���
�$ү�,�t�i���*l���L3�x*�J���C:93�|���VuT�"M�g{\Y.�S�0�uO�T@7o6��P�'�/����t��nP�Yp3���r]�!�P{W���_����w��P�T�U��"gv�[.菵�U����J��� XfE������=+h����N"�gn
Dz�޶�3����?.z��p�}\ߪ�n�n3�����lH�]��w3n���q�'?���V�V�OaB��b��Wb$���'��и����̀ ;��z��^��t=�ډQ�3hDuR}�΃ꊇ�[����|�#|�t钏\a�_v�0A�@a9��}�]7ȱ��ȟA����p9Xu��~������4��v#*� y���%��a�W��"�jk�n�t�G�7�X�
˧�z'g�gB�. �9#�N��ܩ�=6w2Ə������cii� �4����;`К�$����>. ��>6s:�g�*��1<{:�f��31zR�~�T���)�y�\�\�s�İ��N�RyNhp��FN��~�ګѹw@�K�%j�ܪ��.����: (�ի|���ɭ4��0)�)$�6�M�:��wZ�C+�l���$Q� ��ܷ����D�)�Ҏ4+�\�� �5��%��fC��Z=�z��:T�.��Ŧ�Wݧ���PG�� A��W���\�U��3���m���ؘb˸]K��m��;u��G��W�>v����+`, ����s��yUڙG����AE�g���l�NkV<(�J3U� 
��W�U|�@��!���A�������F�Ʋ�o��ۖҳ���&��9+�ǳ<p�g����yg�Ӏ �ѾT��F0Kh��pk+fv�1�jV4#`Q��P���,,�+��������oĽ{���3}�&��CM��J�.�	���#�2(��g0G�^yJ���o�_������Y�m	���q�ᙹ�<yF�-�9�@.P��ߔ@wR�:!`�=f�giF���-!bK$�y�+���Hi�=
30����K���\2��L`:z�&b��/����P�����T���gc�� 30A�)MX�O /������Gc���jX5�����|���?4B�t/�/�ƴ=��p�RQ�.m1���k��W��k��2��VА	��a,p�#?��nR�Jg���Yu-�e��2IYղ��ͧ؎2.g�n�����p�\�Ӫ�o;)Ө���l�y�1
U�����ʹ���ғe�:˘�~j'ʫ@u�5�5(mA��E.;�Y����L	x��`Um��c8bd4ο�J|�k9N~�K�x�D�Q�= �gH��(�oIs=~������(�nG��R��OKs�&>��#v�r���KcJ��O5?�]ϨS�7�܎���^Y��ZY����1��(�=��wb�������t����t��0��c���=`�T���f>q�����ӫv�
���\��ŹY|ސx|�C:�.�������nulo
J�1���Ս;T�U_7�?�k�
���%��!�{��x�b�j{?�Z^��6�6F�V�XIXF4��0:1�/���!}Ґ�@L˙1E�T��b���wĥ���Fh`��Z����A���I��e#]k o�͛���ᰡ�����ɛu���v̝:.=�������F�w8�[�Y5�.�fï���a�Z��jܦ.4�60`V~��H	��n ��s�rOv�Q���"�~�R�0�����<���4;��|���!l1�ȗ����O'�e,��b�`�n�oI�8��� ��)�gN���W���q����2� �1Ɏ�!�UopZ�U?�h�/�֫�4MuNb����4��x��ּy��ρ�%�|A�����LL��ܴ�gW�у�<�&�����g���\R�U.�[[��%�h��Eʹ�E��Hl���?a�4dR &)���G���݈Ƿn	<G�A��ёQ�o�E�ڶO�eCZ��f������G��Z���D��j�/�D��rȆ�W�bzs3f�7e����j�o����jj`a�F��,��R��<�|!Ck����~'��̳>`G���ڪ�ё/d��������/��������HVϝ=�-�V�0�Q�����L'q��G���浠���R���|jWt|�W�)3)?���X+j�U_�n���~p,R�Y������^��sX��+�<�W�:�5g���(�]��DH�~X x[�A'�Ј����k�("-���9L�3P��Aں��~������Əu^�Z �KW���rLiI1���7�w�7��&A�L>��/�h�V>��T�bgT�4�]��:�#`�.|�H�n�i�s�>��G7R.)t� 7(�E���Wm^�
���?��c%/�O	󛀝+�JTF��h�ħ�`��.�)��7��>���>�1҇��Lu�,�v�EYJi��ʥ�B����a�yX�XO�V#k��������$u�5��ż��CM���L4h�u�X�^�@�T�ʉ��<ø�U��(<-�T�&I�n;VD�$S��ǋx(<���x�?|]lr*&��r���n����eJ����!>��@l݉���w��pN��o-�Gca!v��%j>|;�G���ؼ{'6�܊����ގ���?�����Vz'z�ݷ�1�����jmF�������N���K���\�~-�����W�8���1;;��h��SӖ�NJ�����*��>*p��ŋ��ug���ȶ��i��IR���(`!pE�_�b��i��yڔ���I� ��*j�
��cM(�%A]m�c~u#V4/.��Ҋ���i<B�`����)�F�!Mk�2I×`I�Z��-	�.#���`Po6�cK#oS�v[��1��iIP���Z���-@ w�աG��?01}�3�;6�}����=�x������c�#}���`5ɆwJ���L
UvZL��U�ذ�hr?���Iiگ���T � H0JZ�i��O��Av��.�o��(CR�sE�3�i:~>��i�')W�L�|��GW�ˀd�[�$�+ͪ�Jٲ.i�S) ���c)�ʠ�� ��P�;��z�,|x���V�OTGqZr�ߥ�QQ��8i5�=8��6��cF��������ii�3���� 巴����������4?��u����~��X�ɏc���c�g?����4�~��h����z���~���~�h����:����el~�V�ݛ1�x?�V�c��#�����e�="�"$�^w%������	�����\�3���{@xÔ7O��i<�C�)
|+6�k]z�?��$V�v,�\'����BzC�T�Ty��A	෤�oi�d_8c=~8+˱��hF2�A�ѲАx㇕��H3��g�Y	�57�iq�v��*~�Y�7<<s��>�ft�c�1�d	�Bz�lԲM�@����k�0$�d�k� ���t���fC����F��� ��[gP�h-`w:��6K�H��SwW��N���#"4������Vԉ����{v�4 !L�3N��`Cܤ��L-�LaSnӿ>믄L���r6��⮓������TI�
Ӊ�)L��I���>6�vi��2�]/@pN�F�L�%�3�� $��N���-��:�IU�a�d�u�⥩�>��%��W��&��[��O��{g
ˈ���*Qs+_� �������Ao�������`��:��V�{�5c��6��p��h���q�{߉{?�Q����������bM��y��h��0v�߈�Gw�w�a��.D��b�m�D�֚5s�[�w6Cs�����{�1�B���쪪�k���'	y�<|`��%�\�<v����_�ij �*�Y	ăU��}�Y؀�M�۪��d�j8Q�ya�.ܘR�uC�����=�-���?(�}0�e��{����ѧiٔ4��_ xpP��AV�p�� dHӿ�'c\#���T��i�{�t���yf.#P��O(������sR�Ѳ��)s}����W�Z�Z�>"@e��<i�c3��d?9&���~۴" ޝV�%�9v;��m�_�����S��I�?���F1��BS�u�f�[�w	���MR3Y[��O1u��҅�,�|,U`������|2o�xzO��<M��5^u�YpŃ2� ���e���'K���?�< 9�1�1;ʰ��R7��T��|*TL����y��ï��R�f�Q<lN%���om5V�}��7c���h<�{R��6��W���G�q	.��@5���#���'�g_s�~�J� ��Yx�K���|�=��ͅ�mQc1�K�5i�*PC�n��˸��ۢ��ߎ����C�Y��!PrF�;8�2���f@�|�rܾ}���z����B����N?�����׿���|6������I�|��|��$�_�����u��n@Dy3��9�v�} ���>/��hҗ.��TnΠ�H��I��h@�g`0�y���񘘛3��LM{��d����g�]5�����$ԙ�X.#�k0WNyYT�A����ҝ9��ǣodB�?�zJsev�����X�M��𫈕����+m*�W��2�r�Z�I�g�N:ِ�L=T�PTq��s�o� � ��6xT�T�ҩK[��b�o1N�"���ArϟQ����<e��C�J�?�)�]�8i��G1�����1�v�_M�3��Y�� �Q �������a�w����d%�n�t���:����vI§�I��Fܫ�uޯ��v!rE������w����wo�����-wS�|�Nl//Kik� �PLH��g�۽��N�@��I�b���kF�~S�����5���1"ܽ|Ү��������v촶�!�/F�ww$'��L(��|���U}́��0�%�m|l���^v������u�oC�);d��"�=�+@K�~���� �<X�0���4���p���f
��M)p���Nl�����AxC�m��K���I��h�p6.<w).�J��M�Ǌ+>�:َ�ɒ`�ӥ����z|�_�e�hx\�.�s����'�0|�O����iYi$(���htS��ei��G��<���/&m�^P�����u�����߭� Rʣ��믓�A$��⏭!!۲ܗ?�E�.�VuA�M�J�.��1Եl��T�N>�8<�*���V,,-Ŗ4+$�@-;��9q,<�� D]�b��>e�n�h�SK�ˠ�K�`�L�%c���?l��ڼ��r����2�)e:j�����e��u�?��'݇v�ʋI~>%�Iྯ��?�,����@� �O�������
)��> � ��C�}JS �X��t]� ��Gڼ�!�e֣k�0�zo/��]Z��.ߜm$�<�\����w��p��é��_�ь��xS����މņ�_�~=nݾ���a8n E@�)��Y�KcA�����t�d����@�i�0 ��">�&����Go[�$mi~}S1v�x��������0/{x�FB�9�`��k��Yv�?��hdb2����E:�:�^��4^�b���v�x2�Z���&ۏ�Jk@ҺM��[�\.=�:��O�a~e]�4(�(��Xu8�Dv�:��q
\2���a0Z�Vo��U8�*z�TPT�)�fU��n`O6BϚ��Z�R��ۿɐ.�`� ��Wˈ�G�*<R�9\���-�A��x�!�g'�� G+�y*�<]ae'<qX�"�����^j1���$+����_��C�H[�dw��S�'u�t]�0xԯ��� �������K�l���HHn �OZ��~XE1 ��gޮ�w�����7Zq��Ͻ�>4y=�mb~\[��rУ2�uz�9~�S����Ҍ� vss]�E�'l�M���4���-~yKuf�����6X0�����ַ�?����s�;�C��yޠ��-<� W�|o����v��lݒ���)�8l��v	�5	��nhJ��jƖӐ �
�����x���֖b [��έ���)]�f�q�
+n:	�\���Qp�������LhшAy��Z5Z^����a� �{��Ye��1�l�< V���P���S�ѕI�����T�3ΑF�EP�?o%�V�
�6����6f��Q����'�=͔4>(��(w1hO��m/�r�Tg���9u�De���q�)���)oR�F���	Н�� 
��ؽ�> ��gH����t�~~�%�F���e����;�"®S�3ڧ�
M�s\��z��wW����M	L\ʯ\���o:>�HF���S�{���G�7+�F �i�(��U;�-K>4_�Y�����G\��l~R7�����>�l���R<z�@`��|$��8~U�ʮ���Г���|yđ�R$9͑6F{�v횷��:2`�B;�|j���C<���Y�æ��&�
�b�yC�]�"�"�W�Q�l�0�[59�M��&aX�<�J��0;��-/�S��ö�&�ا����ƌk�=;g8.���Cj�5K6�:K0�3u�#́��y`�F�;���[����ſ-0��>#~NUiP��S�Ob��:��'+��H��1rv��;Fa(��P�x�Ai;�
�,�����N)��7��܈��~�<��i&k����+�Y6����uN�r��������a�?�%'> c �<zp�M��R�Y4v�O����"�h謯3kx��oJ�ɟ�[y��]d�B ��i�nk�\},��&%�T��4�.p/;��!wڿPiwv� |�!��Ν2-�>'n��,���\ڄ��9�IZ!R��%%�HY�`W�'�Om�D�N1f5e�� ��M����;��XZ\�q �$h�W<������<�8_�3�\�_��v;ޗ��jx;*Z9�0���i*g�@�#8: ���+
us��1���`�T�4����$&:�d#%�Z�b�ǚgK�9:`k�W�'m=��;����h�l������fD=�]�ߤ|�6�l�����}�j$�}ר906V�a-=�e��� �����;��+��᪵1l	\�^�Ay��`$G(A�H�u���*��6ݴ��5'Q��lؤU@���}�3���o�s�(r~i��\�����f�7��f8��e��D�?������q�g��6+Ee��m����{)L��uCj�"ì�er[�_P��d���'_?�D�(�A�_�G^���[�])m�yْ돶�MWi䢁�$7���2iY$O�ӕ�BE��}�tۤ[�4�����_9���}D,3�u��&���Wx���bW���"� �	���)�N��J)�"k C9���U�ңy�����A{�w�����ݹ'�=i�󱸴��+�Hz��^]ƽ,��X[]uy�2�/�q���@�}�<�6�5>�7'@�ҥ�����ʌ�n�|�$� �)������|[�H`�F��	s �#������q�UǮ�F�ww�=�������vo<j�ƃf+� yMK�;�:��ƃ�>�9��SeOGU�l;_��hIy�� ���<���}^���JF@�<��]�*�)�|��)@��L�`�e̀O}��bPe�f���W���	Fcc=��{wG�Ri-i��V췚��4 ��lȝ<��f�ͽ�Vޕ��C�`���b�y���g��V")�3U�0�6���)Z
aFG��������ִ~���>Za�S�����(?����aP�z�P:4KL{_�X����ݽ�`ʏ� �@e'��$����h�.�DAeL.�H�R��+���sa��q;6��cGe�\��
��>��:�N��-`h�#뭍X��Ql,<R�jN������|>JΞ_F�	��D|m��~�oUR�;�莲��;��1X�W����M�+��r�����@x�+e�� 	��gߡ���\��(
�-�*r�&�&ѷ���z�D:��1�+7=�K>��WyRB�!�/�i����.2���,���	���Rx�W�8Jy��774ѠQ��Z#W��"o�NOMf~�4�us�:1�2�{�D��2+T�#J�V�J�W�=�D������X���5|v�܀p�������z_��>�Mr��ʒI6\��%_��@���Dh_��/���|����ո�qq�@fl��ƅ���y���2xT�\�AvK����w/!:k��(�B1a�A���W��G@�v��ѿ��� ��0~�Ji;.嫹�g�a�u!{��t:٥-�nz0%_�;��Zp�O4w�j2T@�3��GD?��{mx$�`�qY�s��4%K"��!Q�]�`)�N"�1P�#���*��9��A.����(3���g��@�l9U��l(c�d�sdy��+�98�K,q���l���g��t.��Ny��O��TW�æ�o٣��I�
%*�,O)[�^��+�T���B
�ra�	�*���������C�ǯ��t�<�5#@wfY~���T8����y� �gY��5r4�%�񮮬z;cx�=�|���ɒ8�A!�Ax�?}�@��e�<��#�}ؔ�0�mkT���Ʉ
\U��p��4�x��%��m�����%�f	fM�Z��n�٭
cV��6(ۤ�B�%�j@�����8V�/��Nl5 �3I���3mJk!@�+ʜ�J���s'e<��[�d�����W� zip�o�5]$?��)D^vO��\U�t�R.ו<du�D�C��ke,T7t:��4x�e'�0cȡ�%��(�ʔZv�>���>�N�n�t�hu�v)��4�p��G���-��!jD��pwX�cqG�ܔ�*}�x�L����p�k�����r���a;��bU��52�k�I���{�U{B�еlfy~����*��IWrJ]`�����N����u?Qɗv�}�
���)���T�nH�_�A��WK^y!��?�d	ߔ
���hH3G^h��V��<�ad~?�(33dC}+e>M�~����=2��k��r���P�&j��7N9��kd��xpS��8�������NϠe~T�iL�7��zt��_���4�o"�ux5��}��m��k����)Y_//�vbP��4�L:L��f�0
���GF7=*wv�D=�� Ab_|V�
O�J��tv:�>� �U�9�_��}�����}����:��2}W��{lЙ�@�'��\Fl�S�eY��)�&ç�/����8�S��0���T�'J��!7(~�f:,�q��&^�> �E� ����J-���
D���+��+,��������}�B�K���nĞ@�`�0Ud9+����Ӯ�h�<�4��gecJ�%���x�>��
y�?��4�vK���gQ����;��}���i8���@�3��aY"Dg+"/G���A)'8��E����I@=���#ڻ
�~_���㫿�U�CY)�ߖ?�~�֔���=aJ�?���<��|��es�#����M�Uٿ�?;X:�,������!-��^V^wV!MR�x]�����u�I�����N:���6�� m�S�x��s��
�4��@j�؅ԡ=8pҟ:�A=��2@���?���ת��r�6�w^�9N�O?x��*���'�r>��Gyٮ�1O��zT�
_L�sǭ�;�j�JU��H��r�c����ǵ���Y���P�Hs7�6}�f(�>xȳ6�T�Q.��h���g$��fUR��;��`�g�w[ �8T�6�ů|H7�S�Ic~�Ș�������չu��%a����.T�i�o���M��_���8�%�pIy��8T��'���G�PF:U?�?@��A�� x��m�e^jO󌣥r�@��&'���:�>~�";���_����w��-��4J�Y�y��O��MU�CT���`B�%Lap��9|�N3��~�>H��>���DCQ9�qK���aS��n��La-JO99�4�']��(a`�O���Ic��妣C�d����]����:��2��_7��U���Ͻ�ZRӰVSֶ�/���ֵ4.�V*�\�0R�1��q���2A��]�����U��O�J��ҿ��@^Ŷ$�3��_ �����[��N��+�?�qM�S�[��5�יk~n?���㧊f�Ҕ�tCi(��d�3����Nկ �K̓I@�fG��~�~PZ��Џ&^���7+i�M����a�櫜�t�I�d�C��L֩�����⾋<�!vk������VJ���I�:n�*c�*�H��"nձN�Aܽ�)w�i�I�u�Z���^�_�t_l��n�$��Y��Gz���#F�]R�ǔv� E�wk�_��8i�/�A�5�Ń�~�t8��:���,gP����ĸ�(0�̘us��ˆ#h�<_�NKJ)��Hd���sq����[u�������'�l�$BdهL	��:�/���S(�^�PM����z(���y�� ՜v6�=Ю�>#��V^	�T��-�b2U�ܘ�!���J�K�
�����e���g�²�����͵��X�����Z_���j46ף����,�$	����wӗD�:�lA,JU&�{����Z��[r�\�}�t�x����2ɋ4�)��X8�d!H�#��N�ڼ
W¦�uѤכv�͓�䂩rJ���ȍ����N�\Z�"TT��$4x�� �yk*�Oк�Y��-��?�|�T�S;��)=����D��~�u�[~�Iݦ2�_�J+�#���7���,Υ;�>I�4��d���%-�)��L��hǴ�u�+�*��l`2v��x�!O�ݍ�\�΢��n�;28��5���Ⱦv���Z�#�"� �uw����+:ך܄Gkgigrj:����ם��[:`(|��n
o����iJk�u�X�d����0������RG�폝��X�am}?6%�-�Ǟ���2�#?���+�K%�~2�A�h���V.y��	�Q�%��hT��&[�ԉ�77D뱱�kˋ��8����j�K���0�=�Ň�m/�����X^�W��w�费���+!a�]�5���mb;��n�Zv���d:h���_bh{K������x���J<��^J����bX4"���a'M���f'����L\<{&N����Ӂ�fh�t�e�t�I��~��+�:��Y@�34V��iu�WWU?)����B�0죈h2�O6G����,Cfxtz����dy�h���1��>Pj�����������>Bi�פ�g�����|��C�J�N�l��!,<�D��m�gl6������w�U����U��������?��m3�3� ��P�	�n��~a�7��"�7��7D�2��N�r�+�-Z��Yb�!�6$Q'�S������GRտO2��p��h�G��j��Gk�q�,=���->�M��R����Z������Y]�ݥ�ؗ�|�}��v#<ʳ<yO[� ��ILm�
$(VИEL�|���A!�����c�j��!t�N����q~%�Ӫ�ҝB�S����I�t�_	w�.�B��B=)�vѯۃ��!�p�B���a��%a>p�"����'B#���m�Xo;��ve����P��pO����Sâ��֠�2M��^�Q��hPW(C���38�E�{��X�S<xR�y����K8։]��]u�qﰩ�}��寇)&�s��A�>��6,��r��L�~���k���2.by�g��+�)����#�ib���`�Z6;Wfgfcnv�G��Д�Š��n,���=�x�;�0�!�7Y3�S�6�����c�pƕ�1u�'1݂�G�O*��]�1��q�qk{?��V�E��� }�k�KC9Յ�$�zʺ��*ҕnk�����4$�٧��Z�>��<�f��P ⭵����t�V���(�*]PN���'��811c��Cq��95|;6׷��~sm%��mm�k�����֔E�D�|D��g�� T�&7!u�W�0����1�1�����-��F2�K�"'�'���0�ȯQ� \���J�[e���b_1Y;#t�a��ԯHC�T�흶���#v���9`*�_д������sݕ)���s���G�P�/o��[��dJ3Jvym2+�H��=u&65Cd�>,�j�ݛ�%e����&�0!Q����/���/��B3=sB� ܰ�g8c���Be(+�>�?ڻ���?E�(�i'�l��+������Y�bC�\��y �%,�p^�^����-&�h�X��<؜�e}=��Ьm|,��ƕ~�� �?�'�$����O#�<������g}|g�+_�r\�xQ�V��%/ک�A|G����6�?��'�����)�3L�����5��^>m���U�3���G�R�����a?�Qv���	i^S�Ԧ��ME+&E�=��="{H4 ��_v�>�e���F�$Dx8�GFbtx$&�'Tj���J���o|�@It�z)���A�A(��C�N'a,��p}�]L�w����!���Sd����<U�4ſ~�p� 10�$/JkftTZ�d�T�;%�K㢱85���ECI�P���_q�GL��D���A�ۉў�4���?9;�m��j�<|��>e�^d@�*�"%=�W(��uC:�'��R@1��9O䱒7o�/�l S�y�8��-�qZ��C��"}�6�F�^�7}�+	��x���4LU�߳�-S��F�ip�^����)i�33s1-m}rj�� ���Zc�8���a�v�P���cv3SG�WQ������j�4ZV.�Oc
��!͏7T05v�"��3w��[q��K{}��������|��C��R'���ń2V:�̀����]��K۝z���05@��# <*h,<z���^|$`h�LϮA|P)�h��yTd�/�]v�`�_�9A[�j�ٖާ;<L�S'O����Z�66�M�]��]ij��-���wim�쌩�Z�ؽ�Q�Co^�Ce�]9uIg��V|3(V�I�]Z��LY�.]���tH�t������QA>�Qp��j�-�a��&k�q�:5�],�YiTO��iW���.M��!��Z��O>��I> �6�A%rS:���mݒ��ď~y5�/n�v[2��^���4�Ϟ;����Z_����h�/ǆf�M��v6%�ɇ�yD-ZyO�Xc_P66�q��uyꁼ`tU~�	S�nE��Ddh��3,�Nk�*{ig��VT��xSsذ?����尯Y�(rJ��<0��3��>.ߏ3�A���c����3ƚٙ�R@��h[Fء�����?�g��Ɍ������P��H��}��s����uX��)1�|�}<�����+�uS*��Z�ʎO��bt�7��r�� U�k�-�������!�GP��g�A\�4���G�c������>@3O�鑡N�I	脴�1�~�V����# o5��iDscֻ�L����?����	�m������5��㼚��T�M��-lwE��=�������fY�12$��'�nN��	O')j�M����-��h���������@�.q�XK���Pj�pF�f�>\xغ��ڊoVno�.y�I�?nl�O��kӺ�+g�m�Z���$̕�W�ʕ.�&���7ވ/|�^� M���D�����L�l�7�����ݾ�hJ��j����r,,������8�o�N,�V~3����yȊ���4���Mi��?����0e�F���I    IEND�B`�PK   t~�X���  �  /   images/5d57974f-fced-4f10-a93b-7d150e366d9f.png��ePN��)�
�J!��"-<�;��
���-����P
�)�ZH���^�yy�y?<����ٛ�ٽ�۽�E����```+�Kk<i�')�>�~$�:O
�I^�����+Ϻ��4���dt�4-�<�]�1<==�Y;غ�;��st��9��``І(HKhy��y'�n������z5@���I*��},4"H��=[�俜��dVM��������z,�����L�	����S����q[pp�_Et�fe���9���y�я--�V�X.V.�]�����Oq �AA����;���%f0w���j����GǇ��E��0�?���RY�u8� ׫1�MMi����������X���M"���
8��:�����w(OQQ^Nz���V��N�A}}}�y��A_!m0����E� �����%e���#��CB{4R��/��}F�
�f}� ��%5EE�����=q�P�E��W">�ĵs�D���iuuu�����OGk�
��D�����Y���&lW���s��>ͬYŁ0V�/��"��I��	{�'�
���H(���o*�^�I�q�QQQ�s\U�I<����
S#�5c�7A�����ϯ$'���;�B��>��5�ׇRA����&�~@����2c���R��6=Z$�"�y��A�r�����^�߉��IJ	*�0	ua��JХt ��/ő8�1�4B�M����l30l&�^�w�ϝ��19�٫��!!!��c(&fg��2\��f`
�llE%%�Ǔ�Xw��1�������?jyB��Ow??1=������I8\���+ɸ6�_����9b��)�:	i�
�\F�c��e55�[�$�� ��O���Դ�����MM����q%E�B���!�Q&���<|��ں��(��輄.��ʪ��e�[~Қ����Q�;��*���B�Fe�����ܓ��[.?2��i�ج��3㹵��Ժ����%���ե��xbA�ֆ�)�js4�������D3�&S�p82R�;���w����6��C{`ek;6)P�![�%�а�i�������9����_�5A�DIu-����wpI�@��2+a�����h�l���a�%�\� �G俵^%ooo�R��Ut�%����)1L�Ǡ����� �=z��G+�Y%��t����T�hSJj`�����}�v���&�o������b��y1�r)p�/�T"�l�7]�B�������(Tl���E����!50��H���|R�-�8�����`9%e'�l��s�����C���� ���=��Do��K��M��+���J����`C9W`��כ9���7�{�K����t^���3=[QV������rۜ��%	~��}�q�b�SJg�]p x��L���l�BTש�I�'z�>����Ӓ0�]��'��A��z}R.vG��Y��<56�6�������Q�R��*+��#sgý���?�D��J�����v����2�~8�fȟ��J�^�Oє�~a�Iǰ�s�^[��kfs�<y�T�C5!K�'˽�Mv���%ǷH���q#�pۭ愅�#ua��O�n� �ډ�����N H�����i�QD����6���h]�<����¤��w�zv�"�n�}��X��o$�DI1�muZ	�#��b����sC��*�gcs�a>	c �a�ɤU��YH���[u�p#yP��q�sr����*��w��k���24�@^
%?̕�dX�����!E���8z���:�d.�TS��%�M29U��֐�AM(���(3E%p�W�2��V&v�[0X� ��m���[� Oێ� �����������!���X+^?~�BI��01Sxt��s����G�:�;/̉K�p����f�_��	����>���:Щ�+1�-+�2	Lq��@�aD8� ���P[B��l���h��R�)|c���<�����B�l�bˊ���(���_�e=��bE>�L��B�%e�`���
y}�Mb>�+H6̠J�u��ZE����/c�+f�l�a�#��g�~d2��
�hl¢����ɐP[��43�K����A�~��)�^$�~0���oss߈AҐ�k0+����j��S��W|�V����Y�$�/�g�!���E��0&2�������+�"k�6yZ	��ѫ������_?��'K��:^��~C��;e��J�D��|��Z&�]���(l�@;��Ӧ����t���/�.�\·p�@VϫD-��?���n���vHb`v��X��'�,[���|�U|�Ö-;~&���N���p�g?q(?��=H�YP��f���Eka������yF�.�_.��N�E�o��:�`�T";Ló�w	�}�5��k��F��x��hz�ߝY�7D_��{u`4EMJ%d���eXEepbz��Ds\����
�oJ�=BG�~�AA���=���l�ծ��?J� �;���B�T���<���G���8����ma�R��B my�-�J������U�Z��[\�f���Y|e?��_�F�U�H�o���oz�+j�����WX9���%�:	��$#�A��))~��dϢp�����5��/d�C��P*�:�}��oV���sL�Nc�VWèf�%Dom��7�E��E�˾�9ZG�Ӹ[�_;KQB���$�O:�9Y�<�W���S�o�3�P�<��iSuG�O\�(o/�c����-�;T%W md1MU�⾚L��%p��g:h΢uXcI��o&���O$�.D��t�2*�:��/P��x �CJV�N#���F���y�mb�r�x����3v����W}W0~�#��<�Wi4��P��ǳ2$�"ĝ"4�������\(�������ҝ���A ���ښ��%+�3!4��Q:�ۉ�-`�S���G�k���A �^����n�R�����ܘl�װ����S��2�W�\�+g�\��ɾ�I�� .���l:^����C�f�EE�|=�ϫP��.ϴ����bɝ�:} ������{ggK&�&�h��n������4�(	N����+%���%���i��7ۙ�RL��	�1�w����-����Kf#ǟ�'�i��J����K�iǓ��\� ��ծ���l({_�1ss}����!:>�9.ڕ�A��~�����\4xd]�DIS��ڙm���'P�\�T[��6�z��o{�J���u���P{���Mv;ԫ�F9N�6�$�#���J�DI�������y!!K?��/e�픥��°P�5�t:�P9Om{���@,��������)�D��·�oiچ�-B�Hk�g�{QPHTfn���4\6N�;"�����ʚ��cTy�Em�t�q{h,��f ���lllB�q���C�PV�Y��X䃄��3P���׉LbiŠ�C�߈]u$��CE���K��S<�ZҨ���X9��q��Դ*��>�
ƜK�ΡU����4�Cv*���U����M +��BQ(�y�&a�t�UC���#���P#3�$�D��)q�H��$"����<��
D;6;�A��af�Uм��ikC�b"@��5�Z�g�	���)�Ǔ%۞Ue��@��e~p��K~�ߛ��L�-�s�x�d4Bű�K�_?�F.=kwK�2��Hn_�*q���O��K�o�������I�ef�|�&���|���x6�U���n�Y��A��xK��g᪩Y�%�TՒ��qi5R�^����aMYރR.#���v�~}�?~�����Z���)Zp�BQ�,�~qY�#�W���^;^���t�L��0�Ȋ��ddVQSYv��<�xN�*o�y"�)���`�;3'��g����2�*vJȨ�^`��O<��p���f<��05� �d���=m��3�a�Q?=�̈́7G�&�J 7hv(�@V������Щ|ѦYQ�[�d�.��X.ޣ4ە��$#������I�d��!0���kqQ��C��M����#gzb9R^:�R�f\���u_@;/�MNKdlz����F?}���pe���<�D�t���O^��g���&AAYAu"{�9Ec��iRϲ�d/{�}ׄ
Ҹ�;���~�(%iC��:x�<Q��㿽�ɀ��i��>}��W$tB�W=��c�3i��f�n��>..nx _�5�/M�b�3�3�ua3Sg~z�z����]A�~g@�W��.O�QBHHV��w�4/x�R�;Ҽ���G�x}33��X��Z�89��Z���͝oy,�x}FٟH��A�?к6�:܈�3�P�r��O-@��ݞ�F~*��8�*��#$<VXcQjٰ��L�Rz��Z>�����d�W0{�|V�uw}�x���:�M�A��A�O�s��P�U���p��S�a9j;��w����O����<�B i����\�ʥ����ˊ���v�q���Ӊ�!L���M��R��A��Pz$.�D���������Kψ�߀yO_Q����K��M%���z�+���<L�^�]�����<Ԗ�Xo�����ǩ�C!$D��Th1�Zڅ�@������2���qc�Õv�tܒC�Q	�[�g�q���Ka������7S�r�h��vm�#b�7ם�q��ؤ�O9�Z���P+����>�/v���.Q�!��9
�<��FM�0�l�Q��LҀ�h��˝��D�)�fw����DQR7+On�ri%)�3�a�Œ�<���̮ʏo~�R�1�6}5FBdI@�(ݛ1��L�G�q����N�A}]H��Z!R2'�o�1�v.���.zw�͢BP�9
�|��"F��o>�W';K��1֎_��9 �32�,r�i$�W��1�_I�9���>z.�NZ��ml\�۞C�ט[�{^�5g���ʙ����WNm3爛�����'����A�c�2&�q�������KM���f,K{b��u5f�f;(v�C��1~9L��\�-ӟ@��`��%�,Rx�u�l�#1.^Y�"^�?E��v��m�����������)�F�NS�����E�A�0�8r
?|yn%m u���W���t<���>����)���ݴN1GQd(�{������@`V�e��� ���EhXx���pR%�`3p��R4���u�M�ƌ���f1N�_���n9T�����"ǡ�|�~m���w�Y����.hvzA�MhL�[�W+:�~�^���ť��K�`6�sLL�ū=�z~<!a!{�sL����+%���Z��F�mYU�{�jC��l=����<�gbP1�E�GI[�o�ER�ߒ,���*�e_L2�bi�t�I$��b��]olƼ�ju��T�t�L�~UGo\}Y�oъ�6_����gU����=��A��}H�־���F�&���i�ݯ�&��(tiH�d�X�U�!H�ТR4t��mi���ܠ� 9�u~;���\���n��t�{���	Ҫ�k����R�#�
��y�q�b-�3��e"��o�:��es�_�� ݍ�:&�Y�>�a��wB�ls�����
V��?�e n��L�L˛2o1}�F��J_��[�''<���pYOffЛ�j�G�u,�� .�����NnYV�5�w��	�'FV�d�$X޲�nV֔���`jֲW��\J��X��tE��hh�3P�m�N
�A-?X���nܳ�R��?U^�WU�m2.���S
&���"����{>j���;QP�|��F�����2>�E���M��v��
�ohؽ�99\ S0��q�1�*�m䕞��}�?*/��.�]=6����#A��%�V���v��ư�J၃��>tJ��9[S��=���)S"���a	J�o��!�)�If�Z��9z��@Sg7���Dfڀ����������ť�=�"KX]-�ȑ<��Z�N�p>��7�y�l)��/��|����?�}a��Ŵ����[ ���"��E)hOVm�`z#�RVq9wpaط�+�Y��*}��� �=���&)�i�J�P�����+��~]�eܤQ��t�wxx8� ��-�L�[Y7W�<�q���G��kN�QR��cc�Z�Ϯ�}�Ĵ�f]؂֡��7�FP��9�GyW�ŬmYa�V���Accrw���~�S����c�[��PX�����Zg=$�\�ʦ��^�h�w�t5��hS}�T�1H�@ ��4v�RQQ�p-�<�D�_�1&�C^Tf��{���jX�x*sߺF-����n��9e��i��/s���
p1���c
E�>���5G۰��R��,��w������8���������!R��P��R��N���W�T&�j lx���&�* 3��B%�&r�����7+�Q���xev�;��+��w���k��c��G�u|�\�2�6��á�c�Z�QKCS�s�ݴ��;7�#�"7��1����v���.À���Z��y4<�/��>��l=!�n-E�ǒs�
��Ε�INN��*�[����v}��kuu�t�zO�,	������𜆻�0�8KJ�����1�g�w�;/���~�s�\L`��
rx�U�7�Z'�'_1����B��ll��nF�g�'Q�`)�4'E�5*r	�Ͻ�m�倵�*���~E�	{v��F��:�W��!����^�V�۝����KD�\ӽ�C�������;	b�;�e��"����L�C\z�c*Zhä����y�zm-�u�]�<�	�[�H��5��_�D״,��	�w����kˡԡ�]���ᇼ�_2ٯt�5�E@�0c~���_1�%��,l�̮�'�����h�)E�i������뚺�]^K�)��zHG�>'�7o(+m��R� �8hI��Oz!�0�������,��b�7��&�Ҋ�,�އ�<[��+rj�%o��<V��q`�g`_tT�׃z��U��wU�{2i�����啷� ������C�I������C�Lg�Q������S���S9�_'�Q��*W-�����|�\��`�A _���� �*]-i� PK   �yX$�:{� � /   images/5dac6161-a6f5-4ffb-b809-ec8007c48853.png��uX�o�?>�BDT�']�#����tJ+)�k` �]���D���s�9ƶ���y?���?��C�w��ٯ�u^�n��U�/0^ �@�O�<�����@��Ν�������~��*	�x��4���o�<��@��I��s,@ "���G�����{$[{�������-���W���߭y�"���'��-N���&L�TW~^U2t��MJB��ĭ���	|����o�<��.W+�-���w�1w�Y(oA���8Nq{Z*L�"S�;J��_��w�j�A�?���G��/u�_$�w����p��?y�3f=�Bw���u��|w�B�\Q�:E�`������IW�����%��;m����ɒ�}oqyک�\{��s�!Ep�;�� 2�����WH����G"y���k��s�<�������9�r��KI`��6���O�
���22Ĵ���z�
��\ϯ���� }*@���zu����a�<I��_��� �ZL;������م��Z�)�a��[|�ׁ�2R��%蓻d> B.���[a�ĺ�eV�}��y)ʧ`�Xi�2�ޠ��Cؑ���#'�Q��п�?��+I��gSV"-�����a�&Z���j\u��!�@a���:�Ɓ(��\�p�������=t�g�������)�aY�o������죏`@��8(
TH�۴kW�h�Kg!����Br灠�PV�5��P'���*�޸�{�v3��H�	9�
���׶�@f<�yJ���$3^���.�4`pV3���仆:��ɺ�'vZ�\ �����9���+�����`���LA��M$)�>�1�r�_0fQ-�~r�?}���gk �����}���Z�d^�h9-dj�����N��Vf#dn�s����^�3�J����e^�}l���%Y��$E/6/�ͩqN���M���6������h=^�p�97{����n3��d�ó��SD��&�D�z-7�S��=9�����Ͼ��2�M,�#��BQ��}j�^�r~��>O_���br����4Q��_h3�x�!��kS2��gQ>�u�J4Fy<��r�q$'��9R��r��g"������X�G?5(�A�����he0�$Y����� �<>e;�ʔ��Y���<VQ�l��\ܴLp+�H�J%���ٱ��7�㈞�\%����,�u�2�!�jq�b	�%{�:�`�D3�L��Mv"ŉN��X��g��%S�P��F֡eW��'N�c}� �� ��m[�:D>B}|:�~ѓ���<s�Z��H۽�)�x���k�E<1E�	��kH!�G6��8d�:g��-���Ŷ܊���q�|:���y_�d��ӂ���lc�}�x!ѽY&�x
B>{	i��v���J�JM��/���e~\(}�F��v.��Mx1[�r��2�F
��Oe�]�B�DZÿ�p����Q�?$� /��ѐ��� n��׌���σQr"���,r��x���g�t��Y�
EV~�@,+�H���P:��_7�&�PLz yi9=$���0��h����(���〾_
��a���@
���:E����=Y�o���I��DeT���H4�D�Ѥ�
2�%S]�����0�p���"S�Er�
xI�W�¹���.3��5�#®|M�D@�3���J��#�:�u%����� ��i��W��i��3;�c��n���FM�Ĝ�c;��(���D�33�gNU9���a�p��Lc�(6���Y9�S����-�/�����V���N8	:�0�Dib0�Pe�Xn$�6��u��:��Np���)Ȼ��{�(�Q�Æ�1[�~eKa�;�K���O�g�K�Rϝ }g W��yYA5'� ~w挷̭n�����V�2|^����q)/�N��K-��:�bv;�*� ��.������h����gth��Q}ê?�u=K�^|�#P��R�Kp�#L;Ɇq��2���H�(�e{U��j~�qF�q]]���)��\���q��$�~��J������z)\y�;��&���4"ح,�������j=7��8�e�|
�����G��H�����l3�ryZv9<�i7e�K*�* 	��R���%c9���3��� ��~�+0�U,Ώ{=J6�����"�m����������S�s�[B�+]��H*�E�@~���_4�f̘%>mL�˒�gǝV3"�HνJ��lg�E�6�e5�4�!=h��-�J�i�q�f�0�1�n�*��e�Ը�v*r������Yd`=H�XӰ�5���B�p��5���[��0ݯ�_�S�/A���C�"(w߆�-TY˛�`H=Q���5��5�Y��_%
�K-Zk^�c.��x��2hn3�48��u8�'��yH
�ܞ����*,�MB�.���o�'P��w;�|�sW���> ���W�+��>%�0����,�m&!�o�?�^a�K��:�B}nӸ���K�	�Xt�!)(�|���6����`�W	pӮ$X��LB��t+^�Q7�Iy�/���c��H�����M�ޔ�L��r�+��m��V�F��S�eV��E��w��'Vj@�$8��$Q��<���6����R��M�n'5�S:�w��Oꪵ`^3��a>�ȼ�X�#qgV!�/�ݛbP��t`�QLwQ���13؏���*D"�=n��v	�u$p�R9�޻Kkٗ�M�e2�׫�27�1��g Hb��Y�}��U;�
+�>D�΍�b�R#3��U����8�i�z�>��(Y�����!e������|�c�NI`	x���p����jm8P��~�&%q���[�ĪP���O���Dl�M�X�ݏu�M�}&�5���F�w����~zd���*�x휀��v�ט4=k:+Ճ�A�c<�H3P"�ģ�
u���a�e���厳DqP�m��� �I���h#q੶TL�2p� �r��յ��!�x�۸⎏��Aoº���/�� :�U)+��8��j;�ufO.>$ǯ-��U��"O>$�=}MX�SF�9��h+������C>SMLg�|�L��I���x(;��XF|g똷Z�^��/�[{�YP�z	��q�	�o�����K�_l"���ޤ��(���e�����E
w�4-�0�C$^' R:h��&������[�$0��YH���J����m�3�e&	�D#��wD.��4c4/�U��|�S[ؓ�E�H>��8O�N0��^���3���D�IV����a�w�N_q���h���v�$ܰ��X�u�G����G<���F����r?�k�>�m�8�Zz�h����1W��%p��,���	 6���w��b��b>�p���<H��
�4���� �"��)ܞ�@̌0G����7fq��􉑋�ʣ�_iGyc
B�C�����'�gW�n�S��Y�c�/ƅ)-L��al4��%_���$S�Iʦ�X!�\_�9�]g���5��Ȫ�K� ᠿ�T �u�>Эh�件΢�"ֆ�>r���a���u�Kh�;�&j
�_�E>��\��VA��l��"Qf��<�RG���qc?��Ľy����0���e��A(p���^��v�m
AcY����Dx�k�Ä�S��#z����)·��6��6�qw���9�%����q8�W��C�窶xj�-�@�}�#ba�6pUj�q��1_l�0��M^�����K1�5��N��&ܔ	f�y�)�P����t�Cw��p��-[?ʹa�����ܕ����e����/���/҇�,�z��OKt9�&(N�ޟ�Zf��d�� 2JEH�C���y��cA�v����9�3�w��U��y���N�/�ME�S�w���?]��,�~4������/�M�.wq���0H��"q9
ݢ�1�潲t�#η��̧on�gw�Ƙ�M� ��3���yr���\�+�s���>�p�х�GL�)�`ۮ��ˀ����fG.��f��Z�ވ�e��Mzc�����f� ���d��,B.>����}�
����j� &�;�"��8}@"��5(��{�\���?��T���e�p`U"��)�8Y�����;�y�пU�fO�̬.]>T�#z�)L=�������1��'���#�C�W��f�<s�i��y�b>I���H�2�'�����2ש$�~q8%f�}z+����ГX�GlqB֪�#�"��*k3�v�������i9=�X��*��g��+��jX*����_����v���6��ލŜy
)��vSV�$ef�d���9�����P`3��n��6���ZJ��A^I$3Iv:A�)��.W�m�(�鬩�/߰#�����1<AQ�k�r����m�vjN��eF6Tu��Q�.7%�a��K�ac@��o$�F�od�m/���6 ��$O���q!�� ]&������p�X�#RH�(N�S��Fީ�����n����v:�]��H�%J��p�4@*$Q"�ء��hhM��~2?pe�F��3�f��_�4뇉R4��.���m�\&%N�h\��KF��'��S�2�H���;N�W�[q��n��=�A�Z��� �/]����-��	��m��E��;#�F�T 2n�Y��s�_�$�;Փ=�F��������%�B	�JEjN0yH����,�"�]:���K��7���)�7x����)�KM���CE6j�B�����>�>�f�����ZZo{�O� J�_6��i�訮�$9f�&	O������+��,�(��q������p�x�B� ~q�d�
�H�<�(�}=rǎ�X�[�Ð,cƈ>=�D����>�*��c�"���Y}����ם�`�S  Q6WXJ�=zYAB�p=9�Y�ˌ�Er)Z��37���W.��:�c�?F}��켙(�]��>�4E�����b��ᐨ�����FGߟ�B�DWbM��[�c&�8A��{S���6�L�|XT�~JÌ1F�鏀(@��)��K���݁�^E&�����9?t�'W0KN8��A�>�B�4^P|@䚏1�i�C��#���hzĸ_���jm�\[{����%�\N����>�^i��sp?\n�%|魸v�}��<��ߦ��I͌�S���v8�#6wVe�pa�k��`���)ЛrU�p ?����BWO?�Be��~�qUdY��������Ӡ�+��Ľ疾X+\2�(
��#���4�6H�j�#�U����\?���l��������S�D��D��o�hޏྛ]�����L�z�>�8�
U�]i�wX#j�@��m�u��g24o����g/Dr';��}�%��7��2]3;��b �D������S#��L��'@��[��V%�ys|�x�U+���x���Zi���>-ڠ;��W�.��Ui�25��{�:"6�� �]fO��{-��b��)G��S_����.�w'D]��s>㽬�@ ��~�۸�李�ZN�5���w?	�����~iP����3�<�gE����H���x������O��:�!ٮ�߻4 qQ~��}sN[����K�\O`���~7���ώ���ꍟ+�Ey��@��9} ��)�x=gd���!Sc�Ϝ ���T�b����f��`��#i� �|���o�M%|'g>�2�l*�8��H�J��_u�!�#{�Cԏ�+}  2Md{г4�*�N�uC�Q�s�  �Ro0�Blgf"�ö�U=Z� (�|�y]�Yw�_�n+�rh��Oכ��<'�uf�*$IݺR�=Ex�
�h�j�{��T�E���%�5�T�v#ss�;GG���q:�Z��lS�`9 ZT��(���c��|}�O0SA����Q_����|;��{��O���*�)�wuś`Ek�D�n��|@o)�A~����� r�����0N��C����=�8���Kԍ�ˇY3�x����X!�>�D2��C��M)��g� �|��% d�d��yL�)#A[���=>$�ۋ���QN��O�9�]�������7	���j����Q�r7�GM�&�V�RΒ���V�>`b�m��3�{9�������Y�+m�8��������}��!�J�J��XJ����W�6�yul�iF�C���܁��ƩZ i�Sr'�F�w�YHxUb��n��)qˮ.DY�;��w���O��z��U�5���^T%A�"yA��v���w��t*��P �x1e	���n��<;=���"��K[�~H�ݥp�@�ܯ��)���"��$�ξ���͓��N��rf�5J��a}w	�c�y��nv5и��S�8�(S����0���kҖ�'k�BF'5�Ho���A���sv+���}�Wo��$c�*�~�;R�j�;#�yv%L�x�B)�-M�WX����>%KQN9�'@E�`x�yj����SZ�GB�i@�� ��GT�&ሽ$��,s���WIؔ��²~������$c�I���l`+��2���c@�ƙ[��X�����b�ZA��gUe<�Zb#̳ub>R�9,���;���[υ}�r61&�u��J�3�J����L�2�����˔�V�\}��l���	`F8m��`�	�oV���_n�{?l�V9L��hsg�A{���O}b��O'>�,D����E>Ǭ�q@�'R���痀�����GΪ����{�,Uv�?N����ˠ||AquK+�VҨ},,P&aZK�Fy��iy]�E���*�J�*1?���v�Z��wp���xt���>E�}3��P�lpB��Y|k�Q�4�
�)������=׆t��W��K8���-A�E��Fn^�'��w����	V�������/S8��)h�W��P疓������o$ohJTm���E��n~�F+d�'��QH}�A���#u ���=��MI��j��GYf/Kpe��O�P]�M���K�-�93��i �H',^��=sU��=5��5V��~o["�Eo,ٱ����/Q	U���0�ǐ�F^`(� XV�W�A��p��Ӷ�i��S#s��������E�'�I�P�o��L'�������6��<TH9���¿�h�����o�E�V�����iG�S�cd[��a*�5�=���`ގ�iX�{�����`�'�m����L�]����P��,0�S�s�=@uB&o���3���i �5���/��y���k'?��Q}��:[Pe�Y�[ҁ�h��X�Ϳ�5Ѩ&�8�y���m�W�"o�\;�(�}���̍��ē��c�~&%芟�(d��,k���<�oʉ-ׅc�&OG��VVY�?Z���y�eLC}6�{%eY��
���iB�+�� �~���4�v]
J�l�I�G��#"&'�'	ߖ��SX>v�)b�ȝ�o��� 	���?��S(C_�{�(>Y��E�=U�C�I���[g�=_�3K������s�}X��D��*���9Q N���P 9�<9)/̮V�]�Ȍ{�C	> ��d'���˯'v{Af�Gݑn����S3\5�Kx0� �"$��
C�0,f�ƙ�������ʟ��_̏q�#��$ �ig�u����9��%����e������=�Sctu���0G����:fi�x,k�Qv�=H<��2����V{�\L�6���];z�n@�{���{�}*\�|8�hj"%�$8&fJ��޹��������{�2��6!zb�R8P]o)����WS���<�z�
������C�6.�a�J)�Y�� V���2����=��t���ݩ&4F�odw���������Nw)j�/<��i\�j�$ ����0I�cC�а�L��Xρ�G�G%�9�J�b�M��$�u1T :���̙���]uB����ό��+�Ů�.�'�]f���x�g7	���0�2'0Z��ԋN�NY�F�w┏	@3�'��(_��:b��>��=�<����!ob�(�lmC˞��R��w����&��=(�'���S�����3�QZ�Q��)�|��	)_z�5�r�$�]���&��-�ζ������嫭(�s3KG ��L0��T��]��!U~�S�]��i�����Ώ�ݸ����K�>�/�~BjF�|���k����I#y�9t��+=)�נ�pY�j�$�}P��,��5�������gkH2���8O:ep��=�����a*$*w�s�+T�8{S���Se�H}b�oLtw}��;�3g�*O���P�'��vLՔi���&.~�M��u�W[>�Ip��Y�1���v�zWkN��7��#
9v�s�������?/�w�G��AM_���S�6�)����� �
��M���L%�6�I{����L�|��n�_o�G_%$At���<��ȹ�:U����ڝ��w
��+
;�p��̈́�-j �F��X庩/<egI���4����ZEJ�����Ӯ�?�{v�%:��ʆ����9�G��<�l��Q��m/��'��)��[/fG��V��j���x٫\�*�X�ݗ~�A����-ib\�2��R���|��Ưױ�!,w��4����Dp�A
�#����%`�򳛸�
6��Z��ʯ����U[��q�v�+'�JK��Svè!w?���Ş�_�.y��5g!$��~�y�Q�W���,=�"$f?�H�i'e�:�/��� *E��Z�i���\���03݃�t?�R���>ab�.��C*:
v��fڭ]�"��ٖt�M�� �(���ҋR���.��:Գ�����]�U�I�@%i���0�vzm,jߋ�Ь-�E�eDK�� �4R̓�|>S+��va>?t�AF���j,A>�/Oʴ?W�Tވt�;���?�43��b�)�Kݑ�B���ܵ�蓴{s�I�JI}���h�',�����L�kP�c�f�-��1�ڿ�+�O����tn!>F1���u\,+���ݗ k��M$���P����\!W���~f��+�f���g��7�}aUb{'��T�m���B��Gho�B�ĝ�"�J ��Yɼ�����M�̛�ߺ���/l�*�^83�nԒ��3w��R"͌�,�_����h3l�'��{���֥K���iu>L]rg7X
��t�����0���=��I�!_���Rmv=Q�3�b�?�x�f���5�V�j�9i�ʤf�1%�W%�hܨ-�1�)��k/A���i�ם�B�At����R4h��&����.�*+%�����H��3�U~;[*;�{ṁ�}��t��E[d,��
:!��ݴ�,��o+���ߌME��ޘ�Yg�'XG	o\��<��4c�q�	��܌�)d���2�^���&�,k�K��&8=;��S���Zֳ�K��3OV��얟?��+�482
��Hx"�%?=��(���h��WS�5%��tp�?���������I����jU��7/X��No��#ʑ��W�#t�i�2��ćHm�j��7�AN��p�>O��/���tx����t5Ɯ�ab��%�t\i��HǙ�_Oyx�*J�|��n�t��{=E�Ee�.kE	}qiy�R�J��T���P����9�3|F�?C�7�ѝ#�����:�!9�W;!�<a��w/���d��a�r��thh2Sώ;�>��/��g:�s���f�8Y�K��yyO��p�0u���e��>���z:>{^[�-�냤|Ѵ5ퟹ5��*����R��:\����4C�,_�ξ�>�ɲ����`\=�T0t��g��7��d��
?vI�,s�"��M�gX�1U�Yr�r��F��Zݬ�zY 	�T�_�'����ʐ�9����}���e�h�8�-%�Y"�7O1op\�ͷg"�2Ri����w���dG{׺hR�3k���^!���c�9;���s�f�d��KPv@yw��2��z����X�i���16�|���gE��{a��#�h�td��!���&�C�O
]���zյ&�����]Z����An��y!���&X�c������[��j�T<�L��2�}6��k�	��w�����|���}z��N/<M�ǘg�Gp��������B�jw +�|��P��zG���ŠMop�H\��wD��o�s�Y}����6��S/$헰��ũ��]�çQ^�p�1ͺk���X+O|������[	�Ko?�k��rM4|a����M:��"�N$�)��Y �j�UH��L���Y]�&�jm�1ߨ���h�-/��	׈hs�\\#Q7�Ŭ�^!�����s��m�7̜rjg�Q{����x���W�M*�����`SE���n�'&��E����s~6ku�|�)��hM��d=T����"���1>��=��եH����We>�4؍�BPu���Q�[&x���a�V^��ȹ�ۨw�6��W�Y�-T�N�*'�:�W{B�C��Q�_��5�`3�4���7�o���9�U��&�6��r�����g��CM�a�y�\�؞_���9d���9s@���\�l�s az_��|�a�/�/4(�����a�X�޽� /W,��c�)_!|(H_X�$��������T�B�+�O�F�m%�X�lx��>zjQ���Y?���ǐ��O�3w�'� �������@r'�h3�>����d��J	�l,l�m��]��d��.�U%��{��e<)�v�s�����z���ʱ}������%j,�l�O��x���؟r�Aҡ2��A��TWa��O�C#}yWL�$��v��� ����p�a���/��-#��Cg%�K\z#@��v{=7ƈ�$u��'��%q�j,(u��j�
�N1q.ziM�nxq�L��`ޫ�ɩ̲Z;K�\�s8肴�2��M�h���d����/i�~26c6�/�,cke�˙��
�]��Q{�W�S-�c��K�w�eZ7�݊������䵳��_H\Xna1/����p��p��u��v�Hczm��c�`Ą.K��m<ʳ���e�d�.�Z��
�d�Z�V�|c��x�E����ː#:e'��/�>@8|�^�8�0m�V�ҹ����3�Z���U݄ha���7-z�@�n8����݉���kl'�gr���ܕ�I���$F.��A��u�|�-�ܦ�DE�5G���\&���ͭ�BE���W%`�j����3�,�<�����/����n�w�x���cl��؅="9Ӗ�<lb��%}���T8j�^Xd���u���6����5��"�s�q��ȜИ�D�Ӣ��b)�����c��e�F�"y���ś4�NDj�ib=��h�a�0�D�����A5g�_�nr�γ��bdG�׻h�Z�b�=,6L���Fxu�\!+cQz���?.=l��Ш��wM����G~ ��Ǔ�^b�|V�~���)�T}�tP1ۨ��/xN�;K�~�� �ϧ`�������g�r�6�Z+�̬ڿ���Z�͌��2�%}�N�N>�p�X�%�SF�No,݈6֗���D�nK�~�����g��HQ�T}+1���"����g��1j�<��Q��:��v�~[���8R�s�G����1uʪq�YFL�3l)in���n�N���DN�?=�2F��2�` 1���>F�%]�b9~�]E� �����+��Sek�\�0UD9F54 �J>���4�ӱA�Q��U��K���Xa<&��>�c�t�=K���> ��OyӹE��>�>qڅ��&�"��C�臸\����)��,�-T���8.L�#�^�v:2!�a-~�s��O,�W~:K@%{�x"Md7��:�	[5O��X<Ȭ��˛��ne{T�%5��O�܅J��R}�dX4=��Q��8V�Dw���>�z�.���ʼ�k��EW�b��6���߷Vo���e�{>��u�Ρ/�n�b��Ѩ��M��YD>i��ong� 㟭�0#6����Jz�*��u�j�������a��ҵ;�����q~y�h��&��-��8q������?mH_��h޺S u�bji��-��?�OLI�~����=�����B���z�o?��[4c��W\Acx��o��̗���-Qő�X1�ܜ��.M�	��;6(����i�����q�=��E���l�eJ��a\'�Ӣ�%^e�e��"g�Rp<�M�����mHa!��OdC7��[Mj�ʶ�y@�96���K��݀��
���������{w�sF$1Rc�뺑ћ ��;/�~<L��"QϜ���rNK��o���������#]�]�n��bBڐ�Z��h��׫����:���zn�<A��9\1�1dʁ�����HK�G�b�Y��Q`��n�ɸ�p�L�J��m5;��9bW�ҝ�;+�ٽ\0�r���:�Zxb�=dT��*�k�Ơ�.��ܖ.�JZD;�[��O��Ugl�HgR�^x�b��Y��Ϋ�Y�0�Ə�X~MG��|�G���j��G��--}�YK}�}�f��B�{�&i�� ����m8B�`��}^Me�v�����"�A�:靍����0�*'̮���*������M�%����`	{֒^Y�#f�|�6��)�4��3��re6~� <R�n��t��f�F󭨨�v�J���9��D�)��^�%*�9�_:W�Dً������|[*\<݈�8+�L�;����u��~�0����8���w�v��S"{���84l�:wQj����Z䝩�ׇ�S �w ����k�܃���iYC�RWa���F�/�֛"|�B4_�~�	�QH�V��.3���O����lĵ�;3N�[a���-x�\�j��6'�\���8k��ʯ�\C ��*s/�ST�yH[E"��E�Ao��]w��U���#���˙�D�:��1�������a�o�]��������Зq& A�t�p�T��E��5q���Ή���|\<2+"��OtX�u�L�(	�����ΙY�G粽u27�jm��������;�x�W�� ���,ç"��ؑ�A0,:�jY�����pS]�\g�X7�X��c�W������rXg}&B
��uJ��[*�e�s1�G�G	Xz�[��J(���Z���b�K��bmT|c:��Y���O����S���Ok�)N�@3?��d`2D<�Q˗1ErľW�,�^ow�f��*I�}P6�]iR������
����mkn'U��Cl}�6��T��#�A���<-��8H��[��$C�R�G���_��Ko�6���HvO%r�9A�"f�~���[ᶦr�i!qG3��
��rH���
2�G���	�'{�0+�k}ʥ�������χs'~'RC�%�܍7�sƘ���z�cks�k턋(�6�=��xPa] {~G�ۘ�,�rct�b��B���0{O��=!�
ȃ� X4*Y#f���q�{"�p|�Nҟ��M�2ݤ�k��B��/��d�=��j�7�+j��!Y��CnY�U6��+'��$�_��Wo��U�1�!��=��]�h��f�ֵ-�����޶z�x�YY,тM��Y��Ʒ�� #m������DȟC��;͸�MQF���}B��GD21Y)�wh:����T�cSJY��������۱��k	�6�a����h=��A�Ǯ��ۙێ��Z.��ٔ��t����o q�r��,v�f`�(�ܾ95..9>쎪`ˏ��"��*�E)���j��JOn�rø����N|��)}���Cx6��R�_�"����k�R�9
e�Gt�v��3�H���8#MFTm���v!���2��fI"bj��}ta���
�K��q��w�h��"��2���\��������]VAX�U�s�="��:o��T\p�8r��d�K7�i�x�ɑ�ԏ<����%-j�~A+�F �VE{+t��>�vϴ��	��j��\r���z����& f��'(9��y�e;X5꫺"�U�G;�ڣfY � lCh�϶мm�.�p�����ݲz_��B.��G�n��];� � �@�;��Aa��Y;�ȋ�,�i�I��P�Eɲ��ԫY��+8���}���DS��U��7|��B��c������ϙ�@����ʕ.D�!f����{�G����g��Z�Z���卣��;���:Y&�%hMO�Ёn&sHߘ��'�ALǻ��_+G�%�7�²�*���n���%@�+�VI9v1ԫ�\�i����� i����\��--[r�ɛ/Ѱr� J�uvzoo%>���q���(�̽Ƌ� ����%�N��ZX���k�\e�Q �k%����(����V�W��=���qk��3�_QZBGR�����^P�˷��"��:,�����LmgF��MJ���'Dۮ����ǡa0*����Xk_\����}y|F��u {��fW�?~�>�2�E�����V}0�i5�7zo�@{��~S����QT�ep��~ɽ��:v�ƚ�t�w�/#SSK��-�n@�:�h�J/���8w>��t�N{j�ژ���ݓ�D�L��H�]=��"qɹ���g�4�w^�����V��n�2�ς����*��
R�~�Y���F�Y�'�!���@���,%�қ��A�C���	ꫪ����_���X��ă�&��/'��>�	�}�cH}��)J�Ȭ��,�n���;Ő�~��wu㪠�C�x,Զ�-����F�s1�G�������9e��6�t������D;��!k^�d��7+=�#Y>�2uJ_�KE
�mJ�_9ᩢ�)�d�UG����-�7��-��t��Ge�V�����bP�q�Jc,��Xɺ���^�II�d���֣�[�\#Q�л.*T�τ��z�SD�����-���V��娜������a[-N�V�{��k��
� �JT��GI�2���܎S�|K�kAu��7��2a�Ήv壺,з�q�\7N��(�$�"�K-����jZC ����'��@��￠_�AB�h~1�q����߶�T�m�>�r���mvwU`.��,JW�Y�}�����7K����U	Χ����C�7� >E
������R�$_�)��@�D�yٗ�����/
\�)�-����4>oa)x�Q���Fh���������O��5�l�������2Z/����R<j��k���W�}n��ǋ}S���;���D�i�b������þ!Gt6����~�K)���J�ғ<�����v�����,����ǡ�ɾ��)9���w�[�pc�3�-U�����_�v9�Yr�Zߓ\���_�F����w�㒏�k(������G_���%�``����Ȍ��ܽ(a�-Nq����N�����f4H����H�V�F��j�vG��;��/TW���I��u�z"�42&�����^:V��g��k{�x�ړ��`���u^����S�GB�����(S:0���d��tv�4�	���nV!D���� L����;����p��V[ɱ�H�+���I3��G3���W����r��FL��.{�f����.��/xe�D���vuY-�a����Z����ٳu�o�1FRG%8��^���8� �=xO(�&���_�,]�^Ep�	��z�}��[\�������ciH.r<��w�b���[�A�|��9��|�[�6.�B8�y�=�泘J;˄�4rwi©�iu��t�.ᴸ5պ�uD��헭�����m�Yԁ
b�>���#�-WA����8�
wfK�tR~�QM����0�ԛ�H^�+���&TUe��z'��Ϳ�ӶS���=O7�~�W��6�G�v>(�&g
��Pm�"Q��id���S�>����)$�M�R��9
��u+�?x���V�R�*;��;�B���%���j��C��+s;<��I��"�2?��W�j�y��:I0���㷊���(.��|�`3���=b�
y�8�ēNU�ǌO��}{�J=f�y9�@G1�1'R�椖v���&k���K��;�]_X�R/y6��|䣕ǋ��(V��'�&
(�r�1�"Z���p4ڈ�:���_4mMǵi~=�[���M�i57�Fi���;�%��o�|����3��zpSK挬'l���̨�++\�L~� �q��ӯ�_8�c�f����۬:��H� ��W�]���N�FX�y�]L3��g�yٝ��v9�z�>WL�P�h��:�l��Tgv��[[6����B�Ӓ�7�w�!jzH���eP�Xr�e���+��*�`��A��!�[SR���b���y�cE��q����@��d棤��8��^�֖f[�GwQ�-�gdk�OP
�>uH�� �[����Z�Ս�����R��|c�$N|�@e{A�}��Tّ��.��i~���s��o�>�`pp�{���T�y��Vh�=!v����J��%�G��8��<�R�߶��_���o�l�8�O�<��^�V����;j0���+�������4���z�7�6�}��H�u� ��A�$����F�E����D�<B����&�[w�qk/�u��'��ʼ�o%a���L��Z�-Iճ/�Tq������U���X�8!u�w���&�O]�'4���7c}�����U��t��j'�AO��w��%�_@NYR�;�$�yU�Da�V�|O�]]BR�A�*GH�.�>�as��5����)�k=��|e�����!uڿ�Qz�t�g�9��Օ�s3����Կ���$�nН:���K����u� ��F��haЍL��o}eC�I�saU7d=���#ԺM���g��i�ơ5����o����,s��AF�<3��UU��ė�7B}뼾�,���_�ט�K�T��X!�1l�~pB�������U�Q�
 �A��A���R��ҵ�,;	��%���u0��Tc�19��P��8��)������Y�__��u�8�����a�DpY-D4r�����IEZQU��LW��R��+�ڡ~�6*>�l�N_xb��}��&����l�2��$��`+��}�XvgC{]Ju�8\�*���ڰ�2�����
x��o��9�~��G�}��2L�{!�2�&_컭̿� )��xD�'�擝wd�@ 
&s^:��r��²����G��Ø������д�����^��-��T�[f�Û*xq�C������r��dM��y�&PF�ճ��8J��Aٻ��{�J���9��ȏ>��u��i��sz��<6��g�uٟW��-�֪d���d-vos3
�|���LGv�j�����uP�!��&�յ�䛿���{~���Ȋ��TJ������x�C�쮹�F����<�ʕ��'m��7tyw�G  m�Ho�\}eXTQ�6 ")(]��!�)��-]� (-�)--ݝ��J70�03���~�{�x]����^kݱ�9�u.�gI�٫�,/@�I_���9q�\���a{��`���*�y !"�8���9@��&���\3���V�y�\�xa�w'��V'��u�}ڎ���%Ú�hr�h	�*�V2|JR�#�m�~A}/��k�D��aK@��/�W����(�Π�
���/N�f���|g�aW)�cg�[��yy��	dPl����+Կ!,��o7�T�z�SW�~�:8���w#��4���*7F�Nى7f�20g[>4�6����2�9�=C6�z�PwƸ�x��	 T�,<Sզ+�жsAgo��Aw��-�EV�!�ڲB��'��=��l�|)b�䙔2(+n?$��~Wa4�N3璁߫�+J�Ҿe3 *.�F�Hӟ�-��@qlK�Ԓ4�5������'�9"���[������ PߋP��p��"-�2%�Û��D�o����eo�A��kbs D jy�ve��N��nᗷB�,��:��^t��	��w	��R>q)8fY�w��B
��@���~*���l����ppv��G|��#G��o���\�\QZ��a��f唚�����,�r[,��<�$걛���Kϊ�V;urۓ/�yL/NV��/�����iƐLϷ�5g����=��W�#�V�
��2�L��ڕ�F�v*�;�,��r���)Gi���jU�}�:>���0lѵY�R�]1S����K�:�c�gӫL�п�s-f�xd>�͛���(d��hNޭ2]��oo�-̾�3��6��� b�Rz���M.�0�Z��x���Ò����b�~��@Y�k;�C���/äȄ�������P|}'q��s=�8�h��D�\�lo��
+��L�wM�mp��qC�0�P�<�?�l	�}V* �V�̅?fd������d-h+�1���NSҒÄ�o�ZT�s+��jf+�ܲp���(	`��<��
�Nd�ӲC-����$�Tʔ+��z� �%�@�:{n�QiV�?H�ȣGN�}$��}G�ꨢ²[����V{��y�ˑwi�]�`�F��)�������SxݸxF���̓����E��@��x�����2m�c��=�����T�=��9ե8bO�F��P���T����K�E�ζ`T�y5�/neRtGQ�_$�BC��K'�`|U\��I�D&�B]�o_��W�{ۍ�߃M'=�=F'�$0O�A{�:�>�ϸ��Ͳ��K6���<"�6�A-�#��ϗk!	g����h���k��?6ޕ��r��_t2�H69W;׈��QK� ���H��ȧ�a�3���h��\ys��5�@�~��Q��F�}e��¶�����ێ�Qq7��њ�1��(�ê���:q'��G��p��Biw��!��J8�$p�{~��n��6�b���y6��U� �R�-��jL8��H��w%�1;9�49ď�	���b������'/���.�v���#�_6�۲��ƚ9��h�R��ן6�c��2y��"����I�1��R���@��qOX_X���2����|ff�r�QM�S��Y�A�kgyA�:9X� 3>��k�h�V���p��\�^d):�[���3�*Y+� ��' ��e��A��~I��)��t�u^��g>��}��0E����{���0ֈ�h46�QF���E��q�==�k�NA�Rn���P8��Nll	���B�\�Όj+��x7q�:.&Y���-NRC
�>4��3Z������:��J6��o�16���)�:��_��@�k:Z ������]�p�4Zu�ѭ���;8~w���;��n�=86��@�׏����Hϯ�l�.��2:����N�o�=lkB�P��y�oz�JMuR<2�[W��LbQ�s�/�������iW�t�Fb�']��͊�7��R+9����"� ��N��ʭY�(���Q#�
��)NJR�{+wN��jx��ox�Ἢ$�8����>�>[�s7y�e��vkX؜�P.H����E1�ԗ~��a��~�V�?���"[f��2;�9
�#�~�v�I��#�>�1.`^WB�u�# 7m�W���$�4�s������j��b\+��O�W�X�!R`���!w���,%��۟ߙ���P���Gs	�s�����:e��~:�O�Nx&m���7YV���>gj�Y�!|"�$F�5x�ya&1�&EÆ�
v�	�,UW���KG-��t7�������hw�������AQ��;(�N��n� �OM�Vr�?vq�����@���A��~釻��0�D�w����鑶E8�*G��{����/zһ�<�+�� �>���lC���>zu�1=��K=b�O0	1ㆇ�V%�N�Ԧ���-�"���Kiy���t�����7�6ò.�-y�0D��l�����I���u�_�� ��d]�v�+�+����|	\�����C�m���p��g"��g�����j�o0��Y3�s+
�XK6���^�O���U��֗"+��c9��.��T�Zl��ө�P/�$������\B��-��h�~��L-d]���#���&d������F��%�Hg��*���� ff�K�8$BDo�CH����D1���$��1��qig�Ux��24��c��L)G�N��H4w�P�\>��p
��J�JO����f��:�{���-E~�Z�ZJP�JOD2�q䈪�ݺ!���1��^	rΚ��ل��ƀ��"/��#ļ�.���ぎ����أ�_Oy4&՛������W�o���[ }3ua)�CnlL�5F�����[�����2���b��2��V��o]�h�uw���|���C�����͌jg=������}�<��r
�;h���#pI�8�h?>�Vf��][��YiMZ��-�Q�����E!�"�����-R��%��{t�� g��({:�wf88���O2��r��l�;���e]<�8�H۪����)�'�d�\g+W�F'��������X�Y7c���M��K�G��N/�5SG_#��.� Ԋw���_� {�7�k�ÿ��}28BI��H����(���3��a<0�R��9���<Pհ��]�j�Z�(|y��ِ��	�Pj/�a�*�ȝ�&z�3�����%6Q�Q+�Z����<�e����\���s=�"E��~���?����{���AӪ���h����!!Oр]��x����� �&���^2o@�5�������S�%�$6ӧ�cr$�;_�h�i��3��.��<���\��Dفs�m�ߛ�aޕj1������G|�-�I��jm�O,]�~�_�jdˬk�k+L�x�}u���|�f@��&�(�%`bEj��/�ԥ�:�c����â�oq�U�����Z��E�(b��w?����p9���56>b���-x� '�mY�� ǣA�D�n����g�{?*�a���0���Q�"����|�Q���w^y�I�2z�;�}(@L���$x���D"�<H����7���D�ŝH�[dx):�lG���Ѩ7���J���B����AK�9������#l��:׊2CUc��D��?u
~ ���D�]�zB�t��9��`������f�+.�<ؚ�o�/��S�Ҫ��P���9$MK����+����v�p\!�*·΋��~���؆B�!�Bx�V���dRr�AL�+�`D@�0����๡�#K����;�+�¸�>A&�p���1'��oSک��v��V�Hr/��P��{���~$E��"��h�*�e;6�C^P;'~y��!��+ҟP��%P4�d���a�@e߰�?��ob_X��(�_#�K����b?��m�����	�Ŷ궓�J{���0ܒg6EC���P~�[y����k�jK}w���t�å��<6\O�u���{+A�tz�z���k���̣�=�EG����K�W�׋hG ��}��QOk�i����I�3v-^뺽�Q�Pz*l�2���x��Q /�c��R��,��RA��J�7�>�{��!?e��c�q�&�]k�q\�u&��ޥW�q:���b�y(����1&hD�Yi�3�U�Xfg�ކ��_����H���W+�W���"��!|���4P�J�N���_�X�)>/��9Z)my�@�/��`�;CҾ��䯩�4P��Xh�f����fῄy)F�~P���i�J8�8���E
T�+b�V�н!8]�P��)��'*����AS��k����O7�H�J�L�7�Ƀ-�s���~ъ�_D6�3���p�$�?�����ɀ?q%QZn��0���]�@�p�xL
�J��,���y�٪&V«@�#>���9���w�$��w�K�e�)h�bM˥�μU.g��6LU���ba��~v�1���+�������s��np:KX���+�YɘZ1��DV�EحS�?u�9mC�P��!1ֳ���nR��VR Y���r=����|S��|8v��&�����c�^%K�H�v��kN-Nh>�U&��0�q.B@�Qc�O����3�)���n����u��.��ՒW���ڸ��Rdp6}O�h�30Վ#<��H]���mzR���h�Eǻ�D~�,�V�w��8L4fԐs��o� ݎ2���
���Q�yq�m��a8}���up����`�n�I���wBw�bO�a�Sj��JCF�1�/V����o�j��������LR�כ\9���Jw���p�>�j�x��!���Cp�! �"�B���O J瓂K�^Ab!B���E��s��R}0f�Y�I��<��H���I:A����W-�"�5�W[1�0"�f89Iښ�����K�U�9"$�>MQ�����@J�
���obD���լROa�l}ӆjK
<u�Ӑ��uY<�kO���X��=���:�̖B�g�jè+�����O3Z #���眱���X��Yb�w�q~�c�Q�(A��R�57��e�Әhp��bi&N����SnI]^���r��Q��#�//ަ�����W#�t�&^_KqQ\��-.�oV�=�*$�Zi�ԑ�%
��]��O����ߊ"��\�#$+W�gg[���jʽ�8������l���n����j��`A}O�T��:��-���Ȁn{�T�8��]-a���ш���q�]��2
z��̾��D�R �Y�+��Ȯ�xG�Ԡ������^\�v����^h=48�(���hVS^�Z�����x�B��C�^_SD�u�M��-Z�_$�ٗ��nU����K��o�/E)��ւsVp�Hf5F5�K
�J��w��v�i��[nE�ʵ���F6��*(Y���S�a��4L���$)� 6���f�!l��x�E�mf�����m��z�����q���|LGG�}mJ0yH��o��0��X{C_��h���$&�tk�Z�+�%;���?�s��iԩ�I���U���
g��a�e�Kh6��xL~��g�;��[3���<�S�m������aO�%�C���]�Ȋ[	}Ө�K���h�<����_'P�m�TP��< aPu�������,5k��%����ͬ�\
�������HŻ����TWD��!nm=��1p �3���/~�'�@~6�.�ܚ]�d������H:@�V��:������1��y�s{	c�KK���in�I�Mf��Z[aa�-��4Aa!ɶ���>�		��
�?I}��+6nD���"���n� J0�P��u�6���$[��a-�[���Go�^���%]�^��ZP�����V� ��Qgnub�Ώp�BsgQ�,C�!)z�W� �uUV��ʻ˖j�U��M���х��+%���ݮ.��zq;�0>�(j��4���O��V;t#6���`;�N>��-��<}�@O5��iP!�k�[a�m�{aq�Ãc�NRs��Xo`�s�B�s�U�p��Q�&4;���?t9��0!ʓ��@V�W�Z����uϧ�"틥"�>��a�vE��v�� �r�B�@W�	h:�~��j{�	�?��R�k�R�h-��ڵm��XE"�뺮��I����e�G�M>���ە�jџV΢��1[�d< <5��m'�*pK��z�"�w���
u�F�p���}l����?�D�>u����6>��	�A��_߻��hZ*�#�����o�(r���\ſ]8i��/hO����L�٢��;�ͳ7�.������<��M����(۽�M%u�n���T"E"��[����o;�V�����_�?��Y�}0��A��J<������x����ݫ�����:�u���G���_�"���e=t`GIy��MK}6h�� ���T���*}�+h*�o�/�.#"�I+�$>@,yY�)Y�T\:k`y�1tvy$^g-͆~K@8�3�x݁ �Ż����B(�����	v�kEH:>ԫﵚ[�yhǙ( ��}�C��[�}��|�I]��v1����a��oDVӱ����������y�#t�FPF ��y�ɂ�@����b��,�����O�}�s�����j���b��%Iǭ���_��5��Du]4�i:=�7l��q��4���䊌���W|���ϞP�sk���v�	S��ZU&�>)����m%@h�1�f����7�*z�~��ef�1;EEy�qB���� |>�>PA9���j�x;�l�u�m�x�KV�Vgk&K�@��۠�0�)���Y�������o�9g��Φz|�~��8_����6Cʋ�b�_�x�1pC�8Mm��x�I^ٴ(@�/�c��?݋� ���?LB�|/@4� �<v��fE}'��C�F�m�?/��M��m��׶�`8�Z/���rH��;�׀�BeJg�Je���g���b<O����h$�z9�>Gp0Vϊ6��V�QH��$32�ڔ&�ڃv�&�}�$E��B��iq�3Á9d��6����7�;�x��ʚ�0���n93~�ꌴgy�,�s�Ǭ9��'c�Ǡ����C,r���L�I+�����%Oؼ~�y�� -&�:j!U��W.�5�l8�z���g�j���d;��t�)�`S �������%�ἷ�o����3���Aݮ'��`=���b2��_R�ӂ���(���ꏗ��tD��N�_&]�{��޶c�Ox3C�h:LkL�_�����pvG��R߃�v��#w�]�T�O��q��v?�w��\�q�K�w�F QjMmjr�Rno�?r/������I����{5��%���*�%E�BT����:;n�a�o�=�P��t ��R�9v_�iV;Xn�ڗ3Y��n3��<���I���vw-�*�����T�9'��U�e�uN	�Jo�+|�"�)&�d��V2F
��;�Wv��|��[!q�~_�ɳ5�<��<���U��!/[׋l��m5:��KU^T�����XxpY�ʱ�7�����s��SV#�#o��u�_8�4�n��%zY�2ːXd%�#��6.������*��X�7c�?�h��ځ���@P�[n" ��o[$�ч{�u��o�?�Sy;E��c&����=���ퟻϿntې0O��1�jJ���C�*
<m��YXI����yn��x{��h���/԰�ۛ+w�+{	�T�V}�_5�W�l�X�u�N,��,b�ƨ����V�ٛk_S��%������j3��{oU� j�ʒ��^��iYJ � �ɢ��#ם�0��p�_�=V�$2�Ş_n�d\���_�/>���5��w�l[²��Cp���m=@ �k_��Hk�`�e��x[c/�ҡ?��-���gC�~��z�����k�F��M,uT�6S?,Aܰ�����Uݵ�b3,�!բ?�!b�K�)��aN"#���-z_x��$�� �.����g�{��8�f2d�S^���9�눹�|q���K��5�K�JS��.Pk��4^U����, �:��^S�b���C=��a�=��eT��SL])t�{/q�M��^�N��t���5������)����L��o���%��AEbǎ:�N��A�m� �.��\k���Y��u��4�L��6����l;����Sx㩻���Bhq�żGӳF3ǖ��v#�Ʒ�y�TX���r��u�^�8�Jr]j_Lz5��C��Fm���F�jC��
#[��4^q��΂���f��bX�?���c��_�S�����0�g����8r0��"pe�8d08M5�~V9Y�$1F˜�b���C�KcWvG��d�Ke>!���e�V>9>��ׅu�k{
F\4�uz��tZҖhyov�s�۷�Š#�s;����$Ȇv��ylk�o9Q��sz��b��#��ybM���e�%*�0zП��ۿ�U�|/p���F�]�I���-J�;y�\��x��Ej��( �#L�5C�7��u��^�`�}{�1>��Wd))�0�ci�ii���.,���H#<�S0ħ�r�t���&��ɻ��x�n� ��F�^/%\M^�IS!�����n#ٿvW��T��ٙ�Iexx�E���\0!ki�ü�[� �L̓0�)�j�x[�i]��9g����;�t�t����ml�It�2�9�E�&��k֒��P�>���rIt�ݹ��NK^>3y�m�«�{E[�!����bgGM��g���W�8�D�~P�b�����B�Y٬]��$䌋�s������aJ��nE�$���` +,�0z�TU�ëߺ�Y&3��JW���:N\�WUw��z�x�?z����-N�ZU��YЌy]FUq �5�ڻ�=B�T��C�͙��n��OӲ�c������^ �*����;c�W-�"����/S|C;�S���1����ֳ�mg2�AT���:ʍ��?z��e�@ο����s��](�v��t(V�`�A��ޛ���(�7�s&�,��.�9��r8\��,�2[�!�V6S�̟[5�y��3�C{}�T�W
!n�S��Q�+�_��d����s�!���oW�z�׆��x^�, �-�8�\#J"w��N�u�A��GK���a�\g��]�����} y��:�R����&#Л�b}(�o.����d�d#�@X��o<{w�Ĉ�L�����N��f4����wY�_@�F��q��TQ|�/T5FU;���^�ڔtW����[����i���	�p������XK_4�m.�P00�]<X�%+���O"fs�i�� � _�:p�
��}�]��0n�i�ŕ��XԢ���_�k�$wF�v�J���MO�T�p�L�\� ɻ'w4y����_?{�*��]�7PP7:�����o�s=;*;*�s �ք�n���{v��S��u)��<�.}d�#Xg,�>,�?��#.^Z�f
���e�a�������E;�Y1Q�.��77��p��Ϸ.QP�]p��H�v��+�����`��6����w�-H-�_�:��tp��W8�s���I'���֗:t7�b����F]�h�w��\u!�}u5���˭ha]����`��F=�
)��*p�0,�5hظh� Whν#�q��m�V4tb������p�垡�	�E�/B�[�Zb��]�q��b�=+K��׆|�w�t�)�A����5��P���M �����+45'n�Z6wQg��Z2�x�G�z���7^(xv�W]�:"R7��O;�]��u+���_ۡ]�:�w���K"<��f��[78���>�A��R9 �{_U��'l�a�)Ax���>v����aT�;��������.f�FW��<j ���+<��=Q�>�N���������j;�r$�W��Fi7a�-
wd�����������rG
�Z�q5�c�C�g�fܸʖ�)h�/�X���p�f�O�<���N�x۶;.��˒ޱNO#�\��~���\y�Uq�&�a��xf����y�6	C]�U����:d�K]a6�M�#%��"�3Q�x����4R-K����MC�h�%T����Ŭ��JP;��d^�`Z4X�/簰¹�_��{���ϯ�'�����!�y�Xm{��?��)�*@��=c����ɕ��ܴ�ẕ��Bja�!�/����;H��e�����uOܚH��͚�d+,v�$ɇ��i'2��3�p�3E<D���Ȥ��-zD�0oٯQf�\�XX�E�Y��������`��?�9H��������O��Ğ��A�^���W�6-i �J	[`o��#�U��٥%qA�b=u�"t"��� ]p��@f8p/�:�>T�I)��1	���b;�f@�0@�i '�w\Lx̬�������j`�F���jRM��^���˞s���u�Fh�`Z?\���k8��GBWu��?��?Q�#�K�����L5A`Ν��G��Y��RȜ�I�
(���޽rN~��Y��6mjn���n�7�5�Կ�Ӑ�%>�0��*.h6~�4�V!���&Z6�X~�v�o����"���>"O��,I��Sb6��u�D��A�+}f��ܩ����Ni�5�ح�ň,�&�g�o���.���A�*�|���A��G�3"~��E���z�%�r*/ld�Nb|�F����k�U�E4�ޟ-5;�>'�G��=D��m�r�gT�����Y���X��2�U`5�*�q2Ϭ� ���_�vM�p�X�x����F�\�69��Ѷ�C��)k٣1s%���I(�9=�M���/|� l���v�oW�и�WQ���_7%���]EWM'X@&F�|d�#��e+%��q��a��99�7��>�d�`o�"^�oP�n״���y�R�ۏ���,,��Ĺ�V���� ��8߆�ޢ���K!W�����O�l�{5x����E4\!��@�h�Vɳ�\��mRK��g���`��9q���V8��:�TCp�
F[��`����툷S&�o�K��u��kpDƹ�h�P�-!�g���a[�Yh�D?�b�ݔ�����Q�o>Vg^���U�B�&.��M�Bu8�'FǐU��N؂���>��-����D�iiE���(�S17��3+������0��gT6�Rn�Qܟw�3�/��kR|FQ���6�l#��z�d&1���R��C�p�6�IA��1�F�OH�K���/���N5d����]<�p�����j��q
OV�f��8��#Cx�-��nO�V��_�a�!�zX;�-�%��w|��%#S3}�C�o���CR>?WA���o�r z;�Q�Bȡ�Ѕ�h4�U�/n �L��^���aH|ߴM�*�7����lR5ki�Ec+�`<��ڿU��S�}Dd��x% � ����8��*Ȇ���F��'����?���z��G�}.~���P����0��34#�j��b	�R�ݝ;?#���Uy��CRˡ?��=}�#:	ʓ� �.�Kݿ/�q6�;�tv�^�r�sLX���d@��X� ���'�[F]"�M�T�s~-�AV/���3�AʍS�_��+��hҔ����(oj��l/7���4#�_������(�c�э��ӊ\����E��#p���Rh§/3��ݿ�H�A��T�W����1g�h^^� ;0�ܭ����;/��=
_���5�J$�yՈ��"��z�]E�L�~:��k�P�!r6���(k2twKI�0P�h�Yr����⽟�{C���#}s�]\���V-	�{�� c��զK	��T��`�=�"����Fn�%�{���v$��d�X\�ym��i��S-��t�����c  �.��S�B7["ZA�/���&����g[� �J$�ݏKx6��0o\t3�,�	z*�RKBɦ�܁B�O"4��N�w����
i�Ck����tO^�},3vy�)��
��Z�*2#zB����ߐ�⇢��4-ב������%ހ���#bߧ�"����ش3�}����f&�+7ב��{�u��b��B�vc�B�|y@��@��ߟ'��b��+�-���d4k�0`�N�'W�r�Wlu�O4��������|Y���`<�������/BO$�-�`r���]���_k���|5U<Z,!�xe$Ҩv7��� ��'\��U�%��V�q<�m[��5�=W+`��В*�-���m �]�,�����0S�٧������+���<D���19T��$�N���t)�^'s�k�!��Ա���Ɂ/��(�W!��7�W���6c��?� ���Y"�::�����h@#�L�q5�.�Ѽ8=iB�i�@%��Z�\v�^b���*;���0�94:�t~��S�\Z�Vcn�<�Y˩���=���o�k��p@F ?�W���~�)����G�@�Ԇ�,��s0*1�R1�H�b�˕�/�LM��]���/�����.Wƽ�-�W쁀d�C@�iĶJ�1��Q�`�o<���60C��2�L�T'!�7������LU{yr%?>x��C���A���2��>+��/Y�(��Ϟͬ:ư�E��Ar��W[3����	@�p��GΕ�7�Ϣ~�K�W�(=U���S�����c|����h�ɒ��F.���·����������M���kV��a�f^7���Pz�"�����PY�ۙ��JЋ��99����0�lDe{<�.���Ud1|Ԫ,���n_=�r�la�.{�PGA�z���#u��!*@������T�s��?�iXӪ����ޱ���lhT
�
���j�`>�$�^�W��chi{��!��)G5�add�LY���G����ַVydG���tg�,?fѬ�h�k�L�Eﳪ��L���HL�\s�g��j��T8l4ۢ�{�.j������g�g�41f�aΈ����>y8�M�ft�kx׍��3��D��fpt�8q"�dL�V,�,�E�����;<�Ló�m����(���=�z*���f�֫��&,4wO�&u5������L�ۺM�^{�d��p�8$=�������k�1�	�}�ry;��\N?l#j��� s#�g�s�Z�X�Oo�/)E���:��A��\�>6qY�`#57)���L�agx������������u�5Y��1�<���՗��2X�~5�����u�)�f���hZ��	�K�e���,=<����p	3� ?M�|x����N]*H*����{8ĨGϨ!z�}ů]�+����`�ĳ}ҦHB�AwWV�ˈ�Z&
�����Y$����1������0�p��0Ɵ*�(�/)���߶���=s�눏�e�@��/n�4�2��e	���[y�D��<$�%�����z�52�o\~�/W���}%=����S��hz�����"�w�B@��j�1_��=Z��<G�-�7�F[��
�ϭ񞽹9�D����fǸ����=���~�̾�� ��'a���͜���}-"*$�l>as�W�C�e[Pw�٠b�L>�'��(��~uD t��8�K�4d�r�ZҲ^|$G*�h��=@�J1�i`?�t�V&R�g|�����W��+
�j[7��h~�_@rU�{a!>�Z"�(��9?�YJ�\.��,�PfE��w89���od^zP��p?��ۼd�k�|�C�Խ���t�ȳi��)�	݀![�VKs�;!���O�m=�jcDM�������Cj�?�Y,ud�s| =�e(���?� �e�����[$�7ّ�R��I�9��(��,��H�z?*T�JG��D��������ꚾ�wn"���7�f�A"��8�^�t� ;AC?;=�Ci�ax�3�(�R�9Y)p���R�V;�<�3��P���	Nĳ�c\�j)�����QK�v;$Qk�����zv���&��_,�i)� 2\��C�W�ݝq�f5:��5#>fp���N��A􆔟$�MTg>�[�^�9�Ì`@�G�j
��>�Yؖ6�r�19�B}Ae[S�x(��I�����g���P����<m�g=Ϫ�R�Aq��з ��bngy�X�I>h�l( %��L}�, ��Y�o��]�z<���,���d��6a�!���������Q���#U\������;W�7�NpNqY����cZ5�K��r��C��V����=��5�o��/�.9��*�'������㯒:l>S�붦���,�j����o���e��ԏ�3�T���Zֶ�g�F�3���v��<�4�U��tw�|�A�ܼ3#I�/���r�R��@���4.S-�4}�w�Z�m.į)��)��x�E��59�/�Re=�hbb_L��u��,���p^9�q_J�/���]��IK��tvæ��R�H�J����[cz�^�*��|��n%p�N����P<q`y����ĆD?���z�T��:�y�h%�Ud�w��P	�Tɞ��,�LQ`��Ѝ+� �}ҁa�P�:������B^EIZ\S��Җ܄���X"Q�G��GTc'U��*3��zz��������<���ܪ��֍�N����(��Xonz�����#^	�'�����뮬�7�*��gr�;���d:�3K�P�]�w-.���8�`�8����B96׆@>Ę�\���zi]Dv�AB
�]�����:�}�ކ���Љ�����O�\�Hϱ�g�2���гӋ��{�D��$v�)��#���\ŋ�����aoϕ4 ��S�t?�2c7��7��Cf=��D��%���GQ���IV�|C���6���!D��L�Z7S�7�v6]ɉ�{���n���!��X5�1�KG5��a���rM�9��;�[�,} ��v��I̙��~�i�g�
U����\§�B��؃e̔[A�%��8jQ���0(�3'6�T#\#��6�|~tQ����|�s4��a�w9��DYP��R�;q�`x�Dc���	�<W��5)���Ǭ2y��<����m�%�EA�H�W��Ͻ�!��}�Tp"�z�W�`o�Rѳl���F����=���A3�Gg���_��R���v�КR�2��v���%��m"�(WL��~{�K�2�Wz��~ЧGmڍR���T�467�0&�o�������g���q$�'�z:,�ϟ�^i��{ۿ�E�h���*� �[> �
�'�YmKMfԎ�Z�kC��H��YY�
0bU5 �A��_�:�(�b��,��ᗎwJj�~S��P����ۧ�킰o"����M(Ǹ���Y��O�sg6M�M��:��{i�`���u�+ʫ�x|����#�~�eh�D����?S���g� TA(��k��Po��\�mH#��A���Ҿ��Y��<d���ˍOR��n�2O�,: �_���g�\��������"�*���Q�P��\��}��WaOP Jw��դ�z�'*�?;�ͣFLv$l5�n��ۃ�?_�"��7B�ɮR��76��?w<&P�Ow3_�Mu�)�8;xC?/v�n7[*�����U�"��I6��z
*9�V�(y��_��_#8D�,g�s�t�M^�����Qx�(./A��n��9:�bOǉ2~c˨d�m�����kJ�g`$�p�S�b�D��*7Hn��,T��HlH71)�$dճ��c�J࣯xFkjʎ쵗�U�$�m��v�k�����՝;��Վ�^y	������{A�ć�-�㕐��[�G�^'�x��7�3����}� _���]�>���K$�/�s�����;ټD�r�8�.R�zÂ�Q�Sf�����S�|b{q�Q���4�a�� G���4Ri���H��qE��`��Rr�D�"*l�%�}�cr�$�E�7{2�����[4���Z�V��'[(�x6�~��s�An4���c�o{�;-��@�h�N���$�o--�҈���P��K�-W�������ۑZ�Ep� ��8�������y>�!�lT���(dȜ�%$ڗ�γ�h�G��}�(�y<�W���^]$K�&¬e�jE)�/���G�I�ﱉ~�����D�s��:z7q�1O^ʻ|LvC�u�<�#�3���>8�����
����Y2A���?:�YDH��Г�@O�����v �iO}/�A�ʠU��ȹ`w/U�%�Ͼޫ�.�U�p�6ЪW����r�l^;n�6�q 枛�:wu�}��yA�zKv%A]�0S�b�i��U{�ię�B��8�?������Z��C �����N�B�!Wҳλ�mn�'��&��߁��YՆbz�X�Tmʶ��b�ޠ7�}}D^j��r �\�Tw�<�b�J+��X�R�R/<Wh���Zzg�����6�-пJޑq��TE}5�U���Z��:#�M��ܭͰ���X���2b���h�Q`@��lꆺk�MT�_;�$	a�ƃ��y?�i��!AX���4���L�\��g�>+#p��r���r�ԗ Fd`��`NP�
�lj��2��L��',_	�@�R��=#*��6�F�ɣ��g^�"�(��̜��1HF��P�_i*�Y�r�@�=��=}q�6.�|��u�D�D���1e�;��7��{1)�r!��=A�Y�{�܊� 7D�({ֶ����bzh(4���u�]�8V�U
A-��uFYA`(��jN�̓IiK&�oe�o	��>��{6iɈLр���!/��6��T[K~��T���|b�'29���+K�K�[@tz���A���I�)�K���(��<��-�Q�y���t8�c��_C����1�����7��j����Bry7�K\�����h"�[Jy�Xf��3���?��V�h����!�]�3��RU"���Ĳ�����X�F��N`?��T3h�!HL\i2�
|_�nU��M�{F��z�,UЃ�l,fo���gk$��|::	_F�����+��P���+�r�ٺ��ճN��8�{#��x�\�Q~o�]�+Kgs�����Ҳk��:��x�����q��aQGM۠�J�4��tw�HIw�t�t�  J	�"�tׂ�twww������|q]��;g���3�-�7�R�g��RH��"�E�T�c�=�	�Qs�/{5HUE,�J�8��oq2�J
|�ɜ���U��
k`V��a�V�O�wwj�'}�v��|QP�pp�>X��?��bN���rQ%���Z����7�1�(�NN��(�+?Y��o��z�W�q�Sj��}|"n��cߵ���k�]�D0�k.�q`s+�?&��w����c�]+�G3���;�87RYt�����68�)�g��5z�$�!;�͌Sg��	jc���^?���qif�q�t�Cj܇0|���;�J�'�,��ʫP�`f8�7�K�i�V34�i٪u�_�ǋs�T3�6��Y�٧��0ʺ�H���YQ�ڋI����h�M)?i���A�$^�HC�L0�'�6��g������V���F�T1��_�)��F�d�
����n�a�#i����7d�8D���9/yU�;(H�n0�t/��L�CZ�2f���x-��o�9g�d]q/������@��+��|���o7~��Zg`0+�Y�������Z}Գ��o��,����z�+55�y���6��0FC	�"Z&9�>V�.O�8d*�$��?�~@��D�+P��N���+�g7����sÜ�3Ҹ	�]-G�n�4,�H�[e�G;}�b�ށ�6W��o��G�UCV��/�U�(6/E��ĝE�Г|�"���5��t����Wxv�l���|���О
��Z{�m'�{A`C%�D�y?V��Q��{it��<q�F�I���s�˾*��,���v٩��T<B�:f�����eV�E�Tm�#��L+X���F�����6��um�񕂓N)�qЃ��� ��LU��K�E`_~�A��ڒC�H��N�-����^a<Ym����� ����dӚ�2�B�e��?��o�̐����
��������NP��1������O":�I�B���6>3�
b՛��:���#]f>s?��ǒ�V�'a�:��κA��O�-nO�>�دP"pg�ۛ����|hO����p��b�+6�E���X^gOD1Oo�F)�� ��7}�e��N'�dd�Ǎ�ώ��i8�C�n�����q_f��o�c��H���7����um+��q-�H�;N�s_�{����_��ݣ���ý�ѻ�T�Ku�z����c8Ӌ��E�]��]N��_^1�x0�ŷ�S@�v���鄮J���K����^�����-�ˠL^����X��?V�̫8�7~�r�R�<0�a�MVv)/s���Y�u����G�ֽ�=9ߐy\0`�]'&S�u{,�d	�:.k�+��<��ڑ'��Ͷ��9�Q^P�PsK�Y�MoVl�EdQ��ˬy�AR�á�����G+�Έ����w4C��h��L��Cϴ�u�-��IP�� u8Ea���+Y�*��w^�w�K"�z��'�-_Mf^�CPEΐ��~~]C��Rͷ�ǉ�g�U�]�n�4�7BRoe�	@j�'���������XDP�C� ��_M�Ù�RD'v-I�I�N}��u3����8�2�����~x��v#2Ŏ�g��P ��^��Q<h��%��i kGf��ͥ9cCJ����XX!@:������=f\=��	����N�N�Ū�{�"��'����]�Z/;�_FWi]e��4���5��,:�L��5�ˎ���}U���.Rn�|��F����$��\Z��dVk����tD���x��������:k��N��S�:GkE:��c{:R�R�צ�������o�*�w��>�a���u2��9�aȽ6�\�H�o�ha�y�!*�R/�����%J�����,�Ҋ,fbF��Ͼ�h6��}}��7�R��K��OԳ����b}̟v��U}�Kc�R*�
	ә���P�����.�1�E��-��4Tf�~����%.O�3��Y�3����Wv� 0�0~b����A�(�z�i2��`<�P��}���!�s>$��觔%�C��f���$���{h���%���_3�o�iR4�F�>��u��g��ꃑF��nW�j.|M����J���.*�!��0|74�=��L�F�T�e\�W�U���<��l*���W%�Pg�H��ɼa	��V���s~3��Ǭ*�,~װ)&+�sB?G=_�HN��X�AZ�����$���|q�!���|���m�W7�	a@�˽��NiR����ȲB_X{!��"��oy.��+F�G�$�)"1������K���� �����:�m��.w����6��/�Au���/(;80urW:����� *��eЈ��'�6͈t�^�C?��P�;_�r->s����q�УV�.��K�S��6��hʊ���Y�z�K8�H�K��{��
}�6	P��ݐ\z��?����eY[�7�tߋ�FU݊���TO�Y'��G�;�`[$���Q���Q_�[X4�v��|B��G@!D���¢�&bS��<�<��yV���T	ys���T]襘�g[+�%+��k`Ԛ쀣�ݱH�條���d�ߴ]|,#���[1s���7��_OY��-8//��;Bw�5à�W�J���wfWT��S��*n�]�S{c;&�*	�c���;Z�"VcQ�0���"_@'�&\�}��'���4/R�rգ-��R4��}������)���BM�&L�$0��,j-�������tUd�w�Eb�mᑑ�/|�z���,r�e�زy�<����B�k�R�ط���{��"t;n-�n���-�G*j��˗�"���_�lKD��j2ƨu��5Z��.���輤&�3�$�0�ɬq]k5�p�7x���֏h����{�+��C{�_B��OʓskM�y>�[<�ֳ}�h�����r��8]5�k���������Ǿo]�<�v��#��W��:��Gϙ<�3�$�53�";(���j-��N%���/�Sʏ��m�%X�QP�nn9RgO~|.�u ��w�:iZ);{q�	��jkCM��>sݬ��h[�r1��(���ی��WI�_o�h��j���Fz��8{[���D��g�{�������jv%�E-`�hٱ>yQ}b�_���GM���֊qf1�Nd���l�sk_^��}�D�\=_���q�t���x��XǇBiω��;�}ߒV��5<+e\Ϩ��]�20�pz!��9�RW>�Z�ca������%
�/ދ�g���r�-�q����ܖ�Y#��!�R���>c�ڃ�Y��Ha�{��&}��fQ��a1kT�U��OI|���{YS���P�6�FOd5_���	��8�cu�X2����2��[ն8I]�97X��yG�E�ˌI�i�7l���:&�2M���u��X�pH�L�k�L���Im��@N]�J.����sP�|�K��e �V�;���2M��i�y��#���ou@+k��u�]�ұd�����ט�q.�;C�SVp�m�־}�͊k����E?�c���������س�;�#8��g���������e[���u�u��(R�H&�.x�Y������k(֍��=�9�~ȩ�/��>M�U�����b'��"Lsj�����x�S|Z���y��"TG�I��^��!�'�@�ԊS��Y �{� H�C2`�H��:�J�k�Ӆ�Q��7c���xr,���_����A�|xռi�g�F��i����q��32j,/:[b��
Q�[���#nX�F.,"ꊕ��%���~�9ˈ�Ƽ�N�!��N���@у;P+� ��(�c)�ɖ��s��_�"i�zzҨry�Ά�M�;�,�>�g�=#�?�u#9H�a��7�ۓ{��
�2����6f�����[Y���TMu�5m�$��%�������Da\��da3��<��S�>�
F��f�ʽ��Ӌ�����Ξ9�Q�0j�=A����:�����ܷ��S�����ؙ�K�|����Ok�C�5��8 �F�X�Y���Nk������%|�Mt�%Oc^_'����_�P������܆@�e�Z���ƒa�*hG0��+4�/|�σj��+��B����ny
�Ҙ�	3>5F�jM(�3
܈�h�l�X��e��r-�_�莽����re��Sq#�i�Af���GL�׮Ӎp%崑��0"��_���Tz�a�	��6���{{���]B�M�Z��8���o��Q@����D�B�c���L9���:%0=zX咄b ]��{�o�o�-�G\ �P�{�/i:�����!�W))0Y�X*�~��b�@�{��1��Z�a|�m�!�j����B�3;�����\�U��y�5d%K�\X�3�0�̨�Z�<f�v0$��WD��D-c�b�ś�go��H�n%+�_�s������7΁F�����zj6C#R��讄vv2�P�hvH>qv�n����ܮ�h-�M@�K�����o���lA��	%�J�7YIzi��j�;�9Z%ď���d��Ͽ�N����7�ڭ�}LAPD���"��!���W��(��]C�Z��NV�[־h���;>�r��K_�{�^��y���<K��}�w�Ha'7����-�J�����Y�L�Z��N��%�'.�PK�m�<M�����hAAq�֮2��6�[�5�CL�L�m,��D��O��G2���'�����@�;U�el�ڵ�����T��9W�zO��c����Y�^_�!lkf+�x����kzC7#��Y����>0�R���M��-��?�b������sd=w�B�ҙ��HԵ�0��;)�v���5�k�1z�X~{��~b�7��'C(��P���,�d���wޟ㏻�F����l�a�x�'��[ݬ��#G�O��Jd����M������d:��X��/�s~D5������:͉��mᖑ:{��\.�\�Ό
u�<�j��S�X��k��"�g�֬2R��,9R�e��/<�������Y���j+�i0�5��ؽ���gъ�K+�o�-��	J���l/����Ķ�r��H�/\����M��p>�tCh�Wʹ�[���M7��p��9Ҕ�2�Ĭ�F�H��5��ϛ$�6Ƞߏ6��e�77��� ��b3�V+�}�QǿOIp�L��i�����*/!�S���|�s�_�"�h���H>�9Z�r�N�|ѕ~z�r�
;�U>��O�s֑�Dˡ �P��%'"���҅[^׋�h,�u�uWRH�tА��!�6}]r|% ����D��2(U��\����hǠ��ys�W��ݝ����� ������Ζ��,���:�%��o��/�I�?$>�H�������S/T�ӛH1���"姳=��TF� ��Y1�̀�����t��2����;A4u5�)y�����t��	B�1^�'�W]��B,�5��	ϋ�Yb�KB0^Mg�����V?����5�D~������ **�
��E�?&'qpf�y�n 7�c����F�S!?l��#�1� !��{v>@dz����}���]fx�w��%��X�u�(k���g}ʱ�g�r!�����`�vq<+��R!�~�$�K��sJ_ګ��"��nve���v����Y��f�{-Ku�x"�s�~s�0�������oF��2��d	D�E����^�b`��8$+�&x����7�Gl{3�̿+�����>l._/{�V��pg���']~l����[_g)Z����������[��(D�H��d�����n�k�BD�{R?h�;G�w�y���`7@��������:!��P�"��v���m�: �#<#݇���y������=�R_�N;)~ɮHH���6�љ҈ydxi,]�au�o&��%o��d�u�j����#_�Ts�>�	2�����޿���g;������o���C��v���;1�*N*�=����n�Y��מ�� 6ߚip���һ�)k�	B�ڱ�r�K2#�c���9�^v��7���3�d�&ϗ.$�X_�c&�nH�ζWH��\R�W֌3uHSWle�x��b�F�F�����'j5(��/{�(�Gh3Cl������DҊ��*ٲ�{�J�6�}�GYn���;O?�ԍ6���)Z+IQ'g|�I�L��־�������z��I�Hh.��-p�5���K��:W"�� �3�~<;������m0`>c"��ߟ�>=�鲂m{G�s~�������[�zH3,=e�u�x�k)?�����V�tK3w˼��/Ր�/UU�I<!��۲F2g,*���="t���t�[R��bq�&�H|%���!��x�c~eMk`�AT�TE��j_� 6��(�;)����I��i�1E	���ǙҠ�`�"�>xL�0>�q`;��n	нI�[[�<��c&�_EMVy�r��*,��j��@��f���c�;�����K2�d��y�ҭ��h�%��їR�"���U�گ����QŎ�ߧ�!�jR��,���W�{G2c��Sv��p��<?��C���&���陫�W4�o�%ћ�m�N��UG� ��%Y�E��|�O��b��Ԙ!��fK>Y1Ǳ��֫��	��R����;{�����6L%��뎒{n�O�B%&Htl�jKm�5�q{kU��Une�T�ʹ���`�O�䆕���wn>�%��f��S�����a��OtG����q���ny�I�%� �/�$#�E%ޡ�i�� ]Ǔ����C�m\N|��3�"�����Y�9�+���,������c��Z�4D�TP�Z�MkVo��`
���'��^�x���x�R)�)�����k��%e�4�]���Y@�D#����������_M?�˂���+$7���{�Y��;{�.�6��%}b0��>�����/�\e����!�'%����i�)�K��B`GM�i�n���>�J���bn��ɤg�m���J��t��u�ۍ�yozRs�-��ؼ�d�4I۟�pm����	c��=�Y	�w�8���}T�m�=֚���47*XP��W.����~h3`��`��k�B��䬧7��،��=#Ja�u����좜�f1h2��`s~�������GlT�U��Fot�Q���l�u24.Q��ż#p���Q}��ۄ�ʡ]Hq4�YR%�꬐���4��	k�VMu���u�A��`���w��z�V��8M�3��oD�
�������
�&fn|0�}j���\���B]+��M�owAk[~�����r#eA�ݠHγ*V�:2|�ZZ�ua�;#���AH�fҺ��A����X�Ϳ~)�vJ!m��#�/����S�+���~�˩��[�!�i+8��603 �<�:4���򅐭���m
��H��/b����-��~�*�v�ik�,-�΍�f���5F���A�/�|��Ni�"���i# �W[�K�/�Z�ͷ���������0���n��V~?�AFˋU�+j�o��)�}��f��h�o�L{��v��\�嫸h����ۅ֎��z¶�%��*T��lz�%k>Lɢ��퇠�V�3�����X*ö�P�aQ�7���Kn�����	~R���r)��T�G��>����Q\�����,������T����Ѣ�e;��,��4�Gg��{ߔglG��as{�.k�����b�/~�L�]���W���h,�ֲ�Nh�j�	5b�^Fŏ:g��}�a�[u���%vbR�o������٧�+��k�Ӣga $�%�u����L��>�<��_�G�H�/��n���c{�im�
qj��p��ΰR���G�D�q?���==�ԁ�?m�O��V���;�t��Ne[��r�0.�;E2)e�g�2.�u�Z��;&���<\Jc8h������4�!������57�"T|�~ �!E\��:Y���������b�7	vC5
���Q/�����>����4��J�3R�B��6��+2�Q״s�4�P����jJ��3�Q�~�DR��d��pmS����U ��u	΂�-��u������o$h��芰�34C��iY���{U��:��n�q=��=L��?^�_	�D��6�6�'Q�������~�}f?�.�m_1���;�XН���y��No}E��g�s�':�P�y��d7W�֙ҫ~qN��(�q�M��{�s� ˽���mo�]A�B�H�@���!x|M�)��u&<F��`j�L�7u�_��N���0֣�̯ْҝ��Ν�i�C,��r�4T�����K<i܆l�)8m0�m"a����pq��A���A��=�+�dݩo�(��H�a��?)'��2BȆ�;�X�y� 0S�&^tʴmr�s��z�g�c��:��gc��z[,���!�*��`�g�j�gM#9!5���J}�<�����y�O�k[�����M�Ϫ!KH��1�ԯ�/5��o�
�7�ځ�ƃ��N�3T��~���͘/>*�w�|�L<�.����:qˬ�Xε.V�8�q4f����a:[���Y��G!=���'�_
�O@�v5D,x�7>q$s�]��G	
Z��★AO(U��s��O�!L��B�������7���N��qqQ�&v��87J~�[�#o����E�8�ޫ�H�^�&D��ZOIN�J��AT�6v�I�ʲ�,�߯q����л��I��}�F
{�̰fd�F��9?"��d,k{�7�DYj�;G.�]��lX�7>�ڲ���'}0z�T��|�1�ʴ7U�Ab_~����}���u�C7�����c_3�3��0�K:����?�����RweZ�w�d�5b�3�aÆg�,=6ȳ��)������zN��!N7��=����}e��9$s.��M�� -(Nd�wZ-��a�\��Yԣs��+�]B卯��Ҕ)� �dFOeY@ �����sV������B��+��݅��|�V�U~�Ee�qׇ�
! JWU��DN2��;?�aCq�m��YP�Y�����d���՚�imQ���z�/���E��脔�i3�yU��@����1Q�!G�0S�H1��g8r�MO����t~K���>j�t��tx��тU$8�T��f9O�h���e�7��G�oP,|F���	d}Ϣ�lN;��ͻ�+��}W%�g��\��̜Ϣ��;#�=	MV���c��c|��́�ܼ@�pS�e �<��#���1�k���[��(/�,4���ZZf��Dp���*�~?��/�g��;�k�ƫ�I���X�f�2|B��W��2-��s9R(Йj�zB�S�4�)���)lkU�7���*?%��p���oa�>bhe����:�jU��u�ꕭ כD�	�e��Q���m~[5���|���Zr��a�"݈b�f��G��`��=�����{F�?RV��1D������7.���զ��Hf%Z��ǃ�%�$�����؅�Ds���I�C^�{�>�q��ܹ�-�����Ј�)o�ʺ��<#f'���]C(�1=f�����J�La"�/��*�`���� �R���Շ'�]�Y�["!������
J��؏���'����a����MoN�_3�L1w�Ҝ�u�X����a�
��Y���V� j�A1�3��"�MCD�ň�V�>����!D��#���G�G�^����E�u�J��L�H*iK��!�����Mwhi�4�G�I��� ���K;��Q�o���m�ţ���TxH��`��V.�������$>zd�~�|�jP��]�£_Rd��tӖ�x?,���>�
��Y����k�x�oL<C�^�V��d�=����,�C"��N-��]^\%�lőe��s�8�k��x�.#=�o�=�_K�Z�Ⱥp�Qj>�2͢K������ޘ#g��u��B.7��+��f�O/&�*I��7��H�j4k��G���xG�K�0����ݓ� ͛����}��+�#���⅕c��M�L:�U��U��U��
%�b~R�2xqف���>����J�*��{����eEh!��<'@~�>����tߔ[fk�/7�/��d03��U}$Հ%���9��}���L����?�|��-1�0�i���\�r�N��^�I�/�
�%���4��k�u��󧢫�'�4\(��c�a��L�������7d_:��'Mk"�̦n"��֑a��U���������e��*J�������`dF�il��pq�=��Ag�gY�[��,��2pKN��n�1C<Ҩ�<P�J���Y��>�"9���9�b�3��IT���Uz��XI�^��8D�rN�L3,����ԕ�*A�o�IPޟQ@����#N���Q �w���p��ιN���-��!Q0�{ 1eGR/����۷��-5���ӺLF�* {�;�?N���
ŋb���i��>��՚����BR릙2c�-��U�e�&+��N����j�s�.
î}lS�YX���7����}nv$W��R�yL�B`·Dto�JvF35�D��?ٖ�U�j:R�Ď��R�׾k�T�.a�Ne#��߿ Y��y����(2�(�8�,<*���w�0�$���C"^y��J}��k��>��`JʛJ�,�o�����T�+�.",�O��H��
�k�T<1@N���Ǚ�� f�Fk�j��w��	��f�N�D��#�����o��fR�i⼥��m峐U:w)�?��qӶ��*F����`�t������_���$�R5���M��[�겯�A��pު�~����I�F��%.8ST���{9�6�ZwJ����wO~�V�鯊���vKP�-$�u�UvR�H1�{NK}��x�O"�@�Q� �{���}N8��5�?��T_!c�_�pf�5�d�%R9zJ	S-��b}K��u��������d~}�S!��H��x��w+�X�0��t�Ͼ���S'�qTJ�u%"YB��0eYz�Q�7H�Wz�>E��T���l�H�c)��Q��ٙ�h-龜�� �����j�[c'���������?���a��'�B-�������5������N!�X�*��c�9�����w��I�!��38 ����Vh��IC�/�.8�;�8� �
ٟ5d���Y:�*�_�\��x�s�������2����e!�Ot��Y�(����d�?�5І��%�I*Y�c>�Fd��/���n��
��_q���ź�ETq�t�dЎ�������^�tgD���%N����f��S?�'�7�
o���z�4�1�Bc���q�B�Vc�p#�@(�RĕK����f/e����w������UV�R디�ŮW���_Jaː�\��ٹ��Z�Q/A�����)��������@�I�l�Oo�HɊQ�٪i��.��邠��E�,�E�e�PT�m:�.k6&�>�%q�W]�1@h�vc�f���69ك� �G��0��s�
�[+\���H�V�K���s��20��X�u�\_e�ѱC��	��8�H����CSm��^�!�j�л@s$��v�T0����j^�����~1e���L�kh1��Ǎ�L9�r9��=�������`��i��u6j�e �dy�jø_3��5C�x���"��dc�4a����?x&(J9�i�3{��i���o������M��L4�֩ɽ��s��:�_�8
 �����\�W��o ƭ�ǝ�$\�n�X4[@B����応S(���{�����(���eM���i%�g1�V��$�aL��V_Y�uE��D�>2.�V�Wy[S��k���p�ܯ�Ֆ�ԺE�6��N� M�Z��l'Z�+��)$/�����C*�.�y\7�����>ꢼ8be���ő��n	h�������O��D�6<�_"gP#X�B��6�(�JmYն3��E*�>XV��	���M��4�A�kF��$��i��/m]��p^�.\�0��Xȋ2o��`]ӛ(��H]nh�v��X��VnW��m�Jp[��~����>���d+ӻw.S�a�a�.@�%������쿯���m�Bh��OY�;���n��|f|�
���5�S�ay���Ž=�;�<ܚQE�������5�񼠜�|>�Z�3p��¢y|�����0�mxc�W��-�0M��ȆQ�^@�#N���a��߶�X��(�'������(���R0�˶ERq
�E�Ե s���X�h I��;}Z���1�߬d�v��z�P@2�
���������rЩ��Մ��Mm[�!�l�%�#y�F��tM��z��\4{��9������j�=(�x?�ץ31t4z"�3�Y�IT�O�m��k�kj�y*rgFE��/�?{������F2#j�㼜J]�a�Ǵf��8�h�'��7�3���V�rOnt[r7;D?M��{}M�ݚ�*LU���L�z���!�1�QVx��(��n����~���DZ������'緐`m�Y�ͫ��]�P�e�$�^Ɖ�1��j�QDT�x8(xD�Ol����N�6�)����f�D�-�;�L���yΒ���f�9#=cu ��*�ͤ��y+�H4�����y�q�ۻ�Vh�):Y�=3�_��<��}I�˨�;�Ш���p���I��m���K��<�-�>�� P8-3����:W([�����m�4a��wp��Mޫ���R¢�"� �fz����+�t��8C?W�W����RР��s�5�`_���͙����W0���������tf#����*�{�ܨ[Аy!�P)_Yo��8ڸ��j��,����8\��� Th����0�i�<�OP����̷�g���ȓO4�o%����-�]}�F�d=�g���~�${[�����G�����c'X{��`���`$d(d �W��o&�L��N�i��:j��k9�S+껖؛��T�OW�L���|/�l���v%��0���������J���M�bd7��g��g+V�7�/v�$�T�Ϻ�(�����ާ��p�"}�/�~�@B�V�z��w��F�x�o��|�� ���h5Psѻ����Z�����-f3����x��:�x��ԡ�h�C����ԄO�f$��{���cW�ku5�m_!��U�����<Ԕ;����D�>/��w�"ݏ���.]�R��#AɃ��]3X�#���yQ`�֕б9�\�e��.��g�F�s�eB�E����Ȣ���EԎ�ǂɜ��k�����TE���զ��f�\�Wd�?̄�="�92ވ*{F2�F+g�R��L�˗as�T�7������>o�ߏ�~_&UW�<���WMx5����F>���do~r��3�����X����*P�ugV���_>���# #��%%7-T���>||© ��q���$ �o�ܜ $�fZ��x��\��Ğ�	^�2Jݘ�݈ݣ��=E0�N ����)�Y>�ʹɘˤ��-h؞�DQy��"�bd3��U��q��b���[�ib�j�e���׏~��Ѭ�}q�������1~�o�í�Ȏ��^t�*�9�'�B�n徒�{�p�$�y֏m���v���������!�Jw��Ɵ�����Kf+zqU�Q��2`S�1���G� �d��(��"8G!��	�pB�"��fg3}��u��utC�w?Ŏ��c����p�	i��@��Yzvbf�~�~ �� �������\za�z5��ϑ�;�\�{�R����j�"ғ�]t,&��uA�5��n�5��w\I5���l.��]�/�E`�sԵ�W�>��*�[H%���$�q�
��n\�P@��;��p���-z�=6>m5z�(����������3q;�WdǷ��%|:-f5<�kEɤ)���/��_
$U[���t��g��E�Ɉ���1`���k��7O���L�#'U8������֝M����}Jؘ �B�ؖ���OG\����
|JlJ����}gE�'ǔ�!�,���}*�G	"����<��ݯO��پ��"Uu�q�>e'�k��ˁ�&��]g;(���A�U"}37��\�Ȥx4x�/�os�����B�*��b#�¸�Qf7�f�(��S�E�`��V��\��|G8�B���f��9D�/�5�0Rs���	|W8sz��'��Ҝ7�&�V.ʸ;�L�xƱ��+����Z.4��d%��5�\4����ѥ����!���j����p}�^��Ư��1,�da7ٰf-O����\XϦ댜�x"
x�D���(��Ё`���$s��)�qq^k.P�9Q�5{�ؑ��e�Ɋ��3H+���0Q����g��V^�7~�ڐ0*���@��y�dAԳ��7�����(j�r�߲n��1w�3o X��K��͞?��g4�&~��Mǳ����a��� ��w����XX��~�Ä�Ъ9��YO� 7��+~��:I�s۷���V�q:^�eU�A7���Ə</�M���F����̈́_���Y��G�),��zSt��E�˜��m�F�Nu1ƭ6�,��: p �t�*��A��"r߃���<�c����ټ(����>�-R,\���.X����V���ڴJ�%�/��B�F�O�պ�yy~�v}�9����ݨ��=ݹp�Y"<�/_��MY.��16TF�Jџg��S�[X�j���-���\��j?����W�aPcMzF�Ym�8���Lm�%K�k����~&m7����$sm9� �9i����0_��aQ�~��S�u���ne��v��W/����m��0�]��+�c��-j���kr��N#v�Ӓ��
��7V\���܆>L����Y�ɉ����{���0$�>
��2�eF�j3>�Ў����O���<lM'��g�aC;�B�s$��I5>��=��MV�Y/���M�ש=~���ԋ���ra��jw�,����_䗍�n�c%��v)������1ʽ�{g�s<����؟�, K}��b�&F>�v�Lvp��3��M&|e��!�yE� �q�^����ֱ�|+�xj���3�)�B�2�k_����&����~#�9-+���0�p赛�ӿ��}�F��Q�8X����!�s�+Lk�78l��( ���q������Xg��FX���<xG�֞j�|�M4��E�0דRrMXn��m�L����5�[o������ޫ����}�f�>e붗KhΒ1ҁ��̹��޽Kg���v�U"��5O�X���Vg���m�#����8:г_�����>!/���z��Q�	i����]]2Ts�⻭�R'	Ӧ�@ۓ����9,�K_���1�g��N8��CPS���(�!��I��9���9��?���X��9��}BC��\f����l�_&�	�5���2���;1 �uq���I�#S��YݬZzE1	e��z+��ȉMH��[��#�n�)��	�X`��ʏc������|4�h��$Ԋ�܈�5�=��څO�-��V�DvR�/����&��.�~l�P����k<����N�/��49����Xu�+�mg=\��fo%�?}s���vY��-wQ��q������]q�_��D/� p��E��g`��p�]��@����1f8(��c�c��Vݮ���r'�xr��i/ֹb�ґIF@3�����/���S�l9�Jz�ae�^��ej;
e�eB�I� 4'����,�F��.������� &�^�%������d�.�U����[�9Ix"��t��
�������B53~�=����a��]�ڷQ������/�+b��x��#_���O������*��pg��F(kz���bҸ��ʪ`p{��� e�
<����!���<$���X���'^c�e�a��|k2�����}��ƓÓO�k���SN��8NF�L��E��P2+����:C�o�{�A���`_YB!f�s�_>=�G�5�iDC ���^�p^1B��p�k�*������^�I:y�q�X�͈�;���O�N6s�ƛ������`�R���YM"��tv'f ����[fc�jggG�<��V��w?�X����P��5��a�)\u�O,����/S�so�͆�H�=k���v�:7�P�|U���d�|#��?���EOD.�4c"�_$(���s-�KoZ��7D`�&����^�þ�ɍ��|�a^@l�������If"}�᪓���q��5�XɊKʁ
ͫ�Oj�OK�_��t�6�,�x�ǂ��(�#���t"X���+g�Z.T00U�E�����c
5�����W�0�|�����I�_����nV��J��	���[��4�<JI�$����ú"�Ȇݶݾ3������|��x9���_�"΅ƚU�V�wJ򾋟%��O���C`3���WQ���i;{�8TB9� �< <��W�*�����3G�u�3y<#��϶���pe��k#����J�"I��
<U�:x p����b(���^���ޝ�"��K�8i����*�j��UaP�￸(Y{)����R���	���G�E������K�cD�\�|�N�
�q�;	@�ǡ8Q�:���� ���P�����,V�G^�^�?�qt�.��.$��{�*~�4j���b�2� ��m��ɋ�	�-�.5F���jw���W��wJhi^�����$p�}�VH[3���F�1�n�}�~��m�Oy�ŞA�:L�����e�\ϲ�X�F�pY���8�iHF���g�8^�N5l􇄇�55�ޤ�<$��5g;�>Z(�3u���������
$��w�Z�䇘���N\Ϯ��0"='�X���I(�ݘ�9c�%Q���G���J�R|��<2�e�4d>�ݣ�������껣����GD�=!A�^#��5� �轎���Dt��(�F��{�Fu�!�������ƺs�=g���9�s�@�G��R𬖉�ۢ<OՏzy=��ZV�`&�3��3�U��>��l�G��8���+Y�45�ѯ>���r�O�Py����u�� M���K�p�ˉ3}�z��9���A����~X.RN����?�l�Q8h������v�ʤ���웺�[�答�Zǆ������Ac�;}�[�N�R7bN.D�B9"/�ZMaqQ�%bWq%�D�UR�C��-�>N�|s����+y�3yˀ�+\9y��ؽ.��J[-�$�N>1ݩI	6J{0��Wү��*͏e^�q) �T�U�\Z�R(�O���*bhǿϹ�}QOH�uF�Ӵ��F�i^d 3�D�$pX�/
֞a���w�sq6�Q.�o��ζ�M�P�����<^�V����yeM|(�<�(R����0)s�:�
Y���p�e�ns!�X ��g�Ϯ��v�coH���M浗�c/v��2�]q�����>yތ 7�R���Z��	h�,�uE��$ͺ�#������6
�|����R
��7�b�D6>�:�$���}8T͑�R*��jw�X�Z�q��g9F"K��P\��ms(�C�go6�)� N=�.=^��1�����[�z�̫v<F.����Ť�!����v���'�B̺��%�ף�1�oB�N�6�;?	8im�!��B���wU���T�n�;�Z?��HCf0=G��pX�؂��Շ0�������e�f�nL��t�		�=ز�K��f��=�52� �]Ԅ�]
�gb�~p�6'@��R`&���a~��]-o�l���=���!^۟�h���)����"=����Ep�bU����Eom�=.�m�\�7�I�?M�[���W#@r�sB�uHn,�O���pw7�x�=Ɩ�i��^12��"�z�[��h!�c�7 ���z3Ȕ��<]�~�W�6G�s�3��R�{4y�uWM-�u��W��c�����{�28o��]V���%n��mH�纺=�2�������T������brB��c�WԪݺ��~���������8a9��5{�6#��mi'A�'{q��+5�7Bv;n4:M��u}��*K����ȿ�	E鵌�􀖃]��v�Q��:�y�y�Z�{���Bm���� �t��ڏ�қ�6r� D"7O���|`�/	����3f��D�=����}g���@��_����s�,��I�k���������Ej��i�[fF<J�H�_�4���d�E��2��i��G�� ��O����J�P�sl��hͦ�/�z`��������}=�^ZǝXg��#��~iA�co�U�LN��l}0�+�Ϊ�_<�s�YSLv��RF~�T��{H�~Eh����b�0�¤l="�ήF�a&w+P��1��_�E��"��fa�&��=�`���-�S�\.(V�h�wz�tnt��ѹ3�"c�aH����˻*�[,j�#������t��f]�W\;$w�G��|��i��:�vh��犐؊)��L���X�&���μ��3�LGFX.�}>M�mߛM�zP�Qĭ�l�}�i2e����7�A����)��yAQ��r۝����R��4b
�Ӏ���_(F\���O���y��柧_`����k2�\�*����]����`���eg8!��Sf�3�6vs����_�I8�N���>u�*ܚ��/.)����qs
�\m�"�����2%���e�'�6�6�Ma�6�ᚖ�=F���F��ѓ1�*��B��"=垲���wN��3:��F�M�����g��gX_��uQ�G����D��=��bFR8�j!���n��龝�ڼ����F\���(�%�x��z^�i�Q��v�E�Yv�	��kc���%���J�1��C����W�D��`��	�{�l�C��k�e���n
�N=9hT�X��A���w�������˻�[�?�x�i�Ժ�Q�#T�jFh?�7,�\�t/~`�s�*�47�KX�S9�/+h�*b�(�r�ɮ���M'�W�R�3q/_�q�$z�Qe+he�l� <k���0��׻��\\����Ғd�F~:LiT4Xx�"�R�S�HqGh͢]kڢg��\��l��т|�|7B�<��>p}��3?�����!TM���l�X���c�v��m!�A�]
�v�:�3'v�B)��6b5\�rIc�����{�2��$<#x�.�9���b	庭@�c�y�F�0�j�NN;=����$�|j�X�)�]���
����B_��t��l���
&�p܁�E����q~]����1 ��ֲy�~�IИ <1�ޱ�TJMp�/,"@�������;6�?�e���o*��P	1��w�"��-���)3�U��\�D�3^M���L	��П.�7p�xzI�^E�p�������\_�'�U�a�d"rc�u�Ye���p�=�-��+Ӂn�\s��2�_�k{K�eT���+�?-�H�uv�;��Aq��{�_LaBd����%vͰ���3��Tu�H	B���=��> Wt���<����W��Os�
�h����x~�O�� _���
�o��
є~�ų�Y���uy����w��&��y]�c�`�(0��;	ϰ)W^�zV�|�Ə!�nSڋY�v_����چ)9.����Shhi���A`-�n�j�<"׏�<vA�G�"�>=7�I,]�C��Ɉs�{�|�Wa�V�KS�h>�/����Ei����j�w{q�c���.�ܲTM2����.��-?����k̻�o�̙�{�(����"NL$��
��N�='�Nj.�~F$4贒�u7� ����<�����S��t��a[����a�A������?�Gj�'S T������y�k-��� v�����+�I�*uFn�dj��,�i��Ƕ-d(v~B7�����l��{�I�SK�G�44���t�viZ�MA	�y�t]��F��su�-�_ͥ=�	Z��¼k��ǔ/o+ր�/�ԝD7�B@xKY6�2 ����)kt|�F��1Vs߭yz�M�>�m��ɐɶ�D	Rt�w;t�u=�Y*!��U//�=��x.�s��M����DOx��%J����_��Zw��D��ɶ^l?a�
��iw��
���м�BƸ�u.�ur�Q��o
$*�ݣbn�c<�7��Fi=�0RE�\���
�9�����P�V[���
q�UY�Jp@/���8r��<ukr�������@z6ʦ��p�'O���#["�����U p�Nٶ�[7	˖.�ܠg �i�G�,`�by%cSꆾ�x��y<�p�VJ�S���%ix0�-'j�7N�O+W��W'_E��$�yz僧���ϟY�m�^��re��~�kM��q�W���ױپ���g�\�ϩ�={�ʦ-	��g�[���8�����D65]1\���틊��"$&7Ek���.��6��RcA�g���� 3g�0�HӐʉ�K��y��1�^mN���UKt��h���[r�����i�1'u���?P{��x�T7m��o�g�'�Yw{�f8wUI���	���;[rx�����d[�3�%O�;i��_)����z��룂��S�T[Y&�ǞU��/a�	�1���Ï�D}V>��⑬ҿo�{��o����ዄ�"˛�.b	W�>��ԫ���Ky�S9�C�4j���EF���cru�u%�aƳ��$y���r�{��ŉ,�}L}��q����� ���󢌺�����x!�7Y�����(��`P�l�w�X��vWޣqd{b�r>$� 	JFZ�T5tF:$N��~���e�ծ�t�{�g),ҫa׎�:��'�Ґ��jcj��nd%�EQ$dn����FE��X#-���J i<����Bzh/II�����d����Q�V�ra}��@S������YB�Va��oӕ����3�m}[����Ⱦ�n�ӳ�Ƀn��^ue(�#�c<+�E ��{K�M�a�+��˿͍	���
�Y/��\	��B~E�]?A�[��
��n;��>��&9ܩ$�-s�=���j�Ie��:��u z��P�� ���^/�o[G��;��'O�ۃf���y�9��}��0%O�5���\X��� <Uǂ��&�6��?7��_7b��0)��>�1J�-�\�S���H��#���fQ�fQ�$Ce�]��-ުQ�G�A��y���+M�����L��̥�	�͙�O��KY���y��͓�x$P�da"��D��{5`s�F�
��X���1�- �j�Q��&W��%�9w~^��k��]}S��{6/�u�J#�[�,�v����'�u�cE�,�6m�ӫ�'�Fo4ܱV%5�_HO���ĴcGY�}Z��ӈ���WgP���6�l]�_�ڧ�kg{�#� �짯,�6|�*��]��$K/c�g��	i(.3�C�f�_��d�"Ae��
�_xd4����ϟ�'@�kS����̉BO�"$��_#�?��I���^�Ttq2�?-p�� t��#i�]{@�v)<MN��3��H�D�S�1�x���L(�<�-U K���/�a	�Z�S�W�d�f�RNt~�S0��9�Y�g�v����,�����a�ڹWß=+=�BvT���/����wǴ#�h��UD�㡱�:�-	v�]	W��	7;O��㬗�j����D��r,٦��$|<��3�c�n݅A������>4^���4�!L�Aݯ\���-:"}�?y\5��/J.��OrY
�-�S��Z�������c�Y�V�R�Q�F~z�v����o�h�h��N�@s��Y͓t�t7Y�(��uz�����Xá�Rx�[V�U�	V��Z�/�"��6���AnR����D�;b�y_x��<8x<(�6?�mݴ��E*���f�)辏�=[��G�j}{ݐ��^AC}�S�����M�-�������䈩AU��￺��W����z㵐Q5.+��i�z�R�zZ�3��Ft���Cñ��D��n#�9��>%m��>c��b�I��w���o�J,tFt�	�n2�Q��j��n��hh��i�j�'F�Apo*��	��Y�I��au���8�z;T���誙)m�'��UO������P��adMϐn!��d����N�gs��pCC�n��8��.�[,�˧0'��~�\I����8/x ��$7�3B���@�sdglI�+Ͱ�_�=���`Ș����c����a��?��4\��e�ZX�J��?��>��sI��7Ή�K��Û��D��#��l�/=�ɰmM��HG��$q�@���
������5�g��3m�_�1�Wc%�'���TH���'�����",�R�B�|u|Q�x�����J���
�\х;Gu��x� �t�ֹ���_=�� Jɔ���.��S<zc���.�y�!YKT��7��X���P�������p����j��,B�-�uu��3�;���t����qhG�F���8i"�����G�Q�Bj�F�s4��ՙ�5�i!��զ����B�6��������cvl���;�='����ܓ
��JEӮ�H��tqQ#�+�W�@eĤ�@�h�q�麛�$�\��4(n��WN�*﫲�p���|����&A��ߙ��8�����+2f5��	Ȫ��]-k��}5و�%�d�e��+JH}s��U �:c_5�p�T�{vN|�������� 0��V����G��x��$�:��N�4X��&o�d~j�M1�N�%���N�����4b �<ϔԜ&�E��Ƅ��<��Y��dU1�h�z��
�n��P���u���������(�l�-L-ӟ����0�~&L���L�~�����/O�� �"��}��g���iBR56�U�6���6�Z��b��Uc��!�F�D1Hh�q7���翪+kO.ꤑ�:�<ʰq����m}Υ��1s£}��C����77��"t��3�KByj�nd^���u�}yi-�_F>�co��j�)��F@���Ps]�L�C���~;ͥK_�[*���3z-�e>9R��pJ�Ņ�z�e&y����!�y�A����l���K&�m�t��*Y��M|ka��ZZ*(�Q](���ng�[�#��#��w��|�T�x��Zwkw��"G9�@G��k�?4��6C�	z3w�xn2n�`���x9t�̕ώ$�U�}�C>\7P�+���u�]E �v��kVD�m��[#�u�~k�D��_}��ʋ�Loh�J�4�����B
Fp����%�wTE\ V<�Q��2����f���Sݟ�l�f�%b(��2�}��oz�� Ʊ��ؕx6���?�I�L��u+C��|��V*��9�2�֩)u]���#�/:�*g-�]���s�h̑z9?q<�2�"^��Ba,����&S�n�l��+��;��b-��J�Y���1���W�̯��W�x�Y�]H#��7���� �n ���\�׼�a3��W�K@�M����^�[|S���/Q�J�6�Y�uv��z�E�C�6��U��9��-��}����:��,�bz�#���l�2���v�'�?�˱ n��KK�q�^$AP�&�:�#���p���t*�������~�<��RT�MSB�#��\��a��O'�W����_��>q+�8�fHr9�~D��-1�<Q��P�������Wsϲ=W�2h�%�&�h��={极�w�L�,��n7��x5Ĩ�/���V�|�.ԟ��?@�*�E���uv���T�,��a�GH�J�^������&q4$�g�~��]�L1�@l{�́ T"l�S<��2Xgy��H����^)�k����ibR���a3Epr�{A�~pk�pm�&>�����SϏ�k}��y��9?�`�aL�^oT���K��4��C���Lr|����P��Gq�����y����>�+-<v���S��r�p�y����s&J5ޠ�.>�=��g�jZ��3����P��M��'�2�6���4�3��1a��L��]�~"*�l2r�8���� �JOO{v����l����օ�4� �T�l����y̺	M�<r�?gky�y��!���DO��Y�G����_�ӧݏ�?/�%ivF5Y)E	f��V`�S#�(ۋ�9x�\ӳP-�O}r��eq�v��x����~���t�pv���yDR��y$�����I&2�"j��|�)w��.��l$3I`i�:{M�ㅂ����J�/�~��J����G����=�D�E�|_�[�����'������q)�y5�k@Y��^�������(�FO�~��<XL���	q��������P�`��8AHv�ݒ�P�s��n�������/b��5S��ꞅ���
��b�9ۉoܚ���,�5i��b������2�FYsC:Bav`��� �Ҿ��"!awE�"�����z��?��W����Rxd�}
���9l݋��{P���,5�;2��<��6{:z�\$��NJ㑫�TZ��UABl����.�̺�F�sX-+�ί�	�?Ff�m��������F�i�e*Qhشi����.��B/7`���L{z'�1��hd����7�p�]Oz��s=�Z5�G�*�F����H�0s<o�M��i"Tv�t!1����>���N��IN������e1|�Z�K�%㶙�`"<�$d���-EOl6�/~���Z��<�!����*���
-] ��ۊv���5���I_��T�ۇ�=���E�OVh6g�O݈�R��^G��(!�������Oi�(�����*^�A�_�)�[Bi�o?4׿��(b������k��şQJU�s�@����`�9�V�!?Pqӳ�2DS>�XLa?�#
{5����P��qh-��>��)��g�l�*�������%AЫ���	;�vVP��Nx�C��gd�ֿ�ּ\�}#,j`����Q�K�x[��,k]a�O7B�!������*���9K*7/��uX�z��q=�Q��Ҿ�����SU���f0Dg��㣔��ɁOfr����;���;A�C��Gf��@:!�� 	�%e����vԮ��L��P��\�]�0��P$��a;Qk�lm/x����[O�ڹ��Ş�x;cR��~H�M�?��?<k��M�mD���/,�h���W/�
!-~w����+ޟn[0���~;t�6�:�K(�?�y�8�]Bn���<��z]�?XWrBZ<�4tL@��<��1�BD��ׇ��o��R�9�¤�֧��n�B�Q�#�{IY_�,��i?��2��Ŵ��f���#��®��=����r��o�CXUS�nA� ����"��R��j;���[��Mw�+E��A�_!��p����1lv/�YD���%ڶl������}��g��f!h�O#����?a�ӱ�z��{���J�#H�h����d{ZZExSM��U�vC�'r����?�<��oTH!��ʾ&�G򼊜6�J5��(7a�5tfD�{�q����v0/V�B�*��Bh�'BX�X& �y��?���w6	�2lB7���I�ׄ��«���o*Bvi���������MWK�=m앳]g�ߞfրB|�%�&��1<d�Ґ�	�Q}�b����A��!�6n��+E�$����7�<��ӣ ��3�7�Σ�� ��	�Y>��UV%�U� xn6�'_j(�������"k����z�$&��kk&a�l����/�R��6���ڻ����٧ߕd�˃�!g90(�� �/yH���
E#�;<�s��:�-���1� �ڂ�8�%������D�N���t`��p���n!"n(5NV���K���Q������-�i�)���XCʿ��F�<�[�&t�v��&�},��+$ ��[X�dI:~h�]���۞	>��j�q�h�z8�8�0�͜!vH���r��7al��ϭ�$>j�U{aD���(kwE'�������\v�P�'č�o���LYe IQc ��Bp
�9u� ���u�|>�3%7I�v�[p5Q٘gZ��w)+�
Rx�T�W���R�������$����K]\�gT��B>u�v�Ju���̭������nh�}EŔ����G=��#� ~Է9r�%�E ���9d����ʽ� +M����.���L=����X���vo���cѢ(�^��֛�3s��͋��l�7�o�@ٵ����	�1��1�<�AT2n���`܅t�r*���#��޹�Գ�jlB� @�M�� �)}U
@1`���Fi7�g�`���-.m�γU#��͍uT��X��A�x�Z�զzmV0c�،��[_�����z�0�G1N�^u�ьB�:I���  �p9�7����m�� ��W̺�/︉���}�/��������n���0#�C�9"�8�!�:�i�K���}�{��I��RW��M�Aˋ�7�?�.\ Iq��o�V�ᛟQ)8+���b͋B��@�5��F�	� ��y����@�1b�h�?m.}7�q�:-����9��>��I^���Y��
�B�v|	�?p��tJ!�����I�GPA8E�i����z�����{�ч��FcS���D��x'Ei#�R� �C�3D��6@����|�	ں����26_���ɘ]�􆟦ȼ������:�ob='���zs�o���?�.uy{*�Q�k�]��|�dR�g%�k��:s�o�w�Q"�2�"[�U�y1&�5�����Lڜީ%Zn|�&�|�����D�����LҴ绍�~���V_��00�4�����Nf�� ��������V�莵���z��,����`������lJ�pa�;�rO�G9$� x Q��:ֳ�j�Mh�ojh��_n?ݐLLB��>�X1�m�!���_���0ۓ�-��8��΀�He�آ�Ԟ�����H'Wt�i�(�c��cWi�eC|`u���������m�|�]�y�AH҂
	��Hj�X���������.��YO"D���p��:+����*��Q�W^�9�`��P�;u_4q5�"e�+���,ټX[����1���ئr�gOٌ��%�`�����h������3�B�ȣ�� [�r��� ���gF�����$4@Cܚ���pWP�<5p�:�k�w�����t$�,_�OD��'D��a����K�`��<S:�V7�
��p��8�T�I��eU�n*-�6ڰ�����.6�����2�ۥ&?��蕐6�z��G�}v�b4�Py����,�cD*E=�c���z~k�!o��J���8�|�����������>���ߟv[�ZNcL�ζ�2�6m�Վ����3�O��hˌMT�e�楧=Ut�g�.�����FH/�7��a��%�r��1��͂BD N $9�gĹ�?����W��^��cϻ�XR�i�e���KȦXyץ��}�Y?�6���J�>�H�"�R�����ܧ�V^rx&1�I�g_���1�j�b���Jw(�u�@S/e�缕(�͖&�3h$��`�BY�0�	�w�p�d�̯\�u=� p{+��	���k}������^Y�DB�w��]6�*�} v���c���6�"�2��ϰ;��1j���X��p�d���6�WK�I��Z�r_���~�L��>n�M5SA��a�U�����o��8�D]T6_Ga�`�&�&W�7� �0kZF{l� �R��d��q*��ޢV_߄x�L^A]X�+�Z�0��j�I	��D��uUI��6�Xv1�摂�,6��Oh��L)��Ճ��ٷo�h�a�Mf���Ef7��߳o~
Rp���r?�u�-�A��1�a����Sʀ���G5�����S0�r�+?�CO�k��:����உQ�]��&C�"N�#{�J�M�����xj+3!k;�	���IF���o�Hʈ��E����i�g(k:"h�S`�OO��W�Ȥ���%P�f@��ڢ[!賾���mP���Bl����Sڶ9s��̰+}y����&���cK��r�9NNa�1�x����#��#���$�t^&(��V���i@���\�8[�>���>yv!��t��gZ�:�۸�k^�D�S�\ a��:�����vՄ��e;DȂB�$-�=��e%��r+��6���tV�yg�����9��u]$D|��ڼ��j�^�"ǜLԊ�?ʆ6p�����r�sT���`���l���!�%�6k��D����ۤ�89%��'栗ƵL��������"i㔘z��%,�p���m�4Ib��^P�&�G�/�vLT<1B`n('�|����CP��D�+x�{�z�<?F|ȟ3������2�i.N�qi��`�#�t�D�mQ�	�\�q�]=�xpay�?�c���V�����=�h���jW������QQXP�ή�����B�W������B��b�.�����8�N�PǬ���Qмt}�V*��2!�qJ�}���OV�A�w��G\�8���?�86�IQl_�P�Wsj�A�&zV>ʯ��[22�c���
�� �p�]�4��Xn��8Q3S�x�Nz]0�z[�S�@���a��H�}ĭ)H���v��7����qbX��ז�m�[�X5<���]�~R������G�n���~��.QMVa9�����4�6���.S����>c���>0��Gd��:�(��鯷{��Z�^Z���4�Cs\�d�0Y����������ب�����]}׈�=���:TAPR���C����r��w?J�x,�&\��<�g�M�ƟH	l~(ơ���)�3~����4c�G��n�ح��zzb�p��u��P��z)q�f~%1!*)"�T���\\�$)�8\��S�Q�.�jp����s!�� i��c�2������Xx�X�ø�ۣ�$�nֻ����0��k�(�E���o�Dti�p��Ti~Z���V�o���VL�v;W;�V�a�-D)�Ѕ"V�_=T}�-A�B@'dPmp�����m#���&4�e诐{:���E6��E^�f3����4���fJ��y�O���ggZ��9�Ay[�ɏi,��mj�K4�p��h���,6�z]���W-�s�8w���=�Ssp�tw$^N��� �D+e����+����k�[]u%�z
�0�1A�EE_$�e���I�n�ʸD��1���C���L4�WdѾX}����'=*�&�F�F+#+��p(3@$��3�bb�<k9��,[����^�CL�2h+n�a��&��[�x�����M/e�-.sv+�vZ���7��	�.���T��B���S,G�j>1g�5���H�EsݰT9+��q�L�h�v�����	j|��[b���	c�Ĉ֣H	�,=8��~�J[c!N9�R|�m���n.�_��0�"�؅��I5�a"]+9���娬��z�P�S����C1l�ڝ+ѯ�dǧ�QWtַ�*��AQ��OX)a�]f���~��F�ŀ�@�H~,�Tf�K��-�8&����{j��;�oL�zW�F�ؗF^B�<§����1��pԲ�P�>t���_�Ȍ'>�?�^&f�_��]�:-�� Ȏ�%Y5��~*���'��I�x��s� �m���t�N����M��B�{n\|�ag꺈�n*�=�`������Ū�dG'�@�H|�w1JF��V>�W�n����R� �VڜC�$�<�e\��|ZZ��	���-&(�).�d��qeY�J��][2��p���|��ˋ����un4Q�K�I�bA�^bJѲ{�*����)��41T�V��FrY@�35������vOע#/{����*kB����d���S s~jr�t1v_�Дi"�Ϟ��'���P�g5�^����T���Ӽ���>t��y���_���U���Z�vD;.ӳ�I�ۮ�06;Zc�A��7��/M�6��Q;W�V�)�̪T۹t�g�m��\T~t9x�T�B�g%���."�6%���|	�[^B7�Ex�<+U⚢������a�g�GdUK�O�3
�|���*_\y=�i�]�{�7&L���EȒ}��&f�>=#��\J�R���$��U!7��"�ؓ:�ͱGB�'=J0G{��S�<g����ۃ�c��MӤK��Г����n�N�u��DB;���k8s�;�V��m�����P��k�x$=w~����<�x�R8�̢�2��B�zOE���F��iI�iݛ��Wf�X\���P���_�JR��G|y�C�;m�>G?	�c�v�h-��<�����WR�&o��]\=y(�&%�5����̽�Yfrp/�.��>n�������]�U	/�خW��0�K7W^b����>	�%3�\�G��e�����_��8})m0i��yx3��5C�9�h�^40�Ao�&��o���h}���������9�����͕���������� �oy[�?51/����l.b����9;7*��&C\n[ �����w�`�7���fME����%���G��8���+�`��գ+����!�c��֬�D��lޒ{q��`��&�S��f��D�������9s$@�"4jЛ/H�V%x[I�K"��-B��W��c�>�ʏ��'P����-�5;��K?�����qk@��1��O��U<�I��?QH���7^u4.ӗ�
G��jnw�����}u_A��A�8t���~�}�V��zӞܛ�՛� ���\����Li*��A��  ������0�"	�aЅ��5�A_�q\���W\i����'9/4m�e�	}�fz(ĝ�C�"�
����1c�a�~��
����S�^��=l8��a��'�U��#@^{^�����^ ���� ��7+�ƻ�u$c�(�!s �Y�<|k��vĊ����V�RIM�H��Md�ĈO|�`&El�Ɠ.��wER#~>�/��M6��0��
-L��T����}�J��<��w��s=�;���o��%�n�q$�AgϘ"��2��׿Qh�ј�ǌ��Rv5Fͦ��=M���u�8C^�������Q�z�Fe6��>b����	1���:�C�k(xr��"{�O�ΨŔ$�d/i��|'!/ًT*�`&a�1�(�& �g�<tI�C�%��(p]u1Iٟ��<p�I�(��m`����f23�K��I��p�Jj�Ix���y�����wFt榆T�֠�]ǯ��2p��%�A�P����`=��h錁'��{'�I�b��\�]x3���l���G��t�)���S�"�_�F�TE�&�+~ٗ�v��PX��e��uP?B)�HlD���,��)�m�{Q��h���r�>�P��X�5k����M��)������r�6X��u�Iq+�U����H�yMO�:��"=8�x����=�&,��Q����x���S\��"ձ�s;�4�`�%c��!iJ�y�-/������iA�տ��~���p�O{��V/j��|��(f+�)S�u3��h���<��ͷuט~^�Pf�<�]&���t�P�����&���'���E��o�(o�(ש�����6��ϔ2��	b6-ch�� ��Wu�`�>z���k�a��0��'�y�M�B����x�9�(�S�\�xUU�R,�?ѠO�pJ�t�j�S��m�YL��±����؁��L�v�ݎJ��NP!;�{�?�~P��ڂ���[���by��Z�mU����,Qoɼ7.!\��f��j�!�Jm�L�!�ԓ�Q�%���cB�7�����C�ſ�'�8 +�-#�	/���'�]�ذ&'���l��Ϧ<��g��s�qZw���e���N���f�:!�c@��R|$���Q��S�D`C�JP�Xd��O���!����|�W�}�x7�&A�#2��V���� |U�4�
����g��`*4gv�C��/6�#~���<�']8����HZ���#������e��y���{��G0j��Q�Y;k�[P��C��))�b62:AZ�^C�G�wv=�B#��M�'��Y�o@@��[
׌I`F�e@��b�l������������/P�����-r�� #�3��������˧ңIk2R��%�ù��?��;���N�D�o�:�(��v��w��a����H�<�!��^
����Ę�W�P���4��8٬����<ޥ������
�iD�\�_��N+֣)I���3gd��㩲-�m�4�-泰�߅�o�� "���ÎB��qNj)�ǂ+��V�5t̻��0P��|0B�E�y���Z׃N]Pm
},"j�?��U��D�p���P�J����-"��\t|�{��'�.RZ��<���P]#JeT)Z��x�bO*Խ�=1���?�/u����������ۆ�W�X�4 p�� v?�y3���t��gЊY&�M�_�K��9{m>�s�&�T��爛^���i�nz�7],��O�di&ʾ����������+��Z��z5	��y����_Zdh<ۯ|5�;T����������`�du��z�߻�qws5���������!��`�~�I|���"!7��i<���|��0ܳ�-���Y�ʻ�wzMwy&��������~_
%_��y�tK�|(���J$��M*�/l����G�mq�[��#�z.-�⃗�~-V�W�,+΁b2��Sn��(�ޏ�&`rRB��2l���6�asꃾ����D���_��{�a2eN.�����]��(5���&�5?�w�?�z�,ⅸ�z��՝���A����uQ�f�-�L{�yĬ����s�ym��y�^$xn���h�1�(�\�&֋l�/��ɻ��|#p���
Yy�Ϳ��dk�$4�t�H`Ԝ��0#�˚�ј�^��5T8��(�u(�vN/��\'�+dNsZ��bLeqcZ�'��=�a�6 `��n�O�[$0��I�H�Gx~~D�k��i�KZ����K"�mȅ�/��C#�^P��.��8�'(Vnn5"b.�+�I�5ԜJ//�W�$�̺�}v�6%-����g�Q��&�fo�I��ġ��k��Jm��P#?W./N�Iy�X�+�jQ��>��i�"�`�������b��=c��e*Ģ�<*�g��{��7v�Hd��PG�P�_u��U�`���f_�}K_�(� B�	ԝh�x�Fџf>=�T��C�CZJ��{�c
rT�oN����J�7BZ�LB�]�ŝJ�>��ۢ�nۼ��A��q�gyφJy�fʔ��w����S� �����R����4/�Jq&5��v� ��ƻ���d'bT�ec�x�T5)1/��|���^^�3r����:�5�P�x����Kz������u[�d}�j�G� �ۋlZ�!�OPc:��;��
%I��d/��z��A6����>��an*
��#V47"�����->�*j�p۞�Y��l�ރK�P��i ��EYv&!���D�y���vqq�Kq�7o~�c�Uo]o��p}Yk�M�Q=��ڨ B����_�?z2�s����c�R�%��M�|%ښ��;�Y�(G�I�mH��x��s�`���/�jH8�[>�G������U6�j�^�&�s�V�����Ki��4Ë��K��ڥ.;d��0�ٚ Q��&p�b����JtMD����#�ܮ���-���.��2���������)�h����M���̻���}��׬js�DTq��SLKh���1�T��	���������~�v�iۡT���jE^!�O�x2�d>�1CDI�>�?]���@�Z�K���>�]�%�V�D�&Ϫ^�2��˘ϵ���:oq!�Л�΋����I����M���e&E=��f��}5H��|Aauu���0�nD,���{�V4�,c%>��Q�?��:,
&j�KH�J�H��t���HI�ҠtK7���H-��%�t-�tǲ�.��}��'��3g��ϙٙE�$C��3�Z��E��T%$�T�����a3�Ґ���m.����M�pV#�p��o���	��﫳����.�ES�P���4N�Q;��_&i��K��{]qU�Y�y���T���C�:�57��{m1䮴�e#� ]+�R��t�F
�!�9��N<�| G��ur��B�BR`��`�BЖW8)�bn|{�9�~V�ߐ��ׄ�]Ĺ���п7�����g���=~-�P�*�32�t\����yr�^���%p@l3��z�l2�x�p�v���� *��ĬW3囘cFM��^8q����Z[R;_7'�5���Z;:�+��3V���DLp�;M����dZ�#xQ����嚴�e�8#;���}�nJ��	8�qb^�i^���}��=���b�#�Ŀ�C��we�}i6����%eOrΫL�*�3�Mj�\»�P���[vk-�'���Y8齺���D��2��eV��,AZj/�l�����?z�n�㮜��'��U�s
�V�~���R��:���g[{��*�������x�d�N賺�e�͢�h���L��i��{S�!����~��%��]�v_�3"�[�{a._���_ν�˻{Z���)�P�8��D��^�	�Q8s�<�N�-/��Ɇ��%��D�8��G\;Ȅ�r�}���,�,8wF���j$A'�2?�L9�F���FE!}v��Q�c�N��; �tV��Qb��OR����Q��<���jN���J�}�'>�q�Y"F)ȩf����Gz���J#����FD;�!���o jM������u���_�b�n��m�}��䮜	�h���f�ٕrUQ"�"�l\�v��޻�%Il�5,�ve�vՠ�F����okq�:��Gp��Y����A,���V棣�DbFf��CC�J�b$DK�Lڲ�62���:<?N`h� �pt�<��Jw�a���~�h[zB�cЇۉSCnXځ�l��)�B�'��L�-q�{Q~��#E9�n��߫u�������I�n��dn���~�{eN@Q�m�q7�c��¼}�����߹��u�
;�l~�`*/�-�}�c� 	�ײoue�@�@k.��x�D�?���mV��Z:�{���S��ee�dm�K��G?�m�Ɛ5¤��)n����b�g��r��\'����k��3D�ҕ�1�H�8rK�����]��F���'H��}my:ʴ������b^�&�O�	԰��_n�aPC��j��V��8Moڎ��B�Vſ/+	�M��31)3' �`��q� �Msߑ��h�Hq`�R�^l�"��A±~TJqe6揸�%.A���4�=���2��|KS	.���X�ˊ���*xhY1|�U�ݰ�I#f��7�w?}S��1.7�3��Z�%�dRN��ɑ��EZ?c[�����;�i�o0�BMq%���t�\}f���pk>c�\�E��!����b6�y�I�U�=�#lƔ�i�8B|\a��44V�������R�;Z��F+�Yi��d|3E��k:�o
�ۗnDq�J�e��8�����x}w�q-��lK[+�iy���M�guJ.<{NS��EF�&�D���<wb���Q"2��N��-�@!���}h��u����Rr+��"�t�\C�Z��h@�,��r.u�l�B^��}�Q,㉵y�jf4v=s���S��@���O�����B��x모ӂx��HJ�P2�e��̾^�ŨL�	a֜�u��#��`��~w��У�S+Xf�eh���]�N��n�0���ơ��/5?�O�R�\wP,�B#�<�l��1���a�w:M�����geR�";�OԔ�kϥ�mTG/l������hx�v5�}�!i�/��{�}U]`1��w���Z�İ���ѫ&"ƣ��MZ�t�{��Q6�����!:T�=bU5��=�����B_fv;F�f:���*�$J���Wq>�pί�t�X�k������ik�X�S�
��I����W0�,d�u�}�v��I,g�φEUtBr��>4o��Ցڌ�S�L/��� �� Iشk�!\7ʉ� {q�~"u���������;�+S�U[5%r�H4o��c)�����!yO�jo�`Ey6
R\iyN�d�v�j�������5뷳`K��SKC-<��Ss�[�T��whW?�ߖ�`uجY �@�ﯞq�^���]/{�Ty��K�l���y�F�A�`e��Z�۹77�Q3r\L�Hv#��Jc�����'����Ax��J��]f=G#߁�~J6\8����|�}�w�I�0�b�i��x�t�~��ij5a@��`XV���>�����_?I�NL�0��b������ͩ��mG2����|�t����^be��}RV���5��AB�����)����֓"���LR�^�Z�4��&��uK/N伱VZԶNoq�rGlv�a%�K>U?Q�L������t�8`��z�Ƭ�����K?�6,��Ϥ�Cv!E^,����a��^K�&%l*+#y�l�rH�	����zq�S��B7��y���g�A�?��&�(�x�uM�?�:�@	��^
kNz�u�*@n.����s��ȧ��!0;�_��A
~&d�k[1n!ո������U���N<p���b�Ξ�n�kB��wJ�ٶ�l-<�a��g�$�݄��TÃ�;|A���b�x����kƋx�W~9�d�K��V��NXj�)׾�e{����ȵ��|���
 �W\�����z5��N^�[�$���h�k7Wvp-`�7w*,y0�R1�?�JN�\D�l^y��j@�A��_b��1l�H�>�V
f\>��
������e�qQ�Bk
jZ@CU��EtL�~ �u�<7�ef���o4\�����)���d�
�^�����_k�zi�g+>:gk4���]m���h�e{���l���o��b�/�#<^?���zYfvr	A�x��0�[���Ǽ՝�����X��Oz��ߨ�BG�R���X����DR#H�(FjŢ!����������)<�Ӻ����M�7]Mʐ,�K@����L�kr}�.�7��i���v67J��6�Af[��; 25�O�~%]�
=�UQ	�a>g	�ZG�¸���2�����c�7���>�Y�n�:B�͗��*��Fſ���Qm�'�v`t<|*0S���z���o�`&ˡI1��4�Rߘ׭�]�1(`
S�S�+��~�e�����'fKR�,ڧB��U�,��bO����=�I��UxlR��h��-����/��l}�o�������S���ԷFKYi�mp�^H�=�wW'��P�wKt�-aU��9z��:g)��-����l��'-jR�o���'-�l&ǜۧx뺙��@�S{/'�t���ܚ��XK��Y+%���&~n?G�0�涜���Fe2;,)�C/a�XWo6+�x���q���q�4�����B_F̴���EL���q�C�������Wd�/	��j���q��D
Y�ʽG�=�ؓ�����ǣ��z���_��Ulߎg?�i|�cF��`\IX؎lN�� ��8o�`[9l����x؏�Ļ7m�B����,h$�����H�Y��,��6�`uB����(p�����������0.Ҋ�D���#��e��̳��{~.OC\W�����ȯ��I�����1����G\�����~o��O)�h�K���{��4?����?�<����9�'�R�	EǤ �c���sj*3f#����U�����&����ݴ����m,9���^)�L�~8>F&�,m��1��^j�v����X?g2˪��h��<'fR��T�n=u�..L����2�I+�_�&UL��w%F�kѥ��#�JԺ�OML��E��!�DÖA�Bo� =�m��R��s�ba�rb��,G������ 0��gG���x��n/�� y������A�|m[s�����T
����߀�{�o��K��\|�M.�w��r� q^ ��Օ(X.��ʎ�i�0�w��a%E�w���g@��$W�#~�B*�tk]jކ�,�X�Ь���NQ='����I��DΙ�:�������,�G�m���C��X�qڳ|��ӣO��!�����p��(+*���O�&��bv+�a7/4ʭ��Tai�����B��tF��1�ɝ���(�;%2h�N����I��X�Q-'<[�e8�j����m�P��8� U������N�ba����.6��^?$�T���[�O�4g���# A�5A -���Ķ��^V�MA{��F~H@i7���"�&���2p���%��6z���lW������3AHHINY�$$��b��<�rh���0�rf��)�1:�ۤ����C�U�͗O>�`��6<�
L��"[��WJ�i�e��Eo���_��
�*A�Fy74�6��vlղ��.n�T���04D�N=^f"pL rⅰGF�n:�[H�����"2�π;kg3�;+��c9���=Q��B�?>3X��[�u��	���`�*˃{p(�یZK�����/���%��Xr��)�ά��;�N��͵'�˯��#/C���R�cS��]�C�5by۵մ��"���x��f��D���G08H*}��?�D����"*�Er"߼�����so��Ė>��y:�Bd�.@Q�n�@9 ��bD�>J� �R�ps$=^�v��9z  =j��V��sZώ\((��䖖���љ�@���m��˩?q��M��J�7;t�=|�1�0Tf�Q�� �؁e��� �.+��'�u�*)�n@p3?�>gQy����a~�B7#ñ?�CnH�ޑ�\\��R�T���Ky�HqT�.��J����*�v\�[�.;�Y�9!�aU �M�'O:,��$��eN_I���n������F�^���E,��޼,��Z�XWLZ�˞855�L܄?�a��W���ɖ!d �n�Zԟ-�Ԍr&k���#��RO�v$T���D��f�i�T�%�=b�����X#�W��W��Q|�eH�)�BL���X��g�����'f���Q����⤔I<�Y��;��p"\��-+��#�KD�vm������]1U|�	�>�Z#_m�,�[t�!B5�|�뮠�<�,H2��s��7#*~f��A#jᥪ{c|�^�8zأyY�խ1Τ�,߯��+��o_�T�2L�8�y���o���e�L���U1z�.��(��fn�g�7��TÁ8^�r�mb�9���-PT�_"K�:�&�6`N�����%��� ��DC�@�\��?�:*oۂߍv3{R����U�@�|Յ���X�z/�π��	���u��Iu���`�:Z+���ȷ��aR눒�\����]��'�G��ݑ¤�^;�׋��ϔ���~�rALJ�c}f��r�@�<��Q�Z^��a�R�Fi��?ִ���S�p����@E7_�Yq�/K�
�y�Cn���s~�C��IDU&��b����b��I袀� �;�³��#���1-�z�������S�w���Q��n	'Z�Ł�>Y�?�����"v�~q�a��׶��_���~��[��s��jC�A�8`�H�������^���n�>!�AK��X���C�V���;���H˹=�[���LݶMiUn�O��k63��$o*�c8��8e�`-�K�N��?�⿬���D�ϯB�#��cBYݸ=�����F�F�}�c/ѺΧ�[#l���t�4�����0���R��X!��{V׊r0'DVB!���^������t!��3&[׶�i	u������4Nrtw�7Rgչ�{���Ƌ�G�=�48��Qv���X{�j�bP��7�{寮�S_���ø	-�j�y���	5�����$l��/�knZj1��e�Џ/���2�_�=��5�df��d�����I~I�ml���- %����K������.�9�n�ܬ��=Y��/9^�����<�i�9�~{�n���)^;��>�k����{�X�>���|���ÆР�6J��m��PΞ��s���IAV�"���Jg��9�޹0�h�0�3���	�-��>����7�t�}5��<�8��XG1mj���<���Oߦg�4h�~�~G�z��@^(B���Z��X\�l��ɦ������������C�Ǻ#f}6}M�����TWm.���[~�t���]�!EA�S?����<qv��Dc��9��L�+&�O��َfO�{ɐ`@�œL�l������/Kd��u���gq�f1z@cY>���������)�b����7�����^��?����ı�]r���2"�
��F0PT�:aM���@Yk�M��У��q����J��+���������W��&6~ �n�+JKJ��5���O8��j����:�-�x���&�s�h���� ��uf�9��(�Uwy���4he���v҉��m�^�Ӣ2��*�R[#
�ozr�,x�$r>ˑ�v�tu�X�v�-�NDM��b�E��ȿo��Q�L�`v���	*��	�[���.��zd�M�=�
��X-1r [Iq�TsH��c`��,(�{?����D�m1	<a�]\�\��� cܞ�8>��푉�Ӵ���WlyO��zT7*4��f�	M�o�<��=�H�47�Id�pz����.��yG8�Q)�kvEX�Wa�9D�-?Y�y�Xy���o�}�X�����a�Xt���
�̜���uN�Ԟ.�-�WF6����n�~���6�?MG�����L+��iSԭy�(S{Is�z���՛�v�ڥ��۽�R��!>5��/��
��|��_����e��?,�{�y�|f��Y�C|��˟Pj����8�pC�w��&S�
C,Xj�f�Ő����\c�3�/��9�ӆ��nȞA��/��O�6�����uزS���
�G<we��65ڼVY�~�v*�}��0*v󔯴�V`������=6���8�g�;rt�	YWq�G�h�P}���!��!��3˯�~:�K�}�c)�-��֡����"�\_��厬Z��o��>S�\6�!?e���n�<o9��
c���y���*���IbU9�Pd�CMqLĚ���ÿI��()h6��^��;D�J'-��z���[�����[�u�~54�����԰���L�Ҩ��4���|;��8?�O��'��[�.�׷6&��ǞR�ּ<�l�%��I�&d�`p�q嚙��E���1`%�'߽jn������8WZ���hq��:#m�I�P�&}���z�2��^{�ő���
(r@x�%1O|%��a	W>��<y��V�l���EJ8#^�6w?�XYa%g�D+'�9��������\��#�,���w}��Ӱc&��?A6�k��䵠�wx�i!�Fb5X�M�#R^l9>\dC��a�(o����S���u���rbE�,W�m�-�Ѫ'��Ɋ_>��������́�|$�O����{��(����!}�Z�\��x�4`�c� �!Fn=�9ۯ��B�����B��W�|N)��~5}��5(�q�Y�3f��L�}�yVD��$[I,d������_+5��5���O0��(�7ld��=��)�'�����5����7�5{�����>+��g$qãcI
���[���m8����'���޸H��˩����H���4mє������9Q���h�!��E/�]w[�U�i�C��}e�.|�	�Ή�S8/�\���K��Dz�BOI�r���K s�B��vh8?}j�4��˯bw�M:�
"WK
^9���AҽsvQxG}�0�5�_�$��,�d_�x���l�����r��#�q�a��1������"�Vj��[t��ᢳ�SN	�3�j���m������-�um��Eb:���S�S�Fi��OZ!^MD轩#��_���е�b0��8
ꗅ��RkS���mU�H�`�Ql�&.XCWm��r�s1y��P�X�**䑓.Q�;��fZ��`�-���d�P��eM��<k��-X�e���9���������9s�E����%{��ا6�0�����L�������U�蚑.��ۓI}�]0�5��rϯ���ԇl>`����gBߵ��@�� ��׸y/Z7�]���OG�|���54^^����4�����y�q^�@q��uzZ�qΫ,
�W^{���s�L�r�<���������q��5ƃ'OŪͧE�k���r��}�"Ǭ1_a~��t��x7��#���:�ĵQOa �2�oД���1Y�Lˎy�ÍB������-;uv�iY��O�S�1W��Z��`��g��:�奣i	J	2��]:hn������4����d��#_u����ڔ��@ԫ����*����b� '��\��CS{�=#6i)�o�^�Coc�񌃣���d�䡸�����7_���lB��*7Ϛm+-����7ԕ�}��E�z3�͒�$,}�qo:�(�/)��#5��^ ���%_�&���u�(����,���R��MV�����?UTrE����N͋�@K���O+�r�SK�����$�������Ї����dtΗ����8/�e�Y��3�3s|͛G}�ǰ��Um��ļ�<���!��yy�����F,���j�V���e� ��@�1����Ь�aC���_Q���
(��+_J����@�mA��Y�<䂷4����;���N\�kkg�romA������'.RҴ4�����|'?���\ao|j%y~�������[ s�nC݄8�����*ڿ�$���o[�z�a����~������E#m�'�����)\�Pt��:�¦��v������r1�1T����ݬ����P`�X:��9�2S ԭ�݌Yz%�w���T�)�?�`����4��x���I[�Y�G70aT�"7.�] OH-F���Q�V�ʲd$N�җ�g]����yޏ��.QZ8DK(Ѐ{��{����;��"%�IԹ_o�m7 ���y����mT������>�
�	�0w�L�Fl��ɱ�+�AeU�o��ߛ����P���=���C?n����"��%��G�.� :��H�\	m�E�!7����t�^��y��n�)�d]t����ó�,�Uz9.�xgx����"�0e�G�b�_܊�Yk	x�����B���e��&�9D�FI�i�7jm�n0��K���&��T�}�!�:g��)g�`���c3����7����<W��t]w��i֮'**5Ŏ�Î�����T.�Mt�h,L�U̫REdX� d�{��:4]��f�#�����C�h����w�Nxڟe�`e8��2lT��Y�Ѧ��^5��O,�����l��7�c�IѨل�wlX\�m�Ғq�T_㿟��s
�w�Ϻ"�쵔-�.,=����7��S#CIW�?�՗Z�ಀ�@�9nŧ�4mL���Xo���(�)�u�|����lٺY�����+��VP��O-^��
Z�);�O�����N\DrH�����F�p�������fO
Rn�Z�F@�5mEkzŪV������@��,m�u�J���V]�퓍
��OLM3!]����&O��
��e�!ϛATg[V	B�s�3g�F��6�2RF5���8�����A�o��'�g!�0nA�"2���5,����i�u��n��:�a�&J�w���/�"����>�Y��*;Mt�z�3���n�4>�r=gʯ��j����x�H�o���h�z�}��x~�,p�o�#����.r�\&�b\(��[�	�	��\��hJ������V�M�ȃx�@��y� ���W��1BaD!��8@e�!7�~���_@[�]V�cnq:<W)Z݋�#�F�0�ɿ�O�t�8&��"�?�EEH��H�s�992>E��G蒽�Ze��Ȱ�lʇ�2�@�|���y>�^Ưj�{��N��?�=foc�♐	��c�9���22#�`�����a�C�va���Ѹ=���+���&'�;̇�ݑ��NMނI�d�����#�����.�dg8ŧ���R:�L���_g&��_�K~�b�%�8}_�j���`X*����lj�-ȺȔ��� 4q��8��k�?�d�^tf��T��E�ɍz�dх�>w���0������Y�m���P��!w���;�P��J"&��h���@�$�����6�D\
�KF���e��jS�"�T�-v����*k�S����c�\��C��R �����+���<t�?$r��?�}AA�E�^1�C�]�(�Y��ă�F�F����_w��Q��B��A8_�啂6❤����+�.�zV�S�Z�8k��ؿ�<�I?d�Y.0Ȉ�h2/����:V]R5�ף�{���8�O�'u7i��z�M�1nv�A�<�"J��I�؟�c���u�Jk~b�Iu�����s�w�,V-���VCMg�:�>���/( (�B!仢kB� ���R��J�Q��K-��!W*�א�a)�/:4��lb�9>5��=�0Z�R�̮0�jK��a�ux�|7�T�_��&C拸ķ���Y�=�PTR�W�,=�!m�y2�}VY�Q��/��P���o5����c��n�\�8^�dZTR!��4#����:0�7�^�q�C�\1J��,������0�(}�bWxC�d,H<��_�8��]�yꄵ��s������{��M��ݞ4{�N^��?n���q������(�r޾�a�������
�<���+��ФŸ���P�~oOȹt�7�G4?d��I�x����9�o�F���d��}���NNp5��5F���z��e����kz?4��}�ET 3%���v�b��~E�T|�f��*0c���1� ��@��r'��wIGEd�CA� ��"���+m0���Zj��I��R�!�"rZ�b�ߗ5B��漩)B��g�v� 7{FY��
W����2�q������ˑ/o���9?�w��-t2�B����ZC����>��h�n�X;�D����L�U��ߞ��'��{�f}r68��.v$ ���w��˸��A�N�E�*��+H�`�sJ����4��K>V�w�F���p�����`j���#��ƞ��F���g#\;��;����Mb.C��-+�	M��H�h
B�ݾ;��t������(u�ߒ�A�D�;��G��k�V��h�y)㾵�l�C�����<�pg=ʪa-b[�1m7i�"�K�#N	��٣�	OT�t����,���޾F��]�V�sDE��J�=G��vPQ^c[�Y,���h#��E�X,wL�7U�G,M;�ω뙱���]Hs�l���H��7Z�ڠIXgPX/<s@	�=�������%nS7̩dʳK�*���
�Tѧ]72������.���_k���3�i��^�l�֗�ˌ!�(�I���A�U?T:���@��芝�>�h�ź�t�m3���0������΅f�V���5�hw��OI��n��M�JJ���z�n�~ʲ�Қ��`h��G�Edߵ4�դ�K�5�-�V�n��md9j��wO7Ш]su�(q��`	��� ~Z#9?��5��i�;37im��B��1�g�����ݯ��~���Ƥ�cf��^QI{�x�uET��m��I(�P���$B��L�]��!4B�U7�a�F�G�)�J�P��Hr�]UO��0�|��7W�ƭ��ާ�bL�1Y��g#���be7��S�H���}��v'nm�w[�[u�+11?�i���{+�~E^�؊�ը�������>1��;�7͠�Vj��������j$0�{��r/-�I�����&��ڧ�(S�E��nl���9���c�ˆ��Ү��b1� !�K�C�'�|K�(�KhACJٴ^�	l0�=܇�뢱"���z��>۸
��^�d���huY6)��[�ƒ��AĀ��k�7�/\���oL���+v_�X��HrniIk��;�4UԷ#�2�:R�M�����ǺͣI���d�����>��~A~�x��2*'�`�MQxf�5V�n���}z�R2��2X轚����I�w�X�{�߮�zJ�{�~�a٨?s���K'�1~�e>\����1{c�u$8`�a�y'c��ۢƳv���V�0)���@*N�f]�$��!���<�z�^:-U]c?\q����'��t�-���'��Y��Ve_�T9�I�BdY�5"�(��	�y~ܿTb\�9�t�_-u|���K�[7������p�d���>G��M�Z�b
X�y3}a�j��?�m0�ze������h�S��m]��(�eX�R7A�|��Pg�Cpͼ�TpI�x���u�n�u��V��{�%ڌ�bD�|$����T���N[�~k?9��o� �ʿ��Gt�z�Y��/t��T*>��jU�},#d.�$	@�J�� ��?�ư01�)�o݀�e�E�#ndA�sGQ�(�����\�QT-���4^�H�F�|z$0q�ܽ��)eẩ���~a��B�<�_�L��|��і�
4pPF���+̃i����7�܇L,��d�b��*��ݽ���=)�����%�8q<"z{#�
�'}����pT��GZ���;3�e��΅�P��	<�i��q紊�S�~�%�]O�V׍/��x�}c&O*�;�_��7����*��13��I��T�T�`�x��.nͦի����@d�j?I���"��O':�ݚ�,1���ƛ��s�@ލjL���O�{��6^�=ًm��e�����c�(��6�n�Y�#	������x{��g�o)u|>�[y�fˏXw�8�j�+�*n�Z��9����bi��b�g�C���%�����ǀ �)�Q�<C4ܔ�˞�{[W��lo�Lc��J�9^���>��}2Z�J����&��O�����6��_x`Nz��x̸��W�^���i����HO�ҤҔL�u�}���H�_��b��h�O�JkԴ��y0��`f�ܟ��3rO}��G�� � �G�rUݲ�� ���5%1�fQ�~�-��pQ�C�HN�B���K�#SO�EIuS��@��M�0t�Q�&����$�U�|~�v���U��S���Ï��u��u�G�4����Q�&�O�Q��J)��8*�&�&-��� ����NW�7��8�#���Bp�%�F"İv۔K��:xx�;�x^�}E�?��.hR��t�y����7��<��:�*Ow�������#�g�1�jU���G	׊=}��zG�O>�(@!Ċ>������M�#����X���L�uV �����E?$�M�wU�,�%��,�)ruqD/,�A~���H	�o�vĊ�Kl�lЊ�b�Ӗ�h�����I8�����Mh2�u�1cWc��%�����A�Ҝ1U����R��Aj�Zf�*&��Ǟ?P$�@��>FƢ�&�����}~������E���,x>�(�W�Us��|X<caG�e�ٻ=�C�S�ĢK����v2��8y�yz�cy�"����	tAp��)$e�p;�B��|�!���(���p��}�,�L ق�K���W����M�hq"�_�gTX9]�������� ����/�棪� G
B �!�P�W���Y��B�mtRi���]������I��s��^��R�0�k�t5�`��44V�z�iV��8�?�����.���L�Y.��3n�m�Qޝ�v��٭�Q���z�,� �zU�� g��~vEI���i�����p���׷�!��)�ů�APk	��=��9w;1ǧ�P'x� ���	.��h�a�
�0��oM�ʍ��U�s=�����t��{كw����j�#�Z���k3������򷭿E�pV��N���	�M.FG��Q�8���/<�����{�V�3��_\'wj�cG��)Ƿ������[�y�Q�|�o_S�?�s$�#e՛����CŸ��:kWf����ó���9K�_?Q2��h�����:�vCݒ��`�?��[)���u�[ܶ�O)S[���š�1	ĴN&�_J>��-K������^��ҝ튛A[�����f��P\ȩ.���d��f�~�cd ��R�ޱ����>�i������(8�R������&�]"�f�A1.��t�04���c6
�vg�X�b{�#.#ϗϥ�Gs]��1�%f.rzX��k�OGv��)ι2 �;N'���C��!�O/N�RW��dt�ys&�Q�*(9�f8�Ex��mb��K:"���c�y%
���fV��D͸Q,P�5:g����`�u���nZ����_*���{)���+$���W�2A\71ǎ��!R1q����	�G�|�Mn�/[+RH?1�o�����N��^Ck�m���}��M$^�T\�+U��gY�*BQ���6�5�	MPĮcد���2����3=��I��g7�K��(�^C�X"R��}�]��?�}.�hŵ�6S>A��/���Ĕ�4>>�a.�W��AY(���ql�̖]����ؕ�E���j1��/� ��OU�3'P���HFw�~�v��� I���7q�01�-��Pפ�P�%%:��A0��z�U"��~0Ñ����fy����{������$♏�J[ܥ,f�"i}6}�	�_V�D749$펖��6aH;Z\yKeE��G���\�?u�8˰�+u�Ğ����p�COi��)ϧ��x���p�x�{��8<�8�<��&{l��;w�|�[jGˆ&s:#no!�G�^@�8��A�L6'�WB�1�K>���o�M7���ԫ�}��@,��{н�*�<��ئ6Y�l��59�\����Ky�`+�b��g opkw�6����Z�2ӛ0w^3(Gcj26<~7�(���DI�ۻ#P��N=r��G��_$BY=������R���#|Ӵ���s�.�IX��~[�#Dp�bby�F��G��9�`�{2���3�w�S�Z��7�K���e�-<�6W�qR��b��9K���K�V/�5�q`Y�*Nh+:c!5?B11_��V"b��0������#��䩎��ƴ�u6�+nּ�@��!7���^�pm��h�d�F4#J>���S^d[�o�E[�"�C�/�@ˬ�v�%9n.R�-�4�?�|&d�)*�K��o;0�
=�����?�_+ߟ�Ѿ���/��DK�ƻء@���m�>"k0'+�8Sʌ"�^lo@�K����'��Mb7TT�����?p]	�������Hत �ޟL	��] ¢D��9����v(|�CCd�^N��oM�ӛ�Ǵ���j�&g�/_�/V.���f �&ρ�hi���E"������C?����+��a}V��4��= M�b�J"����QI�pS�/RV��ɴ���+i��m�Ӆ��h���r��a��Z�t�Rl��/s6Wl �8�z%�QOBn�����k��;�=�$p��X�-Ϣ�%�]�L�Т`&� �׹�a��Lz��ؕg��!t�jP.�9e����2�è�_���|��L�jh�l��9>� *Xܼ���]c�"��+B52*$���֚�|Qv繒.~І�E~�����\-��^�T�
���x��)�* 9�����}>������2�2����,��{ک�Ӯ�����jh/��m:��/։�ٯ|��+[��1�9��BS�g{���Gv4���ӊ/��I��ɿ�졣��5<wp���+/�5(��5��?���yX�fN���s��yh&�)n�����}/�?�Sq�U�2������_�z{͓�!s�yM��3�ч��>���j����k-Q�?�ؚnGh9���tF��_*�|k+�-��^�.A��M�Y�۽���r��?��|B >Ѯ�B��Q�|�Dߍ�l��������P�\T0%�;C�uH�;����|tr�*�P��r&�l��f^�mb�A��a	0��}���PfR��I���}�e��`�Oj�u@���,����E�P2Ԅ,o��S��٪i>�]j�a2di��Ş\=��6]`��@��e�dw�𷺗��\�-دYYqZ䨳�ҟ_i�,r����LH~�YM0My�5ƶ�(&P�9�7������3�75��a���k|*;t���ՆH6�E��!�W?*�E�)�*�:��ժ�aKl �Ғ�]�M^sJwW�vn|���F��,B��q�ص�|�_�L$*f�f#}����V�n-�:2�O��s�(�������5r���(+�yĀع=Cd2���f�[��2�;S��5�-�0k�Rob��W�r�B���n��Q԰�&�fݴ���cO��9p��윒�ju�|?�s*����K�TJ�+��+��NrER`��0���+6j]�8w�In�s�����~LQD�tGg��խ5^׫5��ғ�މ癰7����qW�;Mg�W��[����6�����Ǔ�4�"$E_�{�ì��unH�&S1���f"�qO�����ݫN@`ڽ7��5�5��}�0��ס�k��E&��I�O�#S!��0䲦,g����B���*M���ۚE�v~E��
u�_�Ɯ�cv�~P=��`����qm,����3���m�N/j�h7<�|�%�# Ig����K۩���z먨�'lE@��YB��n��.��K�������n�ZBҥKX�;��Y��{�s��o8���=s�u��}ha���Ejy���v�|�c-i�S�Я�=u�����	7�klX������f`n�x+]꾖���;�t�q))�6�?V��{�:�Q�~�m�m@�FG�#��"Q�H�mn�b��"�>�R���.�)5�C�3=x˯�j�~+ڻف� p�3%�JO�:�v���:W��'9��!���#1��������n�,����'`.e��V�T�ڐ�����g�������`\�H�)]�y����"
F���M�{My� 
��Egj��[`7S�}Qv4wy���ղ�,�޻�
ԅ�+�s���J�%}��XS9��UQq��]�	U(�{t�s����8>�s�)�O�[U���b��ՠK:��#������g�l�� ��g�$��.'`��?ui�&�4)���O֚��Z�s���ǍFa?���K�P��M�|(���[�7O���΀�r���$Q�?�R(���#�Se�XZ�#���|��O�򷏇ت�kn]7��P{��kx�"������7+�@���2��6��K��:���S�3��Hk��Y�{@��X��z������V����̍^��I�,_�BT�����>eӘ���x�[�6�D��yy�N���[S��Ğ�~_N��󖿌���X�q{Ϻ�^1&��L�>�i����z
}M�����X���(=ݍ��b�w��X*�n�1iI���k��Zj����c�I���n���|$d�\?n����������n8����*	����ZR��|Q'�_X�@�b;��`�
�չ��f値��� :3��zH���9�A:��ށ��X����3��75+� V�<��<���{��ku�����蛦��B(<�/����Ȼ��m)�揰��;��'>5���dl��'��{�5�d�&�ە1x��E��#�_��2��S/}/[�N�m�}d]m����9U!��K�ec`W�bN�]�Y�V�
������C�]����wG=gE���ث��򂱹ٷ7�t��ri7�[m<��a��F_�X���_`�u��p�<�W��0�@��Z%u`~�$�eq��!"+���/!T����8O d��vT�\�.l�L������.2j�q!;��T ƵD:J��Uy����L)�Q�9G�cS'}����gG{�1j������Q+��c�y$(�'F�*��#�䦁oȆNmx[t��]Ɖ�l-�h�l���"g_q���)Y��B.�S��؉b��a���'��>��`�G������F^I�F:Ul��)�]0>�r�����j0?���j�+6��b�5�[C���Du��|rA;wXt=��)(�������g�P�Gx/2_�t`�񮨃v`��HwМ�����gB�zR�s�w�Cb~FYp'�lW*����8��<�pݰ�ZHa5�K}v�>*�.�}����Ɂ�s�o�V�rk�_g_1w������6Zo�ɺ��!#�B� )'-��������e�.��[^ĕ|�s�D���[�A�5:.�8���K�y2hޒk�t�˂�%�B]��_ċ���y(/~�I�n��i-�8c��i���^�ba�?���0vBhK퇈�����B�x�ny���/;eL��r�/)h
{���+l����4��O:`�1"DY4[X,K����J�����+��u�O��]9O���;å�R���]m͚���g��jl��_1�G`�&�.7��c��^$s�Kf��L��9��`?;=طn<��]��+/�L�F��3��ӃB5c��St3�)��	�/�E����������l�1IEc;G�W�.��Ś��kv/p(�_�ׁ�	t�dS�F܉2l���XY���՟S�J�'+�+f���=Y|Gu8ׂ�us�%�!�G6��]	#�W�iXuV"�׼ņ�K��:�N;9H�_x�
l�F+��CMFf< �lT�oze����˄YC$;��pa���Ƈ�|_�����4��f^��d �`NƷ3�Q*��(�KF\�����V��Y4�}Q��%o�m^�v����j�e��B�wyX�n��kc^������]2�@ZN8��qG>���l���l�-�0�?��C�[I�{�>�)	���Z+�-�����ӎ2a1�V���������eԽ��_�R���6��j[�?��� ����%|��v'�����8�~�8c���b�F��>J:[�^�(t4�X��m�#w�����-�M���<=��ji�	�����E)Lg����^�r����r�G*�
<~�]d�,,#O�^d�R�!υo��a�;��J\M���=�|��@`嫡[[���sd�s>_�*m+�ה/�;4���(*���rU�׷��́~~��k��}��@�&N��$����	HP�B�m3�W���6�{ɍN���TP�$��5[Am����#;-����tm���q����~wϯ�ɔ�����x�Â�m�J�w��
e�f=�_V�`�u'������cQ��OV���,pT2vK��H<���oI�),�%ys'���y�㕍� ��O]�$�m&�ƥS��x�?%�V�]A��갇��+�&�~��BC��e��]˜ʔ�Xח���+PDċ��6jsu�	�C�f6+Y�k �1�%��Ӎ�+
� h��Da�BH���k�I��ǖ&G���45[B���-n2z"Մ$���7��~��DBP���K���Y)ဪJRR�s�L#��C�.��;$Ôb��<k��`�c��]$1��*�1��b�ؘ�^���:i��S�㶘�dR$����ݟ�ڣi��j����{�Q��^�)��OjKP���o��z�V�~�M|5�}��C�G�]���:	�rƏ .I8����pﯸ����S�+�o,��ݿfi�˟�i�|ݫ��Vrw��<�����%n��k������M_:�xG����WdĦd#paR{����T*� !���y<t?����!�G�	e��6��r��Q(/$���Ʒ�F����R�f�3������~�op�p�
����;�9�sh+��}1�?^&YQzT��$��+�WifD�uu�˰��X�q���}]e,���:��}A���z�.�2Λ��af��=�M����F�]ͽ8��~��[��)��������_��Lsf�b�v%׏ �\���I���$�
���f%���_l�[�ߵE=|��9����*�����G!�ƏX�	��f����֌rpf�
�7Ʌ�B���OIK^���,����y��.����M	���#A���˩*Z>ߨ��^���[�H���'�7���H/\��~9_��U��3v(�ݐѰ��І�q &�V֝���\96�P�J�73a,U�󹕷���c�(͘����L�d�ߡ��W\Hy��gk��q�g�f]�XyJSg�iI�E^�)�^�j�	o���B����Y��H�XX��cv%����̙L� �a�z�Q����1�-��~�o��N���CP�8RE8��b+;���8�G��3���Ix
�WN�ű*v$>�;d�p�kʚJR+.D��7�0��}^B�}��פi��@���A�d��Tٜ��z�doVt�:�^��N�:����D����\=pJ�	���P�Ð2K���¼£��D>a�X ;�8���v���������47J���,-������Q�[	�s�#�M�uɶ"����l�%��,��b*��Iu����,�}�)4�n[�^�����H���RFJ�ӝ�)�\�ޯH��.��PK.���>:3EK"��&	Ǖp�K^M  �C)�p�^��%���?�>_ ���Z� �g�ܟ�pA��ʸ6_��&~�|��m�;ʡ��!�|Ry�&wpX��6�Q�N�2B����Ĕ�Zx@�Z~�ݺ�]o�����j�ˍ�Ͽ�t��ɷ�R��ˬ�QqM]���<U\EpT>�h���� rz�X��D�&�m�Z}��|1��H����Q=.2�6n���v*JZ�Y�s.M_ը����ExMfG�b����Q-d�:�����B���`�PĻ��m��%7�,^4`k�����N��tȹ������5
,����q��p?�&��[c��+=+X׮	ܳ�m�]iSy�S$�oox,7oE�N��������p�����렄qA͎{���Wy>?a��%#M��)�&N۬-�Ϣ� ��S�)�zua��z�;��:&�Y��U"�ьZ��w�}�vń�Ha�ܸ(����U���dCBr�G��������"��Ch��U��{m���<�е�$��7�&��r@	��qVH�N��f���/�KX�u�r�y|�<�{��2�L�(_��"8
Qu)���?g�q3e� ���ߴ<8�.��H��m��ʟ��ZySO����*���l7/EG�c�|0g1pUz��x$�)�$�/�@��Wi�_���2�?�k�3M:G]z$�*n����ai�+�MD.���><�!^�:~�H�W���3��MXm6�!>�g�[��P6��ߩq_j%�Q�P�jcJә,ۋ��u4�%Ǥ�	42�<��i�Y��u[��]᩶�KsG?��O@c%�h��1�ILr�W��}���x	��s\0�@x�&F@%j�"��z��R�2gc����;�U�BO~��z�ho�-X�$���s�ɭ�F�o`��Z���:p�+M�j-ͣ# �]�Pe�R���E�i4h�:��������3���n��k����;�_��䭹��ޒ���?+"!��(u���/P8vʖtj\���t�)I�3�;�$�v ���kz�LX���s�7~�uv��5iI����o:��x�M8b,�7H��J��Y�~E�H�CS)9_�(�R�8��E��1�g��_�h5Ȩ�����*��,+l��( �(�gG�g�	����9Qż��a�6�$�g�n�D�V���W�;�FB!A����������We=B���Ԯ���6݌*%]�)��]7����e�H���`�L$1(��p�a������S�le)�/�~������!��^r�����S9�}Z��G���pun��W��i�ђr��T{f�h�?]wP"��? #y�{�#��:���7�	?�Ń�%��,��Cb=MR�14�b:l{{�-�����k�y����� ��^2�#��Շ�J|����xev����-��I��E�WmU���P68�5�ȑe[Waϐ��v
���f�c8��� �o�{nnG���y����]��Òk�3�/�+�Lf|x�`�ʙ�-k���	�_���Vq�еAulI��I)<e��"{X��AHv�&���S窾G��&�څڙ�0����WN��#{k��9�K�8�.^�����>LwF���-"�P��>:��{H!��QΜ/�D�l��w�wA�w��p?��٧��*~g�qY���*b�9]��2����ħR�D������#nrIz�e���v����&��=5"�w}%F~��d����M����UW���M��'"�8�fV%源�DY��K���䟑�X��};��1�3�|<�M��k+2��S�Y�2ױ�J("Ȍ1\�Z��?�+�YIa���sE)�'-\��pa�� }8��R1�lpTm��=�)Ij����l{���X� ��������wa��2�X�Ѱ�.�)��}ޘ�C�"��=J�.�>���?���;�sq�q�uAp&�*�wv�=9�=Y�OC�wz����bY;�G:��Y{	-��5 �#�}���<����:P��p���8�x��.����K�46����Z�#�,VZs ��ul{���BW֏�/���9�{¦Ƀuz����۱�K
��At��@	���]�ǩ�.���ʳ4��w4T�$��q��Ư7��Bp��âV?*�փ�� ���&�Kz�e��ن��{��W�_��
3�}����İ�g0er�'�m�O]�/����� �/,�� �}N��{^x΍#fs��dX^�
�|M�������s�/���-|�����=V��i���Q#U����L� �͍\I����U&��~|g��Cs	?b|�=x�p��LQO�}�8������@�(A�qw�+�@�U�˷T��c5'�&r��,�ۍ��న�ۺ��N-g-�x�>6Lq�R@mW#����G�õ�wG��%$gB�ӓ�ݤd
E�W;g�����Y�J��WV8�Ց����Q����lBW�I׬��'Sl��w�� i4���EO�7/BEɰ�*)�[z��r�h�曙��cy�X��8n@Z���-qM�h2��B�����E�ᖼ�L�XwPK�VL�켇���_`�c���s�Eߦ�H�����Gd���<�:��A �i)VX��o�����.���c�%��g����K�1`�>�|�rx՟�9-�A%|g0-�����hRf�Y߁ְ����rh���s����ߙ���RԦ�<e�*jZ{�U�u{L��3�o_��<��h��1v���=�bm󥲭��Su�:^Oې��쀴I�bы�c�&py��ddm�J�CG���v�6	͇Z��W��4�j�l��&Lm����0)��?ղ��a��/��W��1#ďL�n_
�0��5(�S`_i1[72?�P��[I{9����h)�Q;� Qa��okU25�I��H�U1��}N�[�Ŋϱ�j��:���yZ���|K�2����"[i%N��B"q���)R���� �a�u�ka���]4�7��3ֆ������>�RSp`? �t�.R2��������#��I�X�0����m��|��!u{��ϒ��93´�s�dR���TR=)��t>���Jf_��=�����7{�|P|W�y��-��d��K��|�d��e������9�3���pE����K�R�vtv��q	��ϥ�jz��^қ��@��'Q��R�o���	G� !�N]`	 �+]f�ѯ��s�����;���wS���x��pl��)oN�|��@ҩ���8}���:$�H���w��Bw�������'ܽ��'��J.���
���A�5��DR��	-c��G/�+Խ�w˹�Y#��[Xn�3J����.H�h�S������=C��av���$�e�6K���.���ɶ��!�����n�Ʌ���.���uJ=���x���7�=<`B3)�X�LQ2RNZ4���þ5၃A��0&OE	r�����g=/�"��~��lcpٻ���^*t��/�=��/z�z��;w�G�Љ�� o�'ZmR��| �m����Qb�q'��C�+s"}]�X�m�Ϊ�;��>Y�	u�&y���o�>�]e�n�Bj?	����Ñ1���f�S�?$�8��ɇF����xi��C��1z�σ��{~ױ��Y[!*H������n��b���V�׊�Ĳ�tt��O��Xϙ��Yi�����0���!�`��[���}�tR&���}��n6Za�ye�	MK�;�$xC�X��G�M�Z�@��=��;/�P�<�EQ�z�K���^��񓶟�	?�Z���Z
C�:�|&�MQ/��C���1�o����G���7�V��A�~� 뺿�b�t��{���Fd.N�;*�8�+�m��(��{S~�(�k.����q�	px�:���e�d��]�@�C��>J���J$ؕ'}`c#�����F!���������Z�����\�h4��wp�/pLɄ���]����G�?|=�΁A���I�Ĵ��e0�*��[�}��c�x�(���lr�j�����i4������&�7� �/A�r�����nֿ��%�o�f�q �<���.�����pge�CgϢ���д�Ì #���!�C
��{ڥx8:��t��2�"#�"c �w#cnIe�t3F�#0���8:�Kw��*YE.��k��,:fp�6���G�ī��wM�[�\6U�ف�_B����]�!�����d��0e�"�,�C�Zg��l���!����N ��8;sɽP�����l��J�kg�n��3W��w���� ,����7w�߻��>�@���S�O�(ede�2�/hr��?�h$�P#`�!���At�w��W�^�������6��]2iq���L��ӽ�i�6s���񳖜�ktx(�\��.C]����S���e������A�]�a��Z���B_^�sS�"e��FQ�zl�ߛT���?a�����ǔ*���g���9Tkׂ���v9����6�۹�!o�� �2��W�����j��hKW�̐�د2�g �Z0�	����ss��[^Ξ��5^�\���>�H���s���e�/�S�3�5�sl��8l
�ާ�>P�t+yA����Ǿ�}��&:��9M*�O�S4oW��[e��`}��]�����P�?ծ&��G�~�{���`��=����޷�;��I�yQ�{����DbCZ�ͷ?̢y���L��_��:6G"2��� �_�;�u܇�,�b�����������yJ�=(�rAC��l��5�A]�W��ҙ+�M��K�Ki}��C�O.]���jZM�HO)R�PK����$�<L�7�1\�qw��_L7�K��@!���S��a�����␬�5��d��?:�ծT�|����p������	l�j��_u4?*�������_`��As�j,��Hy�>g�X%�^ƒ�Mſ���o���:?������ͦ}S�����G\$]?��ΝahYVіi]P��@HL�o�$��������'d�Y��s�@�3���6���s]�t�cn9o%cq;qa�Dş�+HV���9=��:�����"��g��9���P�}�M�öD.�^8zB�4v�C]�s��-V��(�"dq%6����Hi�i�x���[D��w
�7�qu�)�<�����Y[���������|�=����JɆU���:��8��Ī O�[���W��_^ﱜ�v2*s��Պ��z��i�W��]�0 ��+�>���-��?�b1����֮�p�̗1��.'�h{A����l+=虲׉k���Xӻ�^�SG��{;Na�Zpدx\N��(���4�y���cq�3
��������֗������ޡq�. \�&q��
05>��X�>r�������N��Ω�[13����v�#����@�5~�j����Zs��U�{�H7�E4����B'I=���c�� Gm�I;�ֵ�Ee+�A(�_@�����6����(�K�[&TR@����6���]J����ؚ~���9�	u����]����2W̐�	��Q�]������7U�y8�y3��F��-���o�6�Kމ����*6�m����\Q\�]_:�ӂ�|�\ �Z��)Q\���� �sZ�X�����;�}��ysW��2iPw�5Up6:��?G��3��\c���;_Ep�*ix��/���`��b;ʗi��#잩o�/4�6W����#��H�<n�&dB����&���*$>e��M�M�v�)#s�ۗǇ]~�V���k��7�$��~8�o�q�zc�f��a����3q���.!Xz敳�V^�L/�c��P�u=���(�]=[����M`��F��z�v�{�clX<Qz�R/��R�:��ɰfoR�%�;��5l~��x�Mg�R�A�k��_����J����з�3o0;r󿣄aTΕC���������K�g9�g�vG���&�jBگvx�����鯹L%�2�1��ո�»����-�L�>�ʐ�mó�iK���.��N��W@�6x�NX6�U6�4��Z:�p��_����������nn1 ��q{B��6���������*�\ډ5��|ƌ�1"��l��߱�K���F��آЅ��q�X�Qan&闑KWk����Vn���-�?>}?���6���;{g�ʩ��v�`�1�4R��0}a� F�L¸��s���m��R�C���3<7�g������2_>��A��,�e~�q����낭#�9�k��gy$S����w�{�x��������F����SM����.��ξG-�c����ykR��M*Ȯb��	;�ص�ԠprkeX�"�����}���e��<@�"&��?{�YH+W%�*V�����$�z�*�;�{�!'F��{Ig���<�\<y�-]�z_�ڞ��=��������E�/.M��L�-:)��К'
n���(`j����QZņe{�v��R�K����q7AY��pE��ѧ-�>Џ�-�������L���_��~�[�X�h�m��%�=؈E���#o���?��ל��չ��.��� u/�&��:�m0ScN��5|>�����m�����9���dk�A/�bH�t���:^��{@')�z��yJ�}�d��@}(�bWܭ�(�^�~3�̃���e�Ak�n��5Sk(W��wl�r!��E�y��u1�ڇ��ϵ<����+?}ӓ6%0�$�Խ1�,j)�<2L+��qqo��"ht�,�1	i߳���pɕ�q#%�pg��F�������]��'$z�Ių2���U����������D��b�b�T�Rs|z�\���>����d ������o����WJ�}Lm��}�� �gZ`�9�~�������(�FY�E]���;;>�����&��J��{�c.e?Q��s��������w�n٨F/��\B�8�8U���J@�7������7څ6��xx������̻�[��*�0שf�����5s���^�w5����`4}�f��O�� �k�O7������tZ\�qNŵƹ���*b��2����z���F*�'O6�D��	��B�k�b�y;�f��|��ć��__4���?%`��0���:���h��h�~oH��ޝ��o]��˥{7�{bO죨ȳ���������se��0D��2��?�>O�>3�
�:�������~?��.����<+X��>y�w��ڕ��'���v &��|_3��� ��L
�㝢��B��g?âW��8���@�oջ�S5��tJ���©���eu�*&��%�V�W��=>qN���;̱*;�/���O����g��"��z��,.~<��Ĭ~/VQ�����i �>L��K8j�~��r��`E��G�z�*�Ip_��4�:Yo��(c/�FHO�cJ��x�r���Q�1�&�k�5�C�:��� ~1�����+����Ã�p�"�������ml��ܶO"[�	�Tq��u�<��Z!4�(�G�kWXe�����1�PHP	1��aW¿�ߨju�J͘�4�(����8���x.�����]��s�w79�>��/�������n93 �C�6����g�M��gS�
�ٺ� �	4���.'� W�A�M�'������HNn_���͘���:Vw� ���.��c_����X J�z]�5��u�Y��_�;%��z�}�Ֆ�g�������z�s�C��B�*?΁f>�ޔ+�O�?�n96/F8FX�Q��<��!:��3t0E�a���ѿ���	F��E��/��%̀�k�YM�����Y%G��������l:�� O ��K�����H�����Ԡ'^�:�,�>h;G�8�cB�:S��p��n����y��m��j�%7 �jq���cK���Tr9*w���j�(��b߷����b��,^��r���2zM:���"7�س:��O��' �_��L�*͏����AQL(O?讓��~ڸY邢�T-����T�<;�#0�@��	�Y%,���nX10E�"���dG>��f��$��\�� �;�΁d�if�f��U~�d�Z�ʌ7q�H�.j�����T����T���t[���0���߂)�BU���b�v_{�oE�����,�U��n�i���7z�Jh��
ÉFG�u������јG��Lٯ� nVա¥�f�E�UT��M�6����y�O���Բ"�Hbd�U�����������MhO�D��{�Q򣪷�e~�q�����{���=�#�/�c�ٟ��T�����ۉ��e�u�_� �=�΅x�,y�ʷ��q.9= ����Y�nӸ�����:�9��|���idn��P4{2�9b@��I&������9�#diVIz:�!т��:��>�o��F�Gf�Ɋ�̯��M̨�d�:uA�%�L�s_���CE;��/F�o�%�|�zLC����O�sA�2��S�����w�/����9=C���eŹ�(�6��eP\�ֳ�c&��L��#9V������°'����p��|�i����QP��T�t�@��io:�9�ug}�n�r(��H�,�"��|�GZ}IK݌���zCQ��*ý�O� �y���ʧ��/��n�$p��X�z�)Xj����2�>�V|��/iRɄz,1�=��7s�-j��E$��	ؗ�����wۄ&����U���pe�=�)�)��m%�<9�+ R���V��.��_�Mp1��0�lGG�e�ԃ�Zs�ާ3�x��#��~��rT������q��rR��������r`L�'c������RoAq�8RA�a�(�!��!�=�|�HPo�+��3ѰWy*�!!�����8�Y�X�ϲ1�|H�y�9u,���@�-P$P,���R����]QsJM���^���1vL`8�g��B�A]��jı�|����v��d�AA_�\�z�,�<z����a`gs[�Z,|'9�*��EN�����Һ�>�Ft��h;��m}1/�u��0il�^��d�MQ�Ԓ�P_���uh�ԩ��C��;�8�������q��ȆI����,Dz�����s�����B����xe�{sHl�;,��E� �O�m�IF�-�/��]���oK�5-'@�>��\
�nR����͗H�����x�{�P���;o��d牊�8�����rz�{:�Xg�Y�w�IA�B�Rj���?��f���p	ɺ£)�����â���������L�E[@��a����Ih�3X�Lt��Έ�
�rP�0y��Fr��7�Xژ���k�Cj�9�X4��*��_�e��a�Їh+Ld���ZGɇ� ����E�c�o�tE�_���H��|M%�qU�G�-q�����-V»���KJN�/�7��Cz�/)��-}�Hj���n*�B't�L�)Cu�0��¬�ߣx�Y>h��u��]�޺�`�����/O��u��D�X5��������P�:���M~y��y�n^t��gi�&2�X|�.q[��*�}��Z�!!��㋁����~%��":Dp�wC�,�F�1����+r��|g�ʺ_�NHC'�ToO�1��+��ȼ�F�R|��6�K��t�ذW�(�6�8�|�ҝ؉ۚ�p)]LR~S�Ik�"�?2D�Z6S��p0�!y.G*=��u��gd�P-Y��(��G�+���U���36���D���U���
��.d�l�9Wm�^��탌N�������
ޅ�T�N�� ��k�Y�m�=з��,�N� İm�=���M��D!,����*u\�w��]A�H0�p ��V�/��rV������ꤼe@̈́�L������C1(Co��>�H���I��a�$��Rr&�u�I�%��If�[����������Д"���6�0��&�!��a��}�K��=���Bl�׋<�c�����R���8�ֱ���_A�-�{9��b�>�>�нcKq"&��#N��i���y+�ff��G��޵�Ճ1�|_s)L^�=�(2}#CR��u���!�RD ��۠��G�]����Z�Ny���;����5��Xy����:%^�ˢ���$_���Nm ï�3B��,��&Nٷ�;F�ʍ�� ��jƻ��7�ۈ$�
�QO�O�0�$�%�Ao�s$��&x�k���X�U�>&csK��lSI�7N�ρ����o�K����8�Ǣ��_?�l��_bS�>
+�L�#�Kt)5W�c!��}�H+S뭊Ī���3(�=$���%^=���vX��VWÐ|�-*v�@w{�Ik���%�(ƣ���̌Z�{N�����15��^ўi�R��t&��+��˹���.7gUE�w�S���' xʸ�l�W��e"	�h�w����Θ{rO�j��|�..�[|4L�ނ�vAX|�p�>�n����؟�c�p���R��Z|آ�G�*�N"�{g���g��$?	RB��c5���`� VQ?�j~�~\^��:������F�0b�R�S���wR$�5T�	dh6�hSr.��н��i�,���̜Nz7!���m0j�b��T@��c��Y����مwx5���[E�̍�_��&#�늘Ȯ�G���t��g��X۫H{ʵ��������c
lSJX��=ǩ��R[A	��l��S]�&��%��# Sk�o�[������n�wwO���h���wKӹ��_c����F�����~���DE��yn�[C����u�Sl��������:�H�ň���$>y����v{Sb�9�>�J����HNe�p�������|93�C��3�fʇ��f��'�9=,�6�y{"P/.9 �R�k�,Dq�T�E�ϊ.	�1�2:��8����-Z>��,��]�5�"-#cd�ͶR������}|�1����q�yn���]E�5�27��cI钙ty9R�L�[��.ԡ�/� M
�_ݺ�u~�e�⳺U)�>����Ms���+�8����u	��$�'k��uэAgF��u�����2�4Q<{^�N!er�=V�� �8��WM꺖u�8&;ڮ�X�iv�й��2��vu������+��ƃB�ڡ�]�߹��"�"wP�̟��e}7i��r�{�nz⚟R��9y���o�Lm1\̖��I���;;<�¦����'����?+���|o��L�#V�/E<V�i��6u��k~�o|6� 1\����rCEק�+��F��XD��RP[���Y)�w̕1���zf�w==��w�T�w��mԜ����U�P���{c�.U)X��>�"K�Q�/|Z��4Z��(�����`��mi�� �ͧ��bx+q�&S�[�������H5�I�J+W�[��*t��@��DCr>Na�a�k��*Yt�w���=@����ǿ?�C�:�N���U�尦 ��A�*h77-��э�V�E�q��k=X��n�a�A�{˕����w����e�d��.n�m���<��GXl�f�5l�$�*��$CY�����f/�[7V)�Ѵ1$������|I_�p'}+�tY�������/{��y �q^�v���!"�>��U�B>��)&[�P_>���%�)�0�]��
������RF��Bv�s婖���VD<�(�1Z	�J�䐤�:���P�\�g�w��z��U�j��[o�[ᗘ�x���b�e?�i��z�7����Z��d[��� /���-1���ơ2�x���bC�F����i7�e�����-�Z��ނ�N#ڣ�lWB���{���(^؋e��He�<4c���q�����#ڇ�o��J尺�.�H�I�Ҭs�l�]ފ2D#���?���h��v_ؖ��k�$��J��.^q^1P������ b����}�'J��*��#�I�B��T����xK��:VW��b�xzx����C�r:�.S,��P�^Rذ�\]9������C�	!-��p��п�~ꤳ�n�=�׃~X��@�rz���J�W�#i�/�������	*�	ʬ�}�2�#�G/�[ZO��rU֜b��_E�Z|R.����qn�|�_O�~���o�B�U$�ƹ/�-)�#����P�O:�p�{���Vv�D^�Dt��2��u�0��_�.��W'������Ur�V#�p�������WF��(	������l�.�w�I޵rѨ�j���݌_�����������.�?M�2a=B����-�o7W�s�qy�-���jƏ�[�O�h��.~&znq�5u�3�����]}�Q�lw��BLrQ?6����8�Xt���s�2������hr�Mkrci�Y$�6�!wC�^��W��%����r^��z_�J8Z���ip�y2����X�Δ"%O"��Uc��.I�=��TcS�!���7HEH�����kk׈����D�w���'ݣVV߹��y웃�!]��E�/8�'��[�>8p^Le�/�#Q��Z7�l�=�������i^n�`�噮Xy���������Z���р�����~����ڠs��������N�o[�{��-�+��$������Q���[l:li���ȉp�y����C�8���-�i4�s��[�Ly�@�z����F�cmz'�\��=�G�'��T��͗�ˢ�����b6oR��Ҿ8j�:`�˰P�\�&D֓��j
��-���U0Vi8D��* ����4���߅	�t��	�.��bk��K�vrQ�ˎ�!����*<qE�����]��P�j��vÞ��ږ��=W����Sɗ���x�]7=�mMMF��-�pU~���h��gOv�y��tA�s�O�K�VY�Ҵ"�Ӌ�^�B�Bۏ&_n�P�m����"A�0����	�pb�,y>�F�iiT�}a�R��x�uDnSw��,#4-�"DN�X-I�t�R���(q}Ԛ�>��?|�uT���S�(%HH�Hww7H�tI7CJwJw� 0H�ݍ�H��Ã_���{ߵ�g�����>���u�s�3������2!�~�־V��'��CCR�?Ы�p��[�N�TʄC�h)���� ����R��#�G+֩`�&ѽ�f��\(:v=T�f���n:a����wE͛B�=u{M����~o+�ډ��R�������Kg�n�v=�]�B#�6Dt9�Z
$�o���D0�(���<�wou[k����Y[V8�N�Z 
4h�[F�W��\{��|^y����`q*h�l8�G�Cr�g,JA<F;q��+���s\=�7�z���4%1���!+���g!/bRqy6���޾8�:������3.V��9��������>�io�^W�(�0<8nd3�:�%�
_�r7%��aoT��Q�å�"F�~#?���m镽x��Eh��<ܙ��*��*�������)�5�u���j���C�4�8��}%N�7���<���-��d��})^�=)�DNa�N?�9t�;�H���XVD��<"�F���R߼o#�}�R<>9�?e�H�h�e�eN�P�UPР�E��,탧;�ɊC$h�����gq��	����^.E��@Oʭ�Q&n��M�Q�8�Y�zlU�עoVJ�����H�|#	7�ϟ8e��\��u�a���;؈�Z��E7��M>>V&6�����>����$\pJ�Q�{�u��i| ��u�ћµ�|\�Ik@_L�{�D�3��.��'�%+�^ܹ��Ko�s�h��Sa-⻸�o�gȢt�(��'xVD�T}����={��%0z�����|�c���8���l*'���Poە�N��խ!6ť����U	���/� ��o�K{)�ț�������1���4�.V:A�d�c��7�������aZ�VH��D����G�APb�������'��x��M~���f���I�s��ʤ��ܼeh�>1(�|l�w�w�q��&��pOXRx�R֫�G�ko^ˆר�+�����v�����^��
@f�t�<3))SUȱ<Lh=�W�H�/���b�]+b9��`n��D}�G�F}$�g����(`���&qܹ0�xh�L|�����Kj�U��.[h!���Z�f��D�TdF�Z޻H�w���8�V�i�����5'҅���֗�o51�h���H�W�>V�x?�[,;�N*���|�xPJD2��������nG~�W	b��V���E�&�����&^5%Gy���W�g;���o����?��O�UY>��qTa��p����)�ə�<M'2�pQV�\*���B����G��h���)��
jއ$�AC���+t�lI[�M�n��E����,o"���&k�yJ��PF�lU�y|a�!�`ʱ��5~sMyۛ%�����������KWyef�e\ǒ��&��8�����5��������2B���փƏӇ|n]�9�G���/%5S��l��*Lբ0�Nհ\HL$Vޛ��IT~} �߾A������$� |�,����+S��W6��VP�<d�� � qҋ������������0)Λ8����#u9���l2/�a��~�|�
�P�PD7MI^YY6{��Da���$��t��
T���Rڈ�v{�'i�V5�1�c,����E#�a��w��al �ǌ��?}<��T.u��,�غ�W��4��پ?�ͯXó�g�X>��=u~�����dP|8ebn���FyO����9➚�������:oT��%$�Hl�j�l>� a��b�7t�����i�։=�A�nI�'��}���Y�_�|�?���&1wr���'�,�j�ҧ�5~���5u��F�,Z�pJ�z9�֪��@�s�$r����E&��2�ψ� ��������|���cߡ��HK��Ӳq��ba����
J��t�ЉSa��
�Qs��G�T��)D� �2��g�Rn�Π����+�Xeݒ�T�"Q�%�j���UV��G/kf����̪��zK��2jG<����A7nK(������&�<��a��?ؤ����5��j��ި{��� U�h;�}�&S4.>O���9�Y�����f���Yݽ�>��_Tq?�s��\�R����ˌi�zwbQE��#�����ץ���l<�.	^����ԕo�ni�-Q?�F��|����������>�W[�fL���+53�~�ߵU9T����:�SF��8�m��~�����Z����.<�̫��4���I�'��<������f�8L���ѫm�@��H
����9�o�Dj�;Ձ�g�V5!4I��R��&���2ˣ��t��Xz5����,'�ޱdL�oC�E�+s����v"*�/��/wW�+�ŏ�E�\�|W��Q���,R�ltN4F�n��]��!�s�~��B.���o���i�� ��02��Ј�V�@�Ӌ|�1ߚmң!��	3�j���ݟ��>�x]����v�\bHח�yx�LeR��q5����.�M'�v�:
}��R̸�	@P��f���"�C&�Qy�f@w|��Tdy�B��2�p<�K�T�~_��Q>��f�E<�������.��j��c�Jg\tTZ�xF�^����"����Pّ�wu��fq� AtU!��M�r	���H�'��F��Z��x��R�Y�ެ�;�k�YV��r�Ug� @��$>U��xK�����l�!�hl�?m�����2Xzn��d���jd�LM=���E�#H	_��#a���M;��8������>�Xm�9i�z��O�GTV@X@�'��{�t����L��Yi�m�I���$;��pY&)�5#<d�p����4>�C�-?�HKy��k.-����ðBo/�^�w�'X�?�Z��v
��eS�f �zw��*�7I�?��$��A<gB��["]��X�b�%����L ��{d���Z� �N���fA蜪y� v캩�Ի�$V���R���%B�sB�c���s�Xk��q�=ԇ�=��QФ{N:
K����]/*F�Q��p�VƷb������`<�l���	���q�q\Hxp��(ʒ����&�Pˣ��g����U�7�F�9PW��4]Y��3�T��AV�7�;Y~�G��\�S�{kX����-����n������; +����!����h�!l�ʖ�N�6\�v�@����ݭ�ܝ�y��&(Jv0��G�XMkcU�sN��+��K���2������5s��z�"W@�,�[p/�XHhٜ����?}SNF,��i)���}�J�C�N5ӫ�~	�j�pD�7�5t��Md�M7��cQ����+��TD3�e��T*������]Ftc�U}��xj��{\�8j�S�-�SHV=���Ip>Y��Gb|*��4�So<ͻ���h[�9�0��C�Q�0+�K:C)ojA�T���	�w�.���`�����j�I�����)g�֢1�J&�!�Gm�ïnd�(�D.�x	
�]�8T�G"�,#:�����RV^L��g_*}�z�H"�Σ���}�I0y��9��)V�	�6 ���y�R �J�e�
�=8\��)�QK[��t����\�xׂ]��wuэ���5��w��d�݀���',_�P!m���E'R�B�p' �SX�Qai{���9b�A?'���zP��|?9�OJ0\ܔ�w��$��݉�R?���j��K+�L�a3�=C�z<����m�o�O��D`��XU5��\��!�l"X�q���qAx��6Y�����@U��Z�2���OxP���/�ա�	�n����Ȃ����1�K��1��Y왏@T2����*~:r��~C-	�ܨd}ũ��[A�V4�|(	E�֤���b�n����맾z�W���E�3�Q��r"�c }��6�X5�JCVGY��_����Ah�F�-���4�|m��uF����&��B|~\������W�ɍ�������B�{��D�Bz*�WSh�I��a��g��<�/~��!a�6�%�-d3,��+.�v�D:aM	�Uൄ_�&��.�����miL�a>�����#<Ja���ޒWS��b�ݎ�LޗD�����d��)��qD��nۢ���O�3Xn�P]#+o�@���h��N��/ܤ�_���E^�-Cb�����mK��h(*2G�v��mӯ�PW���(x"1CJ������eh?��߸w�ZjZ�~�N�, �e��w�tF��/TV�M�I�O�SC�q?,��q�x��y��FՋ���3i8T��죡���$���E0�L�Zڙ�I�:�F�[��rrВ`]��r��EG����!,����U�l�+�G�M;�F�/��r� ���}�oq�
S5G��k����s:��2	���sq	�[�YfT<}�a���pp���K��p�^b�b��s�R߸7ns�%.e���I:�ϸT���dj����O�__N�
/>O�Le�E391�m���,3̰��}m�T��_��MK�N�����t���r)��j�H<B�%�,�I2��Bb�Eе��!��v�Q�bB�2�֐���׳� �����E�D����&`�)���D�t�*E���5�u�������A|Z���2\�O��}g3o�<��r7�1�RJ>����
j�������&�%Ei>���s�69��(wOr�\�B;[���z�V[��g
&�!#%���_�+!_ւ��LTV��3y�Zx�s�x�IT��̀{�	�O����5F]�_?4(ìh��v8�8v�S*�]�8F����K�R�{Q����{�y�A���;(��Z-��h��xK!�:>��ְ��g����&����b���[7��!=�q���h�n�x�G���T7/��
�S\�x��W)p�3꣊,��63\����?%�hV��������<�,^��}U�Z<�s6��|+W��|�����x�PS�4^��ߖ#v
A�lʆ��!9�1���W.,���}�&��F�,�h���͐��@2B#d1	Ro���M2���,�)����K�R�Me4Q�d��-�qw��!��V
��خ ��t�ǲO����G�p��AUQ�]��׍�`���C���+��3B��Pv;T25u]Y/���j�o�w}ե���8�ܨi�;�Nڤ�p5��w� �p�va��y�-a\������ ��O����W	^4���XPtrg&�#Ձ&p2���͘O|���Ea�ȱZ<:zTEt36	��dR���}� �����$I3LH�e�Q>M��g���XM���_m0���y$�P�A���D�ER���1�nM�����kn��!�%���c�P?�JP&X�������p��"��t=T2R��z���=����<[t��-�&��B=-(�9*GGeƵC�U���\��K��=-��;uYxZѶ��U�Un�su︿|A��-�����~ѧ�p��i�G0]oDÖ�43'�9�xZ^m�:j�N՞s��_>ۘ��������s���t\���	��i�~OѪ�kK)q�ǣ�9�fv2W��ա�U�l|.�*��J�rQ�x\sv?:߼O�W+l���o�]GP|��mܔz���Q�_F��a�ٙ}���~,�{�l��+*HE�}F�O[�!-~�����B�6������/�rc�ht[1 ��)��[P��~q8QI�s�5!O���Ҩ�9Փ�J�@��y��v�_8�mj�},x���p�i��v��*���iaYaV�Y��?^��o#�."���c+����+S�T|�$%�����Q�X=H�p��Zs&FϬ!��2ƍP�m�l�h6���囨�>�dlu����
�kq�SV�֊GS�%�qa���͇	(D�;��:���Az�]�SK7X����&nE�9x�U�ɋ\�d˾�?ϣ�iQ�襷X�W% iO�,��~��}<P�<|�~	h�H��Vy�C�zO��k�����o)�\4ԢWi�݁�J�d:���I�Aջ��wx��k���'$6=�ڣl�e��V|�!_^"ٖ�D�q��G\x�Kq�_�� ,�"2hU�2i��I���3�q{h���g������d��Ą�D@�?C�m��
��D8S��r�\c���5��� �x���,^� |������y���m|ћ_E��8v
>�'�V��6�>
�:�R��{��S[@�wG���[6)�ԋĥƨ�U�7�k�����24r�w�!7��B�P64�}w��c�#���t�5Ľƙ�p�>:l
�+I�����#�z�͟^`���@R[&��|����$+�o�k�E%��'��S�ԋ{)�jf�ti�.�R=g�l~�W�Ѣ�Z�1�#�H�1D�oC!b�z����r���ͺ��B]�풯>V�W�5<�BQ��2����Uz�������Z�BO�O���8���&�~�`錜�0��x�oT5[TL�b�����ԲUNqp�U���Z�\c���#3���c�-�O̱G��bt�#U��V׷�j�I:����+od��\$����ςuPD�jM8��i����*f���
�:���VK9� F�o�zM��:v='Bn��m�A��3#�W<�4��1d;�����h%?���扢E���-�xk�k2��:l���4�_�V����R�G�q�2�8�-],A�$���3���CB*����S>���Cr �o�E�E=D��û+����)�r��]�\+t ��W�E�@��@�{�Ʀ��JB�d��w)+�EƎ����=4���meR[��]�f%����C��]��-�=IJU�֎��4|�zT�����_/�9܅��2
�d,���}�Hj�.m�Yg<Gت��s\�D��#�~v���m9�E�i0��z�:ڃ��E�@�[�A)����+���
2�"r[N��%}F���m������m3>І¥�k�+�|�K���������kaa���[��6���h����ʆs�E�DI�A���ʺ'z��䥌ðd銕��g���#�Z��2����V��;���3dqh
[�|�����eȎ�U�#�0�sT�(l�g�a�*�@���+�}�Sa\�E���
ّ�4�Ȣ�������dQ�Y��?9e�-`�t�X�<Ӄ���U�����aV�F�A�'I��ޭ��G�Gܱ�(C80�ˡ��yV��]gÕ�������GF���ԈϻO��¾C�}2�䘼.6�ouM^�%/��Q�㥓�aT�uW]v`I�L�t<(�i�'�x�C�8��F������a�
*��aWQ�Ll�'K�H�0�;���"�S�2%[�,��Ȣ��P��W"T1�B��?5yJ$��'I��+���﵊ai�����������FwP�'�&�L`���T.d����d��¶J۶�rc-�*�S��3 ڨ�jʮ`�D)������ ���C_��߾౵]^V���~P����>�jN�)g:��
�暥�4�E�Q�]�o�q���V*�Ǐ?��&/��<E�U<�{W�8�d�*b^?����|�Q�En�S��r���Wv���)]Ř�Ψ�H��M�"5=Iڇ� �W��_�n7�o�S4.Rw��1n�um�����+	���?h%Ե|��:!��ؽs��0lDx���D���� �UXq?ʠ�Hr���Ҡ���㯳����	ӗ����m�#� ��7a�_�HS���i���s��KQ��\�s��=��&4�EJp��1�{u��>�c
~&��W�,�W55�c��ރ���|E3�zrഝ8%���jB��м�����j��bw)�8qGx��m��]I>`�XLD�圯�]L4*[�)�؛���ѭ�흿��E�M�A����Nя��tXF��3�	�K)�|�i���#	q;�G�)3�69?����OR*���I�+����Yz�WZkt��u���N\��־"3z$qٝ_x�b��-mn�@���	��׍Y?�Le�{�z�_W]f��Ib�<|̚��)���a�C�%~��6�VS���f��AS��a����g�޼PD��Y�*1xa^Ë1��KP�Ejf�oVG���%�����t�5�A�?=]E��o�@�-�oL$��50�N��=��Bߛ'U�pk|p�)`�Z�_�[e���6��m�c�^��8���?Ita���� \������S3v���t%U}��\q�7�������K64����?�p�m	��2;�4C�8�<i�W�D�AՃqv��@����C�=7��E��NJ�E��˴��,�@�L"������Z�~��\�f��վ.���Ғ!M�y�>@��҂��6V�E܈�x�9�8��W��L�l����W�}��E��ZG�����[���J�\90��`�Y��X�����1��ZE���}O����8輰�HO)��i-���"/�Ǔ$�X8���)���4����v���F���#��'U�l6}d��m�7e �%�£��_;����^�{�&�jN� �3߿�����>��8�V��2��?fQaz��ȣ�>�d"9�&�k��pQ���5�l�+8��C�q� �.jS���XX��5�˸T�,co�"&J�R"�;�,T�`XN�^$o5��
؈�Fj�IQr�*�.��|}SEg�)�l�;��K~�ٖd�_T^;��&%u�V�HV�܄�5ǋ��LI�=*vПb����� ��Ŗѷ���߷��0���T6�XCK�!�sTG;O��K�!�0���}�Đ'��W�KQN'�k�g�ܥ8V����e��U|�]F��vS<<�*��w�����}�]�����ߧ}���fMsB���8�E��X��^ԣ��-a�1��$���k�<�h9�ÿK�dG+*�-�|�I�
p��lQ*��?S�Z�%�e�R9�*��&��r�G���좇�}���Cu�a��H^����"K	H��
���pR!���$��U�
�]r�J���O�(���OT ��2��mj���뢵�>�Z)�|Y_t�m��n~��-%����J�p%�s��ęE"�2Lb�5b�S�� �Ais�#�
��y�0��)؋i:�z&Hؿxr(��%�����"]�mG�E��jS�ٍ(A��Ë!g��ϱ�l+Sk4���8
�g����H劑>�L�8
��������Rad<�D��h���7���e���ʏ���q�U���k���*�� �r�Nt�K�*� ����0�w���S�/�JS�!��yXO��u�O ��<Ui�1�+9>G���~Ƽ�E:ż��N*�4��}��FU�5FY����+?�+�^R"V��+��W�`��+[&�H��NN�]5[h~� uY��W�)�
��1G��/�O��+�2���#��k�L�)iZ�?�����w<
�ZK"�R�֑��?JH��$4U,�l/V��/Cy\O����&	��w<2=ۄ�UVjoۭ�����΂K��sq/����IcT����U��I�"t.���Z�څ��a@�U���gm�wIXڲ �����YxD=�s�s![�Ζ�dYw_�3�@y�M�U"k���Ťs��X�\3��5�~~�TN�b��)B�ZN
��}�[��r1��ei/�c?�q�΋��!��D��c*_f/���5��L�����U�km{���p?+��q_���^k"!���|Vo���O�����2}�{� ��K1��bw��i����d�:��P�4�x@�|Q�H�@�';h��i��rŒ���"H�FC�������M�S�*�>$��_��W_v
\&Kb�>Z���Pb���T�������3�V������L[���O�Z08~]������uT���S|~�4�\��}3�ٴ�ex?����6/�|D���.(r��D�Ĺv�Ƿ2;�_>y-�L�t������|tgH�5�u
,��4�J<��?M���Yf�e����xX!l�u�����i���_� ��m���Q���"�tj��"�.TB!��ަ�uFF�z~n�E����_�[��W�_��S(�-��,S�ϓ2{GS�g_��I�O�~�T��ğ��1����~�3Ry�! �¨�ُ.���Җg~���,� e*yD|`��󝬉~�����@��m[Ӣ���)7����f;�v�Ӛo�����1�(��H=�R���v�	�_{"�1y����ߦ���|�	\YZ�v�<`�(�,�#dDմdj^��S�j��!�[�CȮst!+#g�������8�C������w��Į��؄/���@��Y�9𰽖�s_O<�5n�\>�O�.E����S��
��D�+�+��Gs�=�	ą��z�@�d����Yv+�
"|U>�����_��1��n�+�.D���v�ʌ�9C�q������b�|Q�%�p��	��F�
�����ŋr?��|�n�l���D�b���ȧ7��i��$�0�=���ެ���$�:������s���Pz��A!�M`��%��).������L���p�� 0�$��!zQ��5���D[<��E8�N�bW-�Ҩ8���	ʼb�J������>�兣*�0����Ǔ������2籾�S��>����t������]b�~_��͘up�OY/��L�.X�	Hv�|�����VĢ_ӳ� P/�#̦����ɳ} ~���-=]�C%��*O����,���D[��Nb���円��O%��f���bd�H����d�?+A�dG_��ښ�`	�=����R�>�/^��`/�o%���OlU�W�3h�*Z�-`��dv��^ur�f��)w4n�t�Ǵ^���U�+mAt1��Ѕʀ���Ω�uS�9�������u��7"]��kC h�������_Zpχo�F�C0ר%?0�/�������*Չ��#I)��?LI�B��N�cӾ��a�$f�v�yn��ѵl6�n����7Z8o�[}[$_�����:�e��Ί���|�A�[)C�ȤԈG�@6�CF���_���AO�����Y��A��Vp�|f��@��^�tSΥ:¿�	��*q?�sH�che)�v&��4)��H�G��9Cl߱dB���$��y�Lj�D��3Ī&N�V�(������8}X^���mz�J�U��t7��Ĉ�8�8���{~d�YU��2xv���i�.~�\?st/���7 -)��Y�P�\�`�X��I8a�6������^'�٧	���-��l�W���S�K�o�6�~~<(F
�)�:f�VTc?�@�<���{	\,](�u�:|n�@n���O��i��p��C�A	���OVk��'5�;�>,��3V��D��������7�trtt��(>:�&	-%��+U��V!�
��?��x���
�zVE�0�~<Dx�/B�"���j��MeĲ�z�6L@C���k�;�"��e��;%���'h}�p�ϙ	[�/.8�M�&f �*Q��3�)�so���z�}nry�뛭�T=�|�B3Ik��"$���@P��Gja ��7�1�1FR�g�E5�,�~�Y<�RҮD���=��6�ټ6��9�LjD=:�H/�ǐT0��!�?.0�*��q$zSM"�4r[�H� K,&��
h�<�b#�.��_:���l#�E�\��d}B��r��I(}P���_�A�����#��zm��6�M;�q2�R���>�3܈,�_��ЅLq���u�U��)[�9I�4V��V3Z���Db�H�gޯ���5N|�F2�W��eیk	U�
^���]�W�s��CZmA����&%e���}�6U��|� ��"6`0$���3�O��'�q�����9��2��N���2`�k�����H!)��!F��8���c����������ѩ*�3Dn�,UƐ9Y:�JW�Qig[�q�q�,DN��B#{��,h�8J�m��o�&qE^�*���j �X+hՏ	O���� �~6K���	�}�W�m��zߋR�w-qk�Z��aS|�#\�3�%���n�`�\Ӟ⹁�>�Ml���S���o�|�!jZ�M*�)�C���d�E����V�ymc��t�4n�wW���"_w��Hj4/$Q����fL��\4\��o�g�}9�*�'}BΏ�[�Hࣲ���1-�@�����r\��`���i�ST�91��[:�ZJ%K7IK܃��F��}:v6	ϭ2�L5~��%j��T���Ƙ�T�����F���)��`��A��5��������S�E��^���o����/��#;�x�����hV/�w MS03��S�򨭧1ať�,r�c�bU����͂���;9B�p-����:�)����:Z�v�k��VS#�������ׂ,�e��������=i�s��8*�4+���?D��!���p��;R4�߮������/��{lW��T6i��Ym�ih����Rw�f��N����Ww�v�"�:����m�a*]�c����+̓TK屑SXS��+d�VD�e /�x��&F~�m/v��_p+5�%� M���Q��x��f˲y�ʁ���܎�����N�0��� ��!�J���P���v�V��3���R�A�&K�ђ�$v�=q�n
f/as��sd��}��M5�e��w`����ٻCLPLS�Jk�Q����GS�%m�	$�J\:�Z����V�+7�X���?}MS�P�/��A��7�k�ۦAEc'	��J7ľ ��@�۳ѧ`�Ȟ1�����I�����.�S̴D�W���=}rc}���;���N��h�j�c�t'�v�eE.X����}��d�?�j8�q���x̊����Ė	#���oO���]�Ȅ@{����TAd��⛽Tdy�!�O`A��p�7���V�TJ6��'(T@�/����?v&_���!�����55
�R.[�e
��%a�Q�0ԕ��B� i�yG��s5g5`7g��#$ݘ���GA,]QL��š��ߑ�","����e���2�PK����t���a��ߦ���oB�A���tri�S�j���4FpɟW�?����%��n�vh�Uo�A~}��Ƀ�daw��J��|1��x�f&e�!�G��<G�6AT� S7���0��h�U�"�iY����H]�:�%����m�#�h��F6]̖�&�wx��Wխ<�@�LXB�~�{������>�|n��ŝ��)��S��� �)W9⟂�+�.,t�2�M���`ɛ�Eϩu̳�r� �`��*K�i�Wa��a��Fi��g7��wT~˫s!������\�z�Qy��dv�I�6vW��LԶ���9�_8���ӄ���X�����c�l���%)���eL��\o��ێ�\L2���%�{�eŭ�H�|�>d�<����趑�IF�a���B��-h�I�+?���ye�H�0L�vk��y���X��rs!gd6m���x|TK�w�{��N*�]���$�57�^�^r͓�J��ׇ"���Z�v�u������g�c����D�%�B2�<��ް��x����Pa}<7�	Tu)���:�O։.����H���Nfڹ��_�CfiG�<���b��n���8;C�
��Ģ�ٖ�i�Ձ�(Il;e�IUv^e���P��\b�,~^@M�	�r#Ɔ.C}�l2�<��[y��ǳ�U��d���A�������P���D���n����@Uqh��$���0_���2��R9_�����،?h��;|ԣA.�:�l�����7��A;x�_D���'%?_��[�_���!���B(�wZU�w�o�7�SͶ_W�nQS�:��q��*�ɗQ
I���F�t��]�W���N)d��-������|XR��H%Q%1_cK���'[B���w�8י������w�1c�ND�~!���^9�7��T7
��h�况��k̚�GyE;���B7���n'�ݖ�[�Ο���m�2T&F���w��B ?)?`0R��r/Y�ك�[	���#{�J)Ga'�<wb\I4�Wm���?���� @�����rU!��-��c�n<ܴ5y�-�gH}��ZFo��uZ;߄]�������WC�͸�mj�7p���;�΃�Yr�G���ܧK�����E��'���a��]�pj�����g�´{��F�����-��/M���Ym�/�rP���c{�%/Q^��TGJJ��g��x�	X�|�6��_��M?����f�i������SO�%2�t6�a�:V��h�f�I�Sg���d{/蚭ґ=�X��I,���xM���IR3�S�=azˋ˥#��x�)2$s\Wv���6	=/��<�����:V����٠�݉;��"���[��z��sw0N��VsƘ�#���-b�[ըIk1���j��v�u���~�6:��  Q�H��c��qS�,IZ���:�v��Y�d ���k�@���T޴�)J�x`>�N�����:�ն�J/O�y4s��5��u��u�{�%=�GZ~o�ZR<fB���3�;���X�>�T}F�j�q6����#�J��f�Y�ȷl���z��v����D��Bs��8��O�Ui�n𠺆��s�h�1w������H�7��n�q䐳"��B
P7�xu �����En=(ǘ�oX��.e��>�%E�'l}	=xҐ����:��%����k�Q��/M�sLg*HK��O$��:j��'KG��Ž{,:}��.��Q_.7nO)a�)���)-��Z����EU�,;���2$��1:It>)����X(h���1W'N]����E�&}������������Qo��܀���.����e��來�iE�39��PW�4�yc�L����Q�mu�{(2�U������T�n��5/R�{o�Ps��H�ʂ�}Ѵ-�:w+U+��Ҿ8H�m�2�4!+�����k>RW\�L]�ş�JV��'�/
J88���QG&��G�]p�N���(�nz��S
���-�E�?�{K<����/Oa���F��p͒Z	?�KF�SG���c��D�K����d]�v�a��t,6�z~'����BH���� �mᒟs�"�����؉�')x5��?��P�`5�a�Ai�R�V�f��~5\�?��a��7�m�t���r�0eC͊����;�<�ʻzϑ����D��Rb6��r�7�~UXo�.��ZA�h��!����{��6�h�6��٭�'�Hp��v�w�eVA�<��;YW�iS��u��@0����H�'zԳ�jER�~Vo	l����G6ìH��
����RG��c�w�,�ꚣ��1�]i������ئ�jS𲎩iD�{�wj���+5���z@���S�D]��l��Ȧ����`����3��FM*����60�z��qq�A�$�����?b�okg[<	c	T7��E��-X��{��� v��-��Z��Z��}qNj-|����tY�`�~Vخ���- y�n���_��󙰎Ǌ-(��{�W����̜O�߼�<A��h���G��6^|Ȩ�Uk5a�m�@Y�L^o`�==&��E�9��2m�� ��%�+dܟbR�{�Vy���-K'=�~���*ޖt����4vH�o!u���xH����n�U���r����zL�V뷜��*�����,R���EF�����=w���sj�[��7A�_�Ph��v�� ��S��|6<[����;DՖth5A��W�$8[?�	I��?�\z����憿����g�q��ҢtE�ߛ��5$y�s��o�^7[u5X%�n�ɸ{����!�������޷6؝鍸�L�8�D�Š�mɀN
��zΦ��6��g:\��(U1�;�˳<\S����$Z��X\ѱc��N�{����x�g�!¨|ZCX�V���VG%��}F��a���C�� ^����GGdm�x6�;D����_�MxJޅ`�O���pi�̎=�U��%�_'iA_�,�C��u�	�}�T����eܑ���T�m�vֶꈵ�{L~�\�oQu�8�o�B��#��W�~��08ƻXMV��h���� �kQ�'ڰ����86�w�$�"�*���%�Ua��G�ht�]�:-�*�e�Ĩ(roB���g�U9�W���f�8=�
b\���%���%P�U?�����f�=�P�?�������!52s�i�/!�e�^��Ȣ��$	 f��(��΀��`7��K�"r���-.���P~��ݣ�|�S�*s�������*'����+��;:;�n���Vd[u!2�	B���S���9�����u��\��*L��4P>�2��[iE���BS�Ƥ ŝ��RS�*�A Q�`J͖N�5t?����ޥM����yv��G��bI��y��X�'��Ga�]w�CO��^�'��d��u'��������c��WlX�N���s�B<�x��;�0u�;�Gv�0�����;�A_1ĕ㖉]�qp��b:�0%�I�Zi�`H�k%?r:��i�s���8�n �K:8"h"xą�K%
�^U����c�2�Vj�a�� ����z߂�}���2��h�
)ܡ��C�K!P��V܋ww+�w+��Z(����{����#ge�%s���9;r�my�ޠ`Ӟ��Z5|ί��='x�� ���^1�5l��$�)�"} ��G,-����n�{��o.ӯBp:�E2������Q�\�ȃ�g[�]{���Ύ�GQl�7#K�Ͼ�N�G��~V�����!�h���%����^��KaE+ly	 �����)M:�WI�c����7�����saNS�%�36�'���iە�!����v�A�h�@��Sg�ΣڻU�-h|�E���(M�~�Ѩ�2v
��~ߟ�%��L|�t,u1�������t�6�Ӯ��UəD��#��]���� 7 "��ސO���
�v�bώ#Lg7�����.6�%]M7�>���"��K�%	�1:_�u�&�`s��1=某��!� G��v��$~�9  �n�v���g��|�1_�j���DdX^�e9p���|	��x#;}���V�������Y|��:�]Mè{��yQϰ{u�~��C�w꘸���	���jA�?�����)����|7z�J�,Zɟ6 ~����Ĉ�]�Ò��:�����ę<D\�d�ޙo^�wqR�.�NU�t�é�?��쩽h_�̔�ݞ>=�Ixk?G��($���)q�D*D��:�7Y'N���|������?��~Qx-4`��4\�1Уj�O��w>iEy�Z[�P��2� 0(���2t����=�r)�h����f,n�nY���,�	[2v�IVba��I��q���F�\q�zΎO��ҫ[�a񔕍�������q��-y�j��S��3���-��g������.}�++̧TX�@�h�2��H�Z2wŕ��J{2c�����x�n���ĳ�P�@ǦGa�2h(��g`V̆�bgk��U�>={}kg]�N�.M�ӻ*�p-�GVAjfq"�\�hN�2�"X��8�y{9v7�������T���m�׿I��O"�5�G�4�Fbq�	��m_r�G��vҪ�;��ş�ò�T��4y��ՒU A�h�U�$`�@��р�FKX9Ah��<&͍��òA^����p%Q�޺K�����ĉTo���O��H��"Z��w@�=x6���h=���Rv�ܞ|/�O�������P�8�A��!�R����uтB�}��[�W�ѓ��+�2��L�0��J���ɲ5������g��.*,�F�l��K����L��a%����:��o�˧ٖx�FWe=O�S��{CD��B�|̟끳/Y��|�I�.�U����(P,sG�)8�a���VaN-���/u̺OQ����n��,2�]q��E�pҊ:x&ۼ�1ߺ1�)��Si��(�c�x��^+�m@0(��9�\z���\{��0ϊ3��h��eɦ&�]p�;'��WN��6���Q�C�XR��'��TdE�-�ނN�N�����g�~���5s��� ��{�v���; s{��~�)�~����S��Yo�>�v�٢�tnD�(�(��&a9j���P�t�b)5�f���#F������l�/֕�Vj5'H:�k�<I�w��X�&m�=��7��jͮ��M��K0�d`�,��c���sZiP}I��Z!q� �ޟ��Jb��v7���_+6����磃���*kq��t�O�"�C22���IJ�8�Bkȵ�Y�S��$�
����0��BA�]Z Q�f��<"�L�U`x��h\F�:\
��X������^�h���xE�{�2Ͷ�e��a�u�N�����(�PY׼� M��:�qQ�˔��m�������?;gi&�)�m�)7�&֚1�5�﹅P��/W�KPwC�ڔx�c���Smė�.?���'����7�"Pv������[�y���rm���0����y�H��O/#��W�kh��g(dfv���f�V��� �F-�s�}���U�v k���毕�8�zK�MĖs�t�f����n�9��dXvyŦ�BD�����I�aف����)p�{�UIЯ��&�?�2�x�.����$T*a���qK��s����-��C�c1�����	,�E���!,�J*\��
PC	B��Λ�S�<���S��ӫ��^ٰޑG՝uW*��r�f���kR�o�o`�2��l?MG{�P%-��^5���\��;���z~���˲A�|�P1����i���㒁n/��Y�����ܶ�斚�yAԥ�n4�{�N�'�a���2<T��")�7�Q(�dȾ��N
���Jxԭ�n@��n����;G�tR$��v�=��+���;��jq|0��ƞ����{25Pڌ�T��-q�\�i�sn�L��0���j�i ��{��k��h���{�Ǯ�Q\�� �N�WAm�Q�3�ԛEhH��ܖ��7�U<"�Uߑ0�V��c�#.��#:j+��̆�!��"Z��t���8�j{���G$ 5�Y�jrz����}�<����E�U�űsXU5jX�,�oe��o�����f��%�'OC��f���"���<���*�K�M=D�u��,G�Uy8�2�f6�x���h��v,�l��E����L7�J�{B�S��u�f?�I��$C�8%}���+J���cR6mؕ�'S�J�����Qv����h�-H��,]C�A��qD�Æ�O�g��z�;0�<���>v��Ā���Ѹy(::Rz�Ĳ�x��\�9��>W�!�l�
˸-��6K@^�����Y��*o�Oe�A�2]r�^~;��|?�����-�	w^q����{�D4mԃ�D@�2J�q��V�2��*���\�5�w|/sVw�xZRHa���췺E�y<F�h���6�ƢkI� Z;��k��y�.��8�~��Z�����k�9\�^9�F�0E��C��gv����~bYQ���{7`����8���us�,?LG��:	��Y�e̖ʒӛ�B{G�W�Y��H�Fw%���9�K�Fmp��Lh������V�Y@9i/*�r)�F������X���ҝ�_7_�T�U{�(RM�U��,v@�j�P�E�}%B q	"w2�J�_%#3�q�dau�Ț��WF���6���E�&�d� /_DH��l�S��w��j����kO;���Z
˸�N+*v,'�㍠�Mgq��Qw��m,Py�ǰ,���@�ɜ˪��2rD8Ù�M������Ύ��v7Ҙ-� �
!�m�{K�*�0q�I��ƵX��e�6z�Kt�$V�vP���%�b��N��*Oh>D�tIuP�KU���̊:��7�2.�m�ܵ0bH#��;>�U�>$o�Qm̧9 ~+o�֋U)�8��른�F/����RM5X�o߆*}q����<��d�x�'񻢜g'
/T��7�͓{8@�[���s:�F������;�{�a��k����A��V�9ZC1��~20���قN�|�&�)����:(٦��j�3�Y�"�+y���Q{G2\w��q2��K���h��.v-'��/K� U��L�6��ۿ$X^����r�A6E�r��ls$��s��?_r,Y�YԬ#:p��!ʫ8���)	����i������^�`Z�ϫ��:SR�	�czIЛI!�K��,�3|W�]Hg�f��d���
�����!Bռ������8�0�x8��(Ͳ֜�����=��hH�k���w��Ҽ��l�p���M��Ä�D�#�R�Æ�Y!�a�ҩ��N�	�����٫<S�QLqW�t�a�s���L �4٠���I�3:�s
���l	5Q�+� �ط7ip�۩>oZ����B�Yy���x��K`��*4z�R)5!�Ζ "fP���&a3�XްX-U^��vqFW�/
�6l�q}#���x6I�/����J�����*�%-�%o��(�)z�/}l��7t��{ͽD!�ml���M�g,s_޴�I��_�A���p��F�_�v%Ի�!i÷�D�\���(��� �ci`�e?Oi��P	��� �2��u�'MeYm�L��Ҳwvz5��>-���Z�c��X�۲Y�Sp�c�O>��n�}>�UN���7ͬ�N��J�3��Y'�')����u��$	�n��h'ݯ?��4=
�K�$��O��/D���Su���ֹ>�a
��:�T��������Z����l4ԖAM񧯛�/zC�u�:��̹Þi�d]�w ��*D1����.�ӅN@���CY��ju��b��m�Qр�,�)ʢ1Q�D�����SƼ���ɃJ;���r2�[��Y��-�w%��x�#p��<���}b�X��R�����Fo�������S��Pk�-f%o[%�R����"�ܧ럗Vz��h���/l�����r��?�J>��7�h�Æ�ۯ�b*�	6���T�����(��~�����L�����	�#��B��]s*.�������( y��'�
�g�b�L��,"5��룀6�p�2�x�!�����ލI������M[et��A'�ؽ��ջ뵱�y��6|���� �$8�el��<�#���+%�m���d�}�l���?;�{�R�cx�'�%�#$J���u����wi�kHEV��Q	eܗ����;"o�g�Ȗi�ʼ�5��������~71��z�ݿ�u*מ,v����%R�m���\�[h�l�(�SA^��)��4�5��$i(<b�;$,��p�߇����V��/3��
7K�B���k	H�؄��J�Q�T@(��Ќ%MQ�[G,�*l�_4{?�:���oH�OId�%B$����Er8k��M���f�|5�=,y2�Z����ax�D9�i��f?���%6��T���Z.����b�1vhg�)�P$�aڡ���_�P�m�j;�R��Դ��+���l�7�7���[�$�Y]��"�?�`Ń*�����T�^B�@W��B�]��Ӏ~ܜn[�ȼ6���l�%�n���9	v�g�mt5�f�-J$o�qĘ\�y�;	�p��_�����+�`/߄���%e3s��lk��I��{5u:_�<�����)��Xő�̘����1F�R�݇������8<2�06rs��&W]����6�f٣�?c��B�}�Nf�K*�񋋣6K�p�s�cS�B:\�Ҫz��?f�|����S�����BV���-Mx��d �򮍔�Vvk�@�5�v�1���foA�2���.&��¼���A����������p�Ly����t0�;T�x%L�����Ƅͣ�7����e���4B�Xϴ�S��5�� JX2�J�r��P����H��w��T;��G�T�4��J߾���f���Id>��~���bur�t�&͑Th�]��@��u�e	Q�pq�N�f�6m��v���Ps�N�A�I
Zd�L���C�)�.1���ҝ������D˸�K��>/D�1ܡ���T�s!��w�$�LdD�z�{�9&��?����a��j��/���ʴ�k��������w����*�j�*�(�K*��9����}�«!�r��9"LwWo�$�;T�u����_K�mA���������J�! ����{����y�	͚�A���4s�{�Ae��0�3�i|�|��U��A�w*��άW� �>a��F����q��t.�\u9l𝒦3�>�'\�7������	�5��,#�w�L"!g �ݔ8�/��#��r]>=u��� ����#��d��U^�H���xTT�����T�IFZ�_���LԽ����O��l6U�oQov�I+}4�%WS36�@�����H��W���F��"�-�X"5�*�F��X�����`��q=6.7�  �D�~ LX���$�#��qv���d�O��	���?����F���g?�8��X�z�BB�|e<�U����I8�t��*R���w������۶Xʲ���ނS�	P���@2�����O�U�Q\B����{+== ��^˯_2�q�s���\��9��q�+>�C�������6�A�L��й�R�N;���e�%r�+�TЍ���gik�}������k]~������������!���
���h@�(� �ٽ�w唚}��{���,�X���jJH�J���$$�6vL��w�}G,h~��U`�g�i�}A�l8�O��7K�=����Ԣ�y`��S��)��8q�W�ǎ�5L�ʦp��6�|"Ӥ8�⼩Z;�H�k��C=G;{8�b_Dmd�*S�)Q��mZ�Ϭש�;Az>d[�9����7l۹p�.��vo��@���T���Sdr�hlB�_TM{X8��x�X1��/^�X��ok�36�?�0�RD<O��v�h�������)�Ѿ�[�M�`�+�WM!P}��ZW��*�9^���q��j*:Ⓐ퀶 ��ǵz�:~�"�#���J_��]��i��ڏ������b��U��B��q6��ԫt�d��i��DHCZY��������5%�CJ�1X'�;����.I�U��>�zGi��}5�s�X��� �G¬f��W�̗��p�=���Q�Uͺ��}~;��$_����kg�j�q��@��*B�-u�*-&�8��X���۪����ך�wu?�}ߗ����4�1#ju�O^�Y�^���6�O�#H�3��8_?��>��F4�L��� ���ss�ф����1�$�w���ߤ4Ѓr20��&Cg|đ"�`�29�g$��Q�Ƙ��f������T�nzj0rO�i#�sg$�A��!�h�`Q�@]�����i��>��X������/�F�~�SNaE2�����}�Òa@>�)�Ȣ��@����D���6��|?�-�ȃ8{��lߊ����������H�-�'�A�[�ц����9V��Z����:�GdXܳ�Ԣ�:���saaa��.JC����t/�]��o|�����7�w�*�&��g�v�:f<���Y�7��g:�h)pI�ZF�����|����<3�;��"�'�M�����!>U��I6�� �)�W��⃐^�W(�$i�0�T�����d�v��58zf��E��͛�˙4
	��,M�Yk+�.<4���g%���!�[7V�7�Г�_��l�-�� xD�Ho���kq�T��y��ع�;� �Ku���n��rI.p�}�)�v��8Bx����(��T��<��E�o16�|Mޡ'��(;��r��)�|�@e�7,X�*���!�Cg��Քo�.��L�u6�l��9+�����a�0t��i�J�HH� U� �}a�;A�^��9�V��H�U�%l�j�zBgH%����:f��E�N$�;�6lw����c��ȧ*f���X�d�z�;�C5�`m$��3,]ԟ3�Ql�y�'�O�hg����'���G���{{�T�g=9puXv"��3"��67����Y���=�w�oU%T{�߳_�'�yP�o��	_%R�~ryx,jO9���{�pG���e�{���G�dq�"�'��SQ��.��P��)�57��e�]u��+?�/&��v8wt���A��Ԙ��h
+W��j��7}���`�,�7�:#-�1��b 7ٔђ�6�H}��/cj�{���I�#Ӣ�\י���������0<c���<9gQ䶵�$�f��/��x�EoWAsf�t�<�z=�e?k�p�z��r� 2|�1�G��q�b{o?�����z�I���!R^��c�!F�F��Șׄn^�#�R���!C����{��XC��ʟ�,fh�/���ۏ'�5ܗkV&U�Cd�Z�)j}>�h=pÒ���eu�4���)���Sf��q-�ϫ��z^?K�����E=h�ݯK�ﺜ�L��.IA�aC.�B)ט%�.ٲ�"f��q��/��V����<�7w�l7�a��f����Hֹ
~�X���G&�fy�/;�	��n[�17\I��h�v������BD�E����h�ҭ-O5g)��G6�z���~T��u<O�V\���\�$NX�bK�,t�ݵDw���J��'��lv)vc�D��M!��]<+ӨK1.,�i�m5�Z Ŀ�^Hu�����,�^�4n��x�������.���)���¾�F0�>�Rc��1���OP�����2��Qh��'qL"�W?Q���4���-��<)���t-���%���9S�p�l�R�(��n��Yd_j��X2�s��Vt�+�Y��y�A|��*x�x��_��?�ע��_�y��d3�iq;��T���E(�9�q�ϝ�:s�ɤ����91��}���K��pY$�v���z�a!��r&��k0����oL�|)��ͣ3��k9�2��}n�e2�lCa�g1�}�qj� ��J�*O�Q��٩�B�ヿ��M����qaP�����g�r]���M��-�5E��Ua�U�/�oh�L��3!Ѧ�B}�#Z�ݮ�W�R+=�َ����Le0g�9;	�R��͢)}'d��Y�d� BCۤ�2���-w 
�k�)8�ᦠ�M�f��[�nX�p��2H��;g��L��k�Q ���:m� ��
�B�� ���+�{�����=h�!��e���(}�	댌�6
o��9���W��Ǣ
��*���9=\y���ib��-�X(IG�25�6��E��I�9ˠ��ۆ�^�qk	��E\=��k���LB�yM�IA���Q=�.�,�w�Kf��f>�>�|�F���j�����>�7�E���鵵���<Y�^,4y��Z��4�4�8Q�*�<����/%��\���.�Z^�U<*֗1<c`�����D2�#'� N�}N �dT�	�ٖ�t�$bB��+��	j�/����w�Q�o�ZN�L����b��y������Ri�Ѥ��
~��sHZĭķC�`��:�$:��}�H�]x�:�Q[�53�I �fnT�5iǹU���ͯZ�m_-����P�c�?��@;��|�q+]��9f�(���:kD6m��b g�O��dї��E��+,��5�ʨ��4nK��G�;�X(�+��?�\*\���������ȯ��ͭcB���[x���'ҵ���9]����:	��#�r�旽ՙ��R>E��챰l�;�3�*q�^��{�a�>D�L�u��ٗ���a�)�6\�54G4�N�G������N/�k�~K"Ub[]���6tV���L�Q�����A0��	
;ZK���$�&����ㆰ_��Te��U���ӔoF���:�/�b!�4t�z֋��l��_�-��l��rg!g������eאo��ߘ=�'Jm���Y����%m���/�s!f��Cz���Vݘ�;��n��5�:?3�~��҂��)�:�mY��K��C~^̫��y�}{�˰g��D�و���/9��b=΂���
Js7����/�A��"l'月��mYq;���T\n�A��T�J`�ʋ�N&s�g(�(f�=j�P�'g�����+���v�U��}"�����'A
~�?�P�-j�w�?��(�ף��Zn!6�ɬ�@�3`h���,oA��u-�-CW<�3a1����?j��i=��Ы��[SM6�����gsS#��8��)I-;���?�e#uDw�=��u��{�Ps�����x��}#�'ک�$z|>�);�|��n�.�z=\��b\HG���T���͚۷'�$J�%q*t|��G�5}g���-�15ܝA�w���է+6/ �M�`\�:�f�=��g��u]}/�����,��b�9��]Q|.��J�Z��#��ƺ��8�.�R�%���_iGON�֜H%���'���塢UyմQ�K?��Y ��Q��ti��B[~ڈ߿m��ΐvv�k��G�7Ȁ՚�p�D��%�  �V����Ws�Ldp��D5ٓ�]��xV�p/�(}�+~&�j�
ɾ!{NE��	�ʭ��Tv��'�4�����-�Y�~q�hy���n#��e�9���lSnky0�~t�5}���!~%�^��#���9���jg��bĄ�Bux����w�J(D���}o�vSF(7���u��+㼠��O��f�bSc��[��َXha��;q�q�������t�-pe**�':��"|D��;���~���Ƨ�OX��� Vn�-� qZtHpP�i�F�^�+p��͵yb���bSt�NYY�~Su��R�� i�|t��>;@@ld?�Ӕ��S�[G�@j��3��n��S�^���Q��T�^ K}�[~a�֮ ����\�cB��R�(yc�"0��3�8)�Y$���9��j䰹�����^05k����|��z��C��(���χT���w����e�N�^�*�-���.�U2�I�BF�M.j�4	%$���f���X��|��ل&K�t�\���7bϽw�Ws�wekY�DZ��0���o6���]� �A�W�Zr!5��z֦�ޔ�����u`��_g� 8�7� �'5��?{!���,X�'i��G�>/�В"����ء�b�H�̴�	K�ߵigE��ڑّiQ���,:8W�z6>W��
�����qB�"%�vD2=1�Fɉ��ȁM��(�|�>~��?�)ckR�s�_�?�VT+r�V{x�֭��ڻezP�r���ȩ_�>ac����9^z�em���0Q���Io����&v"�#����@>�p����a����Z��cC�����?rGS��#�Y�J%8���!6ÝO����:h+�΄�oLƤ[5ߙ2uR��F�XpQ�����Ky�k�u���sW8�F/���F�R�;��'JFy&b��-^Eue���G\ڿ7.�?�qg=. �4Jl�`�Fmg�ɾn 8�fE��oeg<�x�%�|�]ntsj����F�.��"bw�.���ytS�3����$����c�h|���/C�bK��9����왴ǔ�b�;��lJ���$�D=f����څ��3�k��y�x�
�m�)�d,v���3����Uʅ�C�扚��s��!��|�H��k��l]��<k�"�q��L
�t�8���"HIH�k��bf�x����>���"4����tkDr���t��v�����Z�S����!fm�|0��V0���
q���L�S<9�Rtq�¦���.����?�k!#��xj�pdG�~�Y��3��Ǐ�L���F6c�9Vqo�v��eQ�|��U�f��ZC�:�N>���yo�9:8��#�i��1��F)[<�Gx��{�(���{<ݸ"����t9M�2f����3陈&*�I"ˋA�6����%*�5�$9-wn��+�"/9^.S�y#+j!mE7�:\��3ݷ���*=*{F}A	_۰�N���G�Z�����=�ɒj�ft���,�Ot]v��ǈLK�5hv^�����ܗx��D���Q�3[�;��2.Q���A�m��.^����A�����x7H��e�p���X���jv�<�d*�J�!
�} z,�f��hQ��.n� | E3�n~�5DȰ��D�.*6��J��L��Z4D>�=�V��Ֆ?z��G��FA�0�*�+_��T0�!$|�V����Jan�<�/G���yS���ۂ���2��wE�N�;�Q�=ϯ�?o6ݑ���L��W7�b=ͪ>�_��b"
�Zp>h%��QǞ����e��h�,{�d��Tg��ha����m���x�5e&�J��M�ou�~�4XF���:9��
���-H����*���W7��r�;O��(#��j
�[��!�4�p<@^V����%��~���JD��)�#�����?N�e7�e�������i� GkQ'a�[緕�<3͒�����tf�* !Gl�`�Tr7� �^*�T��J:�|͍\rbT3s�砣�[&|�?�z-u����߮�w7�꓊��s�1N���*>4m����/_�z�gy����nt!+x�{D]���65�Z�-|�ߋ��~o ß��ѬD`}`�EVqg���斯�Nu%w������KV�󃅅%d�0?=����4E��E�t�Nu��Y���YQ��T�~�{�n�Gy'j�vZ�%ES��; ���l����ھzP3⩴J���7d��NV?2������V��N���{��~��Y����Fa��Q�
�j�eR�]�tA����+��0�-���*��~A�ŨX:�Z�����JU`���ܷ��>$Y0J�m�$Z@:~|�t��V�ʖ�@U!^�_��R^&��a^0�P���Y����N�"��pcH���@�ݺZDb�����'��龘��Γ�>�����}~ ������ ϙ��rM�k����L�'= 0X%yy�l@���١�kv��E�U1C�"���*AXD�G飱�_u�8�ǧ-�T%��$�P*=��Ӣ^at$s|���x��K�_�g�B?���H�:�����>q��H?V����?-x��2�'��crr��ᗎ�(���VO��fup��ĥ���vv6�����X���-많���"�M�|�:��<�@�$�p匆F�F��#*2������f={�=����?q�>����@��%���ңk'T��@�c!�g�\_c� �|>e)���k�?-�^��_z�qD��n>����S�X�9���޲BƯ3������k�����dɞ}��ZvU�v�J5)LPկ���c1��s���;Z��릧} ����В1aɰ[r�AX�������k<y����pLp�N�N�Ê�r�r�E}��rp�Sʩ�rr}k�����v����T'��盇\AUP�`Η*gXD��(��9������1�Q��mP���87A��9	��A�=r�֯&���b/��"�lYh�9�a1�H	��	�ұMd�J~n��eH�O�F�Z$�-�=j��C c�M��`��ך�[���&��{��^'�{��RLh�F��n� �ą/�u��q�סZ`)���M8U颩�m�����z�p_���=��7��֜���g�zL�_7r#�-�P�xRV�����k��;"(��c]��f���\0�8R�)�/�5��>���h��#�֞&�:������zG�5e�۹���O�cGS�yf���Ff�{����!N��e�#c��L�+4���8���2孡��P�_/� ���e�NY��a^߰��v|���YC',���,��0̉���-8!P'1T`r�u=��Q���w�|v��+��1H��*J0o�H��\j�yc��0v�J)j��|z�""�W}"Hߴ�h��ę��?J�N�}SH�|��,_�*�*7�J�A�pE�^���1�w��U5��H�y'�* %$]�x���?Wb��l4WI��h�/�¾2��◿�i�ֵx���sVc�ݛ��x�G�o�{�ND4:�?JM�#�RC��*U��1W�) 79kS�c�?L�	+u�
�b�OX�H�C�$���S��r1{!+�~��"�B���(�=���L����P����CC��w�u���\���5���yͨ~��~.��h���M�Ս�9�3l�َ�*���/i��{�l��ԣ�O5�A_���Ϛvo~c�p��f^�.U��ݦA��3�y�̣�6�E1�b�x��d��m�>��:u�2l����@����qI{�t�\�Wp��}��^nj�6��F��N4ey���G�<�ނ;n�V�:R�ᮘ�xb�ヿ ��(M^�� �M�i�Y2����;��}r��&��sj�)�]��TM��fY'͂U)�t�4�ß=$�����h>������AswҠn�|x�T=v�G�$U��҄h�@9�?�z�7�����ㄺjֆ7�j,%�Q�Wq���u�����n>���ޭ��;"�A��Y���Y�b�_W��j�%�v���A���n�	C�v9���y�ƈ;��Jwy�2�J�b����5�����v�x똿�R泝��������������/�M�|�$�ʥ:I�)1
���?�O&[X��O��!/��w��[�CfE�e˧n:��@��El��">��{-K/��~�lx�_��́{٨�0
f/���?}��_1|4�k�w!�B�O��*C�i5Ag�	T�:���c�M�z���o��R��qݻ�w��=к�4��GV�����������p@�6�l�af���jm��ԡ�ٽ�:���G8�������A�KN 1)�^Ļ{;�eT4b��zZ�k/������y�����q��W�!m���y�O�56�����sw�/'���^s$��ő������5�s���K�7�C)�,T/�H{��mL+_��7Z���Y��J������-y?��V��E~���2����<�!��}�J�i�.L��w���nNU�:�~�\�h�1�9�r��%ǰ�X].`�p��*�$��7��E>��j�"��ɿ˝I"7�Z�,6�^��v��av"E�����d.� ���ըÄj~�)eg@�]�~�eY!)�_������+�M�c�N���s�Rb8���tt���S�1R��ӟ����j�y*��6��G 8��~���K$�s.���o�F�'��^b����ܞig�e�v��]���&I�����]N���B?��4a���Q��œ^��:d�^��:��+أ��9�����V�[���w���"�u�)�n�0k,~tP�؟�l�ĦaB'��� �x ���+ �����KDB�/.]�'J�>��z���K'~�?��+Z���m���}�h4����Rl>����M�i�?�=9�w?-6W�b'���LBǹ����￳�tԧ�-3�������H��7��v�+5Nͣ��vR5C��\��L�,#�~	��ˑ��Mv:���͇��U��z7�;�B��}ϩ���y��JϪe�����������,���gq÷ӌK��`�T���v9��쁗
���"����w,G���<�_�2D�OY�|b�8�x�{���%���"\4��|]���b�ӑXX���]���>b��D��|��eA��{� �,_�2���#�}�t�~lP�3<µ�d���������b�߂*���C~��2��vy[���x��|I�ONt!\@�yk�)�'����ow>�	����t�e�����[>Mrfw��e��P�=�L�s���z�?��t�⫃G��N`����ʿ�'��:LB��O����ۨ�8]�O���C�����/g�؁���߮�t$2��Q�:z���^(6Ʌ~>a��3��K`7T*xӰ���`��ZWkK�m]:�u�?�E��<��~����U�Ĳ^��vt�?u#��S*��ۼq��4M�~��4�����Q�+���ᔯf㠿ѬH,�|�������ۯ4��.�v�:��W�:"�noB�6F\�����͔ٿdR\m/�r1K2ՠ��7:8�o��!�w"�9��b�u7��hj�{�~��&�s̋]�d]��WF�&�59I��m?6�o�3�aJ�m�� ���R��_Q���C\�ų����g���� �WS���T��7����2J�[xHߧW���������Z
����Y���{^�,=�w��Wp�Rӷ|,6j11����i|��7	�}f����s�y�5�ٰ�EU�V��q��������>)Q�?��ᗂ,��+�������q�7￀�_>���eR�����vEz&�����z��$qq,;n]sT"�v�ލ�C�o�9���_,���6���nW�6~�c�sdu��˿Hx�@�!`��2�~��nB`��7RT4�j9!�����.��W�{+DP���<q��A�_��Ds�ʀ�[��`�8��M����i�"i9.��������g��k.?0���w3�T�/<��D���5;�� �Otop���?E{��ʸQ�n�m��5y�Q��D�I��6�!�3�=���M�jfY�&��\3�q�.��(��z`�������nV�Y3�p�^�C�8���ռ��H�	����|W��C z�y��!��3�yi﬌H ��������%H� �Zͩ�P�/D-3�Έ�c#=��+�J�.1*|��XK[�~��u�ʢ��>if�����|�����H�����?���dV��Q��\��HK����p�Vr%vjT�ى_��N���ѐ  �Z���x�>"H|��BHԖU"�|�D�d�*A�Y�6���0
�8�+n�<�QjGk�~�N��t�X�u�u�/��S�tFz1V�(�jb�.�+�z�h�s"�^d�ߵ�Dq��Bՙ�k%5�C̈́y�=���"�8���F���{�:�/�4���kb$˔> ��o�����6�o)��R���:���t��~�W�K��W����1�jnބ~�f�}�����J aZ%E�~͚�}?���T�	Ig�D�W�{��5v��>	�NkrJp����_#){���G�[��`4ܐ����r&1|Α��J����&�%�M���T`/�����/�u��Ɉ`0S'�w�sr0��ٙ���u����9c�v���>U<�#�n��x@�j��\5���x#%]�g}!��E�~����H(��c�-���ްQ:���	�N)		�A@��F�EzP���Eb`�{����������</�pֻ�Y߸׺��Z�=�����O�V�A�;Ǥ��n-���d�XP�g5������L �ً�?ʥ�H�j����!��1��n�$���V�DM���I�b[����V�s��WO���];�*�S+`և3XI�+��ZBV.�xa	&%w�?��51Rf�6�h1_��ei�`N��e��ʸlGo�r��|�:�2S�h0��,1���	��=�����n�|�?�&�c��HD��,�$y/j�D޵[X����	 .+�s��#-�����*�g���4- mg.�y$�3��L	Y�e�wBpIf�H�&3�4SU��:��o�#I,��ݫH�<�h�첷1��ٻ=�3�mK��� �ɻ<����S�>Ӓ7�#�C��T0�ʍ�������i`���n[#���t�؞��T�?�5G�������<�'M��E��^�Jr}[f��DFn4��:���D3��#��j��
ݷv�t��tܢ� Ѱ������Bk&���o�����2�,2f钀�֟�w�j���-��x��ME���Ѝ�$ƿ�T͚o	�u7\*)s��R�/����ۏ]=�u������0B杛����\X_���7��p>�	?�*+v�;�5���<��}u(�ס
`G�F�������C���:��5���z[�v������k�ȬO�0��2�����-���q3��[�:�*�ƴrVB�[;���O�3�)�h3W陯��3)�7��B�d����j��������?�V<T�G�ؙ�[��)������E���Y��Kb���L��~����"�r�p�<%p�"�Cr���F�݃�XjO�B��`^��7�JP��Ɓ&�L�}˧���As�\`EiK�Cռ�y�Y�8z^�cxAtUz0��_�{�"�·Z��n��0V� yD,UM�V��](J���*!�xԇ�4��Q����+���$R+���zQ�/��g���]r>�I�V��+�u�ˣU�sH�/
S"x��}��>�B̢8�Q=ݛ�]�	�1��ё�Ⱦp���uVGͩQ�Dx���Y�I����Jh��H�u�#�%�����$��R	r�a{��aٗ��)M������6K�K����G9K+��3�iU�ڦy����D�\��`,�F�;��&�J4K�;N@Z9��$J_�i)6	�a4�4������o����	�-af"گ$�=Bl#3
;���0�Ew����)O5�-S!J�:���@�&��*0I�����i�o��tP<@�
�Y\�7��9b^�V4s����<k�U�d����ƾ��dw� �
J���k���γ��R��zL��^楮6K �N�W�،C���}<��#���~�C���T9�r1�L)�Mm��� i%$6c����?�I��`�y���#jT��P�W ,Cԥ���Z�:K�n����Z�KnF��_�7O���f��CrTq0 ����,k������&��h)�Yf����&�bg����Hr�cj��W��xnI��˄t��z�*���������cK�W�_4^X/��>���/�բAN.Vy�yIs�3�2�c?$�@z�/_��5��׷7Y�<��{�,e����jӹk��<�Ӽ[K�	||E�_�� K�(�U�:�F0}ޣю��W� `lJ�����r����5�3���.�d��ݎ�;����)�gʃ|�1*?��Ew����8����/X�l��X���%m�at��h����7����2{4�O��Z�7�Y�aN��v`�4!�nNT�7PF����"�7c※�V9ۖg��C00g� �)n.�� (~W?k�]J}���^�q�����K`��J�\hݍ�DT*�J�=�Wܔ�Y��~��e��؄��[ 1�N7�Z���ϕ��o�9TR������>�*[�
�w e6O�s)�#���4�?�x���ZW�	
�c_$֦���`���nPڇXt�p��>|�A����gj��/��Uj�L��`�уҥ���${8Ʉ��$�����X���ƕ���K��1+���S%�Τ�ͣ\3���c�	X�c����Ϧ�Ƙc6K�!��F���~��0���T��w���_�{� 9��}K9��:2����\���Cb���ep6	�p�W,�:�������+�kF�8`�ar�%LD��0�3��a�d.�2M�0�{�6�)�@����)�ٛ~Wg 'yj�:�Ӝ��qz�_�&&�Ob�?��Y�����MUAl����u����9#}�Fv�t4=:-%�jKŗN\&4+Z�f� ���~�,6�O�>5w쥳�b!d� ��Z?���R����&�Yr���Ǩ?�w�z#7�{ę ��3�8T�w�u(���}F{���%f�D�D����5PD���!�Sr�ĝx�G��k�wB���l��z��̶6�q��x�ob2�JA]����N�/pW�!�_m�1���55�l�_74R��"&\n�*�.s�t�v��æHg��Ig�j�����2�������¡T"�����'�0�N6�?6�=�[�:�c�UEF�i�ޏJ���w�G޹��,��z	�`+�&�f��q  R~��`�.:�(�f��ִ���1LHk'e�i@1���󌦂��n�?%������X��L����>D�)�]���l�>|SKUJ�b�pm�Zzu��2g��"`|�;̳R��ՏP���d�ou)����"�sV�w��eBr�ڧ�9n��Dwqf�����C�:���T����3�_��W�_�5��Q}cU�E�:/~-�ف-Ҁ4`ҫ.i�����[o��h��?Ϣ����(��]*o���J//C����S�$�Q�1 ���(�^ܨGznv֛e�������A���:l �a�Z5<&�D/��		f����&�67�2��pk̤�-w
dE�Ok��e��]�kU_5gC�1>�
�}E�����M���>��^������U	bLf�Y�O�srX9�*�[�wp��vZ���X����[������[�W�������{�&�"r���}3�����	��A��H�	���z5a�'eL:��\����TFSvv���0ػ��	*�D �aB�Į��I.,:��4�(E������k�,������i[A]��X���A���{ޔ���V�Ɖ6��z�s̲̫�iޡ��D�|�`�������F���a7�[v^m�Gۤ��V��G�����U
i����k;ث���"�פzѻ5Q+	�aܫ[�p�9"��2����b��
f��1@���=��lqЗ/8���>Kg��{��V�����"� �����>/�BD�
 �_�3c(G
���������z[jӲYRyw�,�%2@�8 ~���9\�K��NL 	��I�ygL�@�����^u�ki�#�}��8T;S�d����j$`��Ѩ�?�=��2�2�ƹ�^Z�VK�x*,4ݫ9�  Z�k�7�h&p��tZw�;t��|؎=��R��㻺�;)Y�`� S��D�&����'Z8�;E���%)_U�4��r��	����T4v��#�V0ʽG�C۸�ш���_p�B�M��g���6������;8[G@zֹ�B�[7}S�,�E-���4��á�������r���4�;�s:G�Ч 
y3R��S	}N����jR���nk�ąܳHk������UsF4���F�8q�k�X��}J���]���%��f����}A�Zg�yv#A>|��mHc���]w<�ws������<�z�L��g�fڥ{
�P8"f�*Mv�c����wH��qr�����tA�$ �8��TU��<�"��C0i����O�.�s9��y2�rI��Y{-��^����m�Ö��)C6F����X�{D�.�41�G䎑&��IY��m��z��e>��Ē�}~H{>��3����r�~|S�l��ϩkw�(U�9	�u}��4���+�!%�N�n,��l ���)6�R����=�T��Kkω+���I~���[�y ��(o��-��/�+盇~k��A�/A�V����愬~�D�1*�G^��+�/�n#�Hի��螞���|����c�����v��Z�_��o+R����s�	n�<��R�` &Dek�n	p��Bf��\z���2�Q:�p{���% �le�펻謒b�haL���K#����+;m��@0f��ͨf�h������~H$d�����op�şAū���߸�)�!���_x!$+=���Ur�?5����f��t3r*<H�bT��C�}:sY�.t����ig,�(�)��g"!C�V�1ۧ{�f�����S%�[��hui�� �Ki������c.*���h���e�� ��b��#P�U`���M!"FN<$�/+h
�q4��^p��� ����<��GS]D��8w�<�;�'���#�#���`�1�]a�F$�{Fs,Mֽ�?�y�Kk���]�r�{�0�*����af��C��vפXT�_�2N��U���p��6ٔ���WA좨tSo/�A�/cJ�јYȲH��#���Ƥ��z��}��R��������%�-�:K��+{'+��ߪ���0���:��Nq�> �"����՞MbY�/:���Q���C� Š �/5���U�-�&�*ykz���`��X �-��o���r`kN�����r�ewv�M�i���5G��Y��4�	�FN<1�\}yh��tt����!m��	S
s�hw�4� ��8:+|����#���mߒ7�c�Ō��3Hˢ�K�vU2�i�ݐ �X�Rk��wiC�?�;w�����t�n�D]����V�_B���3��E��5�z���o� �ٵ��Ar�kRb�"���
��Sta�pH����ٲ��_{���]��ة��éw8P��$q�鼥fۜ[���Q��|at~�Å���C
�$R;�[[R�Fp�`��T��Ej���7~��ha��X��Wˬ ůF�a��F���l�c�f6�g���O;}�*:����d+}
[�䜹��W�1�\�N��)�iT���a�vt��ov��}�Y�Η�g�"�d�@?u
߯س���y�xy���W�_Q�����0��Vp%�݃yТ�nX�9�vV�q���_Nۆ��hѭ�"~��ː܈����do�tu!�8} �X�T����C���+Z.wE5�TW4�|��<��h�l����ܟJ8A^Hc��{��Ppu`�9���z�e��l
��Z?�;����N � �����oL����ߖ;˿Y���H��d����(����$1! �_q�^��v����B��%|���ꈇ��{;�h�1��ԯ�J,�쀌�)-zI��R(�/�+�m_gٸ�	fn����5�
�F���Ԙ]�,T���o�����Σ��(�ɱ]N�������÷\2���'��`,U����L�$�Ǝ� �U��Ɂ{HD���댆؉;�qW�dD�U:�QNM���bZ�n�qI������8�h��`��5`A���7�>�p��Wz	4Q8�>	khޗt)1�q+�k_��A6q�N�m�=���]���o/n#'�;*�����٠�D|c*���{ܦb�IC����ga�fSn0����c�]�����tw���Հ�w�O� r��>�Ja���:��x�f�iRf����_�ZҞ
/ia��:�rF�2;�!ٳ0:�t�	,[�v�L
Ӧ�8���|����
�c�D�����T��N
���5�hM<K���}���`A�&��8H�"�ʠ�����B�=>qs��7���D���8� ��4�V���}5l�@	�� :�CqQI�\��+��KN(�A��o�}%�O���)��,R
�����/N�+Xg�{�x�i�ѸD{�}����/� i%NrV�÷����7vS�Z�^��u�.5L�㔷���*���i��ˈc�<_�;�CbxT���]�Ǝ���uV&�AaaeY��kG^Z��p�n�g(���V���
g�o���a`��k^�x}y��eoP%|.� L�$����\|����^�[�s���A�y�� ����82�پ_l4:}�R���r����ɠ���Y�a�x:q������9��H���],k� �AnЎM/�#ͩ�I��������W�-�w���K��2re܉H���`��u\WZ����Vg�兝��f{0;��5�[��1G{>�����YO�׻uN��-Z�h(�����С[+���v�Eokخ���n��Ĵv-9
����@<�+
���sl�i����EMn'�_��|7b�Z�L��F�xY����|������{�k�~���A�?8=�:�]4{���e������K�:Q�=��=}Gm#l��k���|%��G�vvv�z:|�����w��㘍'�����w�������J�-�.���z;T"d�7%�}�S� ���g401���=�����U�U�]z���C �>���
(;hHw�[��F��^���a)���$�u�G�u�sQ�����T5H����j��_�t7)]²X��F_%׹N����/_ތ�;�x3_�J�w���������WwT��>�!�7t�� @�����%�vԟKySh�͏X^����� ��*��2��A�A�%ŷ�ݱa�ۣ�n����^I��-h�}��Z�wz_S���?%�a��(7�]�`�ي..�/���a�mK�[{4�:��Mžx?�<���#�xÏ�qm��?Uj����J��뚴tGVN�l�<lDt؛'��Jdrk��ޅ�oJ��pq��l�ר��siE~0;��0�3Et*�}۽�(��Sr�ODN�+�vt����;?rˈ]Y�g{ga���q��b���{[e��z;1U�n���^��`��}�Y��j�\h0�����A[�X��Rc�4I�9k��k���ұ�xe�q����_�泒����O�GG��I�~�ȝ�G������
��/~>hKn� vڄ\=��n�o�H�2u_g�a�\�K����l3̛�!���֕sʧ+�L�����N�
h�g����CU�>G��dL����ElxmAd����u�\��[��Q�����Z�J*�.p��qH�h���Ld�_�!Vő |�D($�-^�j9nSw���Zؒ���q�����}�%o�{�yYp"�Sz9���|VS-�g��~�<��6�j�?�}?F�%��G�R��β�5�Af|��N�������A����JN�W��M�/e��˹7ؿѨ�ڎ�^E��ѥXU��!�^־o8�ۊ�R�2M9�,8�d�8oB�V��y�N��f����sX>[Y�O�=����$h$(��C@�T�Ց���N# ����>4�b����ҏ!Dl��X��ְ����#ļ��&K>T�n���JuoR(�%m�)�x|оų?i���uo���/gI�O]��!V���b���^�o�PA�{+#(v�%�xb���xK��W��T�}�,c8q���Z��U�������r�o�����l����8�fc<��/�vQK�If0�^~��V�Z!_�ߴz3g��]�������?F����ae�Ōu��|�m�8/��,7��I��atC�jl���RD����_g��QI�:_O*1� k�ɡ�_�r��p�s�����ҟ�1a����u�_H�o�I�����v���d	ʴ�w!����W` �O����k��Q���BG�Q+�����x$�,H�4��켱<|��m/�Pp�%�?<�����JEN����+%a��5��2�Tl}��zK�:��o,O-�RҐB�X�nn����32Kx���/o��xS~��0N��u*/�*��^U� �%3L_/;�3{^�M���0+�o��E�j���:�s�j��ls3evM�xY��*�t�
%X�5g��\�a☽q5�O8��M	Uǁ	�w��9sBYu�$��5�}ِR.!2�\ۻV�;�_?��cr����A<%��`������O���.��~�͎#�"�m�.�+�c�]����@�Y�!��Y�'��׭Y�#�V��$�5�)�ń�^f t=b G���h��Rs<�:*z"����lR�ubc,�L�:Q�z�8�2/M�ዃԴ���>eϔ�%,�� ۬��˹�C7�ѻ �&���@/����[��͆��*��PM��5 ��!��������wV=���Va�;K���BW��µ�i�'�T^����2@o������G�Ea�B\�I�&���~y9F`4�C|VCTރ�ăj	��G~:Y(<s�"��8�������=�-$ht�SJ�ݖ�@��4���/�
R��:�!Sn6?h�p�,W!e��yh6-��r�g���Z2z!�!toKAEER~ԯX�]�E����2��i���ޣI��WDfddy�{�v,�1�� ?�}�Mu�������=�ھ��r�THn�����w����0B����Y�pY:^A�u��<@ird��x�D {�q�4/�m��U�Ny��?�]^����D���,���%�"��4*U��hT��CW5�HK��Ԫ��6��ׯ�5��7-�*���X�J�g]�`N����$F'4 "��L�������� q�P{�[}w�\rW�����>{vXie#q���t�췘4D��Ԥ-�����3pЎ�ks.[�aȭȵ��iU.Ґ_LHQ@�>���'��)��%��,4/`]"��~� �]�I����gtJ�0�M��ta�8��-����.��g-ঐ�hԛ�4o��� ,gѨ�b�.:�}Du�zuI���S�-{�)S=W?�~�c��`sfDWD�CHc�=! ��K�Lʊ�r���e��*�J�}ǟ�}���N�Y�5�?���c5S���=⺇&�O�U�p�y����0�IrTUq�V�����*�~���jXxc����/�&t<9�ve>6b�'֊谷J�>ת} �XM�35�8�i���A�2�I�>C{�X�E ����C	���&��=s{"W(#ino���!��n�`�sH��Ǝ��޶��]"2��X�	�~�= ^X�u�'W�vk���ɭ�����#���nZ7m�[FŇ*��r�O��ʋ��3"V
�*��e����Ұ.�����+�8�G]Z�KǍ��yc\���$��d�J���Y5�6���F
�W\�+, ^g���D�S� �Ϳ��U����J�wCm{�y�R�5\�I#�Z*��M3�Y%=��|�u�fc�LD�+�c}�.$���8ۻ^F:V��� @c馠���$�c!Ѓ����k�J�75��-�(�DM�14t��;�Q��e��G���Stf�i�[͗������Ҙ���u~���>�-.' w)�����v�`y��F׷��(�h��,��}%삓u>Gkm&W:��1�<�@:0'��Nl`I�g<a#�̥ͳjq�i?�g˫�+Z����tʐ�`H��37?�L:Bc���I�Y�,龠�K|)v����Cτtaq�|�l�����]k<<[; Y�^�F�nz_,|4�G�ڲ��@���m!`�,0'��/=���gA?��y	㉟(O<2%�=m]7���V-mUm(��Gx*��D��W�F��a��S�Q��)�_[5i�O5�,)���׻,S�ؓВ2�V���9�ZS7�rJ����A�!l�,�<�V�w3��J�P�l����w^�,��n�Wk��_�mF�``��R������Y�����Lȸ ��*�:S�Lk]�R�@�;`���tݾW4�}}��\G$�:��J*@�[-�F�&��Q��2aB>�w��7�]VP?����c�Ɣ�vy)]R��6���8��\`h�LV �����%�{߮�}�fǄNo`��#W�Z�ɭT��va�ِ��,�3i�A\�#��Y�Iǧ�Z�I
7�!��I����\�=��Q2��C˧�I?�AV�\�d�F��ԕ��1cH�ci�is�$��V���ڗ*O:m��J���tیR��\󆐅��-%ɵW�A�������ʮ��
�#�w g���!���ӵT��p�Wi�չU2��E�Z�ͧ{ ��BO��_} &����/�{��3\G�HZ�wj�v���������T���X ����_P���ا)�s}�o8Ɂ�BԼ�b�c�uN�ۖ�,�tf�ս�.��>���T�?Kh/���3���t]���1�>W�{Ը9C��i�{��e������=������@��G_���EM<r�&�:;��5�	� ���v�v�M	�v��IG�Y�ZTL��v�F���Sю��bfѦ����J��H1mI��{�~��@�o�|Ft�Ҷ��Fg�� �Ȓ+wj1�,Gx*4�y�L����L�_mEO,˷Sh>�O�Y���ٱvYd��h��>5�[Ӫ�&�[��I�����AE]s�&)I]�����߷���ٓ�<�f��p~��� G.)I��Ƴh���J�E7?Py+B��T-Q�-���=\��.��;	U���XK���K�g:R3(?���c<mj�w,��X[�wG�I\��밴�Y�yť�35�N�\��M*���-{#�.��W`#�M��pߍ@'�=[/���Ή�:I��n�&���K�U_e��d�g�z:�B���Q�{��m�7��5Oכ�ڧ$j,}���/�eNl� ; �`t���T��'��0�s�E���h�q�lY޺��=�%�'�sSK����ŀ��E���N}���ܲ�3Å���[и��9t���^�,:�hT y���Ƿ�u�?}Ab��b�gU�G�E�X�K��v)A�	�eҘca���
g�9�=��[�$=�H��^T�-��E֗�9w�H)��������Ti������'.U�B1�ӎ��z�|d���9���1��&L�O�P�?P3$h��r*C�� `�G7�(՟�(�������bJsIN����m��-�	����J�������~I/4/��|�T�Bn6���
>�q�i��B�0~*��3su����&�t�C�5H�j��^�8�뻇�֮AC�����{c������ҙ���F��%d5���;������n��v'�7c���γ�>D���1�� ٚnz��̵-�4�S���}r�?��nn8��MF̻��ʬ�׳�������O�?��WD}�^{��p�5.\�Gx�(�1\�P@|鯉<?�Z>Z���u��Z;p�f�����y��B7��nU�R��8B�5):�/�0�m�v.S���E\8�������Z�Y]/iG9���
�=Y���tS�Z���1�\�Ƽz
�j��+
l��2G���i�'�waj�?{���T}��m�3`;�Z���y �$����Cn������w��	&�b��
�e]���6\���LZVn���פ%�eu�Q��f?�vCt�a�ˉ6�.1�yK]�+����m����菨�QP�yٽH0;�[�0��T��/k��G��%t{��{�ԻZ�u�y��������'�1b��`�lia��і�l�"�ym�jc�֮9�'�rz��zC�u����@��q�x���W~��^e-K��<���5�j���1�����:ܼŨl��˱l!R��x�V|�b�̸A����60�e����DBٶF�� �4����w��C��C1�dS$��e��.�?�_�Wiw����To����&��pz�˽�������Ζ��Z�Z��O�!Zo�f�}��������<�-�"�;^��`��fU7%u��P���UTZ��W��]��N6�xX\W������{3M��^o��VO2�,傣�3�9rfM��&R��er>�����a�@���P�<8�f;i�dW�N��
�����߿+ '6��s�1����<v=�Ŋ�]L6Z?`��;��}xfq�T�'�ا���i���!������?��`�y&�l�����RUhc�#��Z�u�~%����l���?QG�!\m>c�2_�^�7	kg39��'�KI���1���99���)7���s��}�`Ϩ���JN4.��5�"�G�ҋ�t�Յ�3�#�%���(��L�$�X�DN�Oc�V���M�L��>�8({�eR��I]��XO�����r4р.�%��w���Y��e���"�I�NV��'�p�7n�����\Gm��� �^�IiT�zA���>��)�#5'}:����n��壮���G�l�J�ŧ���	OT���}��	 M-��Ov>����v��b��\�q�x,Ԅ��e"T-�+�n��[bq���헄.����)7峬�;$-,��в�W��S�*��.��ie�*�{-��\b"���ɧ(/˾���[�ѣ�[����MzB;x��'�́�'�Ep閸&������_К4x z�~0:�j��R���}�+����)b�z�,4[��;�tc�^��..k����Y�[[��K�T|��r
D�%�8x}]���T��񝸬���ͅ����:����o�0W���<0���y-�G�����C�M���]|�j��E�\!�	S_"���o�KȤ��k��f^%V>��ʍ�={�5T���bتu���پ�٪�2(s��?���c�xs���]�T�I���W�{�0[��v@�K̻*���Q������+�!�ME��k�.ʛ���kk���$�͂��Lюr!=��0(Ml�z��>Y�'r&��G�q- vӗ��"�_6��V�4/�M¨�_�F*� ��4
�+��5�ځ#d���/���P�	�,���˨2F�,9G�>��	��$�*����N@�[f�OD��أb����/W�E$ptW�]8/)_~�x5���?��UꛯI����ʌ�|l��Zy1���|<��œ�Fu+Uy��}���������ݶ'�m�}���y\�c�����㠺˘ψa�C�p���'�X@�_A\���W�w��h�8�d/
Jo�-2���G��F�U��F15��v�(j�xk[�u��P�$�8��0�^w"�}�Ԭ#�V����l�u��Ɋ�~������d�'�UvY�"
l�*��S����L�	h�9��V��ѹH�T#��n���Fgy��� �	�#k�-���
se�H�v+�ۢ�uo�����G�vq�O�;��)EJ	S%j���}�l}�[�v>ʪ�ؾ�f2�0���T(.^.K��-����T��eb_���W�w����zY�p�I~R�b9W[E���ӄ�f�'��R����B��_��Ά�D{��u1�jO_K|�K�"��(�I�G�c
t�'4��yXXئK��Z���I�:����9YC]�o�2D��$	��������a~㙓kQ���]����ꭅ-
�E���(��j�f��m\ng��σ�e+�H峮�y#��B��-�p�!�D?ǧ�KIE�5�٩�kHҺ��-IC!yP�2��<��RJ��:x }���#���gj�u�W��3��Z��~�2W�G��.]����*RVr+����-:��	q�ۭ�ڛ�N�a�Ĉu���V��,�M^��Ar�\fO����aZ��ŗt���D��hXj����	�M`2�m=�
%��r��?�A�l%L�fUS
�~m�Cz��m�N���OQO�~�P$�f9�s����Vn�E���JQ.��_J��ɨTǼ�u5;+�6�Y[�>0Ę�����ڐ���)��z�Uᢑ'�L��Ed��ϛzO��c��U���Е��}��q��rJ�cn���=�)���r|>՚}Bw5��u�y�]�T�1p'�G�1��Q�n�?��H����zS葊�3c(�jL+��U��هk�+i��U�<`[�(�Q��}��5j�4�~�'ٗ�s��废A�t�PߕlM�D��	!E%G�rڷ�I�v�C�E��y����?�z���2C�ͥ)V�dU���+H!�ո�x3W����[%��p�?�#��Ӗ}�+�@���8_\1��r@o�X�N�<�`�קy�7��Kx;X6��a�)ÖI�����~�����ʖ��Ľ�������f��eO �_Rt����n��~��}��q9lnTH���SO�v��d�j*�<�8������wnbuR��Ÿi���a0+_b�a���}db7�+�L䰗��i}Ve����P�><~�e⫇�uf����[O�H�����"�G��%,.گ+V��0&��j�)͹�q%^k�$K��_d��>�"��,vL��M2^IBr�n<�8`�Ky�������_�{��O��S©�j�E�Sl��d��}5��]�� ��0���f#�ke�..���v�/%�P)��3ߒi�[���7���~�Gİ�;����8�2���_�1zM��tg��'� P�}��?��r	.`�ڎ�r)8#�aG��#�v� d�;���d��;�R�S@��Q_�sˎ�\o��Vu��~�1;7_���u*��Lb�_�,��S���M%c��Uh89eIdcz�(��rM��q���1Eͦ��v{:�6V��,'M
SÕ�7,_��^ͱ���F�Y�^��l:�%	�'Q-��:�,����)���n,ͱ����q�;��>-�:������Q��T/�1�s�̅Z��j�O����h�W
|<������"Km����m�p��&m�Ş�2�ޘ+�O:A*��ܵ�����Z�K��2��[��6���O�꫉���~x��F�3�%����F���/�+})@��u�z���z�`4��}�^��I�PS�B�L�(���:չ	Z;�����?!���=R��ײ�3���e�59m��
׏����������)��K4��v,�b~E�A7��ܨ�0����<��b$m|�=�ȝ�I���{�?�}�J2��/α�#Y
[���$jBx��GCO�.��β����P��!Մ��#�{�	��>��|�5���&��Y��L�oD0R��
��Á,��K^�ɯ
���e�"��;�ʞq{S�r"�x����@�j��H�����>����M���.�/1��@c�������<���ѾE�q���=Li�(�v��1Õ}6,ֶE���U6�7�"/���Q��������Nxu��"�oiR�F���lD8B�d� �ޅ[���^�k���	�?Gj��"$z١���b6v�(�Sr�;��o����Fp�oWKDsL^�=�u��q�󦉶�FF�$-�(�L޵J���o�5�f�7�דeؽ��^4߬�����+Ionc�������[�<���?
�ƃ�̫��lm��%c6�M�Qd��
-����E�m�͘�:P��M��.6��I�Ƕٕ�����>Xat�.��_%��<���y�x�*�7e*Lo�����⥅_K/�������?�K/����5�����fc�|���Jl��z���#��>��-��]�ߧ%�����U-�Sz�I�[Ĭ/�뙬�ڧŵǷ��b�g(3�e��/����C|��g�(�*YN�ɍ�4p�|�����aܧ�V�����G���!|�q����Q�ƻ5����j6n�����l�u�D����?����1V_�R�&��F*b��,M�m��4Q����B�_Wi��r����[�z�1�2k��[ҡ$���s��aж��(�.��3���)�Z&%�	�_O4�#?�������t�80?d~�� ���K�MZv՞X����[��FG1���{�-t���fD1nA�����Ȝ��fe@ob�����}����M�����n}���7��茮qEG.+O����$�\6��,�W��c��pD<����,���,�-|kNbIm)�oo�DgV:�~+H30H��2�|ﮇr�Ӊ$k��2���Մ��5XcO�`��l頜�cj�e�>���8(���k�ï�l/��bR�����v����~�m�,=z�hl��r<|�5��K�#����u���$�̴�V2��Ts��$/^>��A �Ee�ʷ��^<)���\q<���S_z�fi��t�|�o��?Ľ��<�U����S#a��OU+����^s[Ss[]�2Ӈ�z��b�k<�5�֜K;����Vl��1cg �x�f������/��p$6IŘ�*?��Zڏc�&%�+Z�+�d�w���g�g"O��B��;B��,c9�����Qiy��Y����0|���xjW�^�[&���*�҆��'?�]%�A����n���z�U"M��d��.�<���xy2�[�bk�ꖄ"x+�دl�*VhTg�s'������\���A{�,	Ω�$'U��b�C���7�ܫ2ﰜ�4�S����=����(���L�QJ�TQl~A:�CϦ��["����'�&>Q���#��9���	Ӧ��m�����!��?��'�M>�\��*�E�[��f�
�0���pW/��I,���٪���)��4��QNf39t�XX~f���r.�ьN��?�M��3�K�4�r����a�=��j۵�(�"
A)J	AE)"U�%
*���(((!@B@D)BDZ�""�� -����$!@H�y�������������c��W�d��9������yDpg���Ql5���.|;��I��nܶl85��ϝ�?��q��R��j����g�T����E�,w�yFG,Т}�7����.O�8eic[9���!�P�*��2��r5*����A&��Sl�r�?���xA!�D���oF44&U�TZ�5<ٗ�b�l���H����aO
��l��_�ʊ�z���v��*���_EKҖ�)���e��.��c�%PK�Q�mT��n�ȡ /���}�'��{�tw��QZ>�8��o�vɛ,�����0�=����γh� ��~��S��'2�o,zI,�3Z�W���e��]��p�O���/m�r�X��+߂�_����7����T�Yem�:omM�/���s\�qļx0h�c��� �Rƺ�
Z8!�r�x�U���*�a��@ϟ���]l�;��G���ބ@�.���ֹ캏��s��g�A&JF�M�o'T�gW����_p'cO�}�NL觻���G6��>���|	Q�Wf�.FChQ��O/��kD��K���~l��b�� �yZ�0	NQ/*���?j�a�����{4����/���W���.@�h��D�oF��85�(/�}
��|��ኋ'9�~�����*sW��7�P���H]R!;T���BM:�����U���ej��S$���c�� 4��0�uѻ�׮qs}�w����~;�C�C[-�����5ܻ�M���6���f����� ?IǒB���)�֜����{�O\�YՍɆ9��μEbk��ʮJ�
��H^d����s^��4N���v�.լ�J��ר]�[��/G'f��"�,��~��nj�քvT��Ub��_��C���dPb�����ܸ�����[K�-^����Z���,�����%
���d�j�Y�jL�eiP��>z�9������8���O	�������d��Q��g4������&s����,=`�ƶ �bXe����d��:���	��B�=��������I>������(.����K�����?�~Wc��oG�+*ƉsN�k(V��Ҟ�P {�ج����J�g�4?��1�I���8Q�A_���2R�>̓L��*�C��Q���3�A�ջ'Z�c�j6�滴�]K�o�ڧ�d��%���/L�w�n>J�
�[]��j��[m�O;�%���ռ��
	��h���'E�`���Ȣ���=�� ^w�
O(�����i-w��L_��3��VF ��� �7<#?X�$k�qh�+b{y�9��N㶽qY��o��1�' �=�K�r�� ���삊�	{QQ?d�l�`�_�)3\xt�7J)Hd�T���X�1����y]1��hQ��G~\�7]����n���_�C_�n؂��޿�F~Px���7?P��fuv m�����O���؁�������B�k��>�f6��Z���o,�?|x�#����ѿ c�u-���~-�&�M*�i��qg:"a� 4ϯ��4��B�kE�=xf�2���2NѢ7C����@$A�(�Ӄ��¢�����A���nCg����*ܖBx��PT�~&V�89k&���{��Q� k^�Kj+ �S�r>G$�Ŋ�$��ڞZ�qo��/�OE2���f?���9��	�o�G����Ri����\6|�'<!�ff��'V0��|�܅�TO�d8�xj�Ե���ÜLTI0��'4Ν�*r�\z+B��4��ૹ;�$LƯ�Q�����i>�#�
<+���{���˔Ou�M�{��M���r�G�O��.�:!��T˞��4P_�;�L7/��`a�5W�AI�-������xB�H���-�e��P�ƖXN_1w�/�	���jY�a'u���p���+(�[<��ST%��@�h��6R(�+X��CW��?i��B�h!q��49^�7fh�@���=�E!�f���uoӎ<�	����M��w[�o9��y&�*�&��\��5��w0�H�-�Wz�zp1���ڲz�V��j��tFq ���E�c�p�$r;��a��1/��>ȼ�E���+�Y�k�O:�K�74&���kr
�W�ȣ ��3����JXm"��~\��b`�~�$9`:��S�~�_c�9��?g��wo�9�B�i*!��s�_��5}o����Di��}����}�T�� �a�C�7T$2��<j���i��)�}
p���oy��u�fa)0�2	Qi�~=~8X��7NeW�v�	��X.i�i_�B��`�������o��D݂���#���n�;�n�������=H�6W�0��� �������~�C�����6�l�
8���m�>���M�9�m��l��%�ő�:ҶaM��������2����M��������y�pj���:E��>�.�T^Z�B��ޡ'ڱ�r �C�5���z��}yH��\�O��.�Bҝ9oH4����SJ�K��uUwn�3YC�7���K{��M�w�Ԉ�Î�]�:����ّ����5�V2�bI!Ma�hg����vyO���Ϲ��Ҙ?��J�h/��Ҟ��2�k����Qq=�����bK�	�Ӏo�\(��-#Ze��j�����~F>�V.I�M�"����-A�7�j����s����ѭ#�g�	��l��>��{P�O2��;Қ+�e�D,�)�2|3�y�91z�$}1��z�tR����E�	G�e��I��C�c؄$�J�L���1k��woh�Γ�E:-�} ��������g�w�����՜ihu|X���ʼ �Cp�����;�z������8�0A���|+i5�ڧ\��my��E�E��u�8����\�s-�}���w�I`'u�*z�=���v��֬��#[�0�u+��(�NP��+�}É��`A�_F��%������E�&����L���_�o�2`z����2��8�5�g�/�VZF|Y=� ���+�W����4����Ѳ,����gz^�7��z+�2\�J3ÔG�?��3/p~�ϗ�S�\�US@�<<�W�Vwt�=�&7�a��M�jT�W�$V�>�vw�	o����[=҅[�߲�H?>M��|���o�E).Z��#���'9��*����ZҰ�|:8q:��3]�4�"OT��@Zj����M�3��cdP��vU����k������Z���`����Z��y�����-�����^>p��U�N}MXYH�u��M
4�T��3�֚|�e��><[��xO�w��-�}t'p����/�C�T�fOv���
���!;��&+mY)�6r��1׫�ʚ�d\�+:��-%,{��̔���IV��.��a��C�t����J�%��ҡ��I�J��Ѯ{z�Jճ�q��:�P�ڕ#���e��;!R�W��&J �u���u��9hE����S�{�<�σ�� [�`�Ka���&sw%��Xz�_F}����1hW����[*�_g��<�8 ��m4����P7T���j�%��0=���y{Gs��}�Չ�K�����ȟ.��8���L��n#z#��ǧ-��>5XێK6ue��gO׋�
9�ҡ�W:��'[:ɻ'��N<4��� 3.���:N��k�����:Q���v4�r��<��C�b�}�U�\E2׳�B�W@k�@�C�/-�Riu~cR�R���$��2�+����AKv�{Йb�7b�����g���(%�x�;uk�`�R/V�9�Q 0��Ew��h���N�Ps[2�7,�G.���m<��˻�h�j8����e3E�utK���ÁǞ�z$��L����d<�h�?[M)��[�2T�n����d��8�sH!揀����6'}���:�ݔB��$ɵ����j�pgj���a6}U@�Vkқ%�}A0`�������8H�V�+�Yc��hʉ �p�/�����f,ph�7ɝ����!�}K������B�J����gVM&�5��\����]��D�?"}���gYI��t��kh�V�jJOGI��#�6B�=*��4'��i���[����QI��K;.�U�VCl����U��>����ϑ�-��5�w������:X�hl��M�Zl��T���48w��r`����jt��q����;:STҵ����%�m5�[�V��-���f:�<����{�:\�{�5DZ�:�����.0��O=�����e�7*G��Sw�Չ�*���3p���!��}U�ǥ?�)4��N�tb��..��⿄��I�/뽱_��F7��'N�LoI��kvKrǇz����Vw�^�&5�Jw�W�D�(�sQ�-/��<��R��l���K�I��:�1h!���$�MT�=X�B�鰉R�ԙ�.EԬz�7��� �W������G�����5K㶳gֆ${�KU��N��K��]�a��Zwe��a���a�ف~��<��L}��Ç��%u�9�g�e���Q��,��?2�������P�k�/�����`����7l�B���p�����;?�i�w8���އ����(I��V���H�{޼�z�����e6���ґ�o3)���;��ؘ~NF�Zr� �|�?r�_�� ˞	��ב���Q��4�wQ�9͉_O;�:���N��ܓ`�l��q�H��9z��o���A/�Ðl�ܬ���>�]洈��2\�D-jS[Dҗ�p��կv�y1�3`9�#p���;����I������Zx������y|w��y
?�.(i��/[V����U�&��'�)�6÷��q���í�:7U�7�SA��O*,��,.�*~ѥcH���gw�ӵN���Ɵ.���Q�VPZ��=y���j���>8�bg�
�E �3w8���F����Mi�iH����r��^��kIؽ�VB-ֿ}wK���5%�&''B��Ů(�L�s��~��K�Q�Y��F�[>&c� �7�����m�F��'��U߬A�pw�W�*�Z��z�-a���W��Z'0ҫ�U���ʸ��<��\J��&�d4�g�s�3t�A����Z��ƘmE8����b���#x��~|^��2�v�JZ޽sLϑ\?G�u���,����?�(�~מ�4���6�i�KN���g����6�2�nD>0��nk����i�։�+*&�"���?L|+릟���R"�y��o�H#8��^C�L5�ة^�]Q?�9Q%*b���".%	��g=ғs_�nVw�A�֡�
���Ryԁ[}���UҼ��{�B����Cb�HYn\�� 8�j��|���@��1vM�*])L���i,ΛE��dDGE��w���O��e����k��;��]F���F��W����K�l�G��x]���5�Z&N����6"Z�6�d�_F%mY+/����g�^���^x�7	aa��_���Y������ֈD�9:n�)�~	����O*[�O�VA� �,�����+�g�Uf'�Җ�^!F�Q$��!eP�����Ԃ�Y4��n��/�a��؁ܾ���h�0{5���I{֚��`FL�ר��%[s�4���d۴�n<��x��lu��B�Do��p����h8u�G	/���F�I�aWT�y�����BW��AYo�Py%��+U��8*5���lf�L�_i�t!������&Qk��EίR�;/�a�<"���Yg��R��Frx.C��q����{-�<9%���5��D��/M1ZB�L%Vx�r�Ϟ���c�|�-4�`N�xפ����;ARp��]����c0���am�M�S;|iM�>5^8�3QX}ٮG�'6����p~�ZxY�dt��j͒�����r���Ȑ�N���J`��-dNtK�r��\/���3Ȁykm�9r�U�1��Ƀ����9�AWF�_�	e�t�9��Y��+�[F�$�,�`���s\�ϑw��B��+���i���Êq�X�媐��$��:��(.���L6���jO�/�ЍhuH�Oz_��� }|�I��=ˢ����#,I��FlJ���=XX�Er*�l,4aRT�3jh��']KK6�?t ��Zt�w�F&�$�g�d���<;�ĻɌ=�=���<���q3��l2������ˍD���۠��8zʃ��´(��g���zUnD+�Q0�v�j��ރ',qJks�7���} �wF��%�z4a�'+`B��'���,���9�
�b�ի8ߡ�W�Z�xtn�L��X7d����:&�#��u�e3?C�e\����*�G���)�Ÿ���I�*�X��N�{�(�&3؂$��B}NK�#�ƼC��e�z�;�V+�S�2���H�(<�~�$[�vI��'�1ܸcV�=\���y%4"
�0�\,X��n���Ø��������U99˳��C���Ğ�Y���W^b����[�f}/�q|��E�D��A�&$��u���*|��3����x�7�9kWѧ���=�=T���:�bl�������e-N�fr���:�E�$v��S5K�L�p��#���jY1�P��{�/>�	��*�*1xi�>������芈�N�BX��^�q���0K�F�33ؑM\��J�@�-��i��`�|�"�FA���>������'��`e�3E!��g"��^	B�O��.�b���:�T�6�n�8jZY�E=r�� �Jp��z�Zw����ߏ�M��F�EA~��{��v0K5�����_1���������]́��%�V(L����J�vvQ�8{��|ErH�g�09�����x�{g�^׎�ݴ�Z��N���Q,���Uև����3<h� v�C�}-��V~k�G ?�M��\���~,4�;=].|>X��pAeg���V�*�<�r���2���oE��|�{�<w�a���`M R���/�{u���f�]�h�K�b�����29�`8����|0�UEXx��o�i�UՕG)��� )��:U���Fe�O�M�;��toŎG����FЖ�źD���rW�ռsM:���Dn�����C^�u�W<@�׹�m'��X�4X�Ҡ����7�1�V�6�H�����o�[[�U� ҆�1�j������i��&�o�H�ig��o2��L��x�n�෡���31v������!����wf��/��o�V��Y�I�a��/��H��+D�5�\����B�7v��D��Z6�5��ߵuν�a�qJ&J��@�9R���6�g��=�J����J��%�8��*�º���8�H�e��ٷ�s�,�~r�~����ę��x琾(:��kǃ����Q�\i�����+�vՑ7�)9��O�U�#��9/i�����b����$��m�HRW����˱��OPS�Z;ᗊ�T�7�J��OH���[Ͽ1̝�0Ȧ}���,'���1�TQ�f�Ɔ�k����<�|6����iZ�����d��~� A��:��]M�#��.��	I�ݐm5��M\^��<�Ǉ�	F��4�����î�#��fȇ�µК����(H���M< �����n��fQ �(����}���yȳ�'S���ۯ��G�5�53u�"E#�R�$��RR�B�n���?�pE6[��K�����X��D��#l�</${ծ�0}�ģ0�r�ќ��(���GI�@ͭ���,]b�TG�gV��j�+�ے��zt�u�1á1QE��|��p;�x&�y�'1��/�~��4�(������Vq����	��WR��w�,�"����3I*QGu�$�/4�]gZ�/bTf�b�z��Q^������;R�I�B�]�;=�^�<|2۾��ӭ���s�	t[�%�Z�UD�7�@�c�m������M��q �'e��y'�����\]�oz$k]!)��w��=>�Q�[��������=/���	Y��*@֯����ԫ�㋧�E��(����3#�24C����<��?�YQ7������#
����������|�Y�g��ݟ�$��<�	��[nK+)d��%�M����3��L4����m�i:L�G� FR��~;�Hpk�+�C7�S|`������Ҍw����?M��`�����v����� �&�K��C
F#�d��_n�/��Ō������k+�|�hĿ����7<F�s�J6#>Ι(�82����t��s婇ޙ$�І���7��5�4f��8]�)��Ӄ�
������ku�M9H����
�,�@U�Wl�О�8�}������V�@�*uݓ�b���8�π`���;�����7�S�tp��5���Ј����{`�
'Nk�F�W�C�D�R���C!��%o`9�,��'yQ�0#z����\��lu��g&%q9Ƥ���(&�����TBGǿ�3:�.q7�Gu�+�
و���S.���Ј��/�8h�mP�eؒ:�@��t�rg��ʇ��/�2A���e�♏C������>w�]� ��l��E�Z�F۠��h[S���W��t{��l��|`���pc�Qf�m�RkKj�x�5�q���=7�EM,3,*|ih ����Ո���?rKP�������ZC������dNo2$��G��5�z��,/Nx,'l� Y?�۾�x��~��i�NgU��Y��Bz�J�ajzE`�Q:���&R�Dvi�٩��QaUL�"Z!��:� ���d�w`(x����l2�b(0K��;�g��L�m:��=�23!�j�G�]���U�7p���ZӘ�f�A�S$�_�M�W�Q�o1�����n�_l,�q����4����ZSF^I\G�'��5
ؓ��V�ܓ�|	��JNo}g�0�k�V+�:|�&E�;:�H%��n�_�.��5Jhl�Q�)��h��%l�6� RhW�TDi�홍s.��˴�n���G�e�s[2�S�����*)T�s���тҏ�8��e��~6��}.����|<v��<��b˯��?��/�s�~�CA�I[����.	l��|����n n��A�wO"�爟 �z�,;:��PlyL��q���?�;P�|}���h�@����`(�!�o	�����B�#|v�<%���W��y�����ϧ��p����;��������Cw$A�Rv�Ҽr5��[���綷��	^@{�4�"��}
��no�� ����󄏷���܃گ��,c�K��Oa��F�E�i�옞H�3T�oճ��&������ez�#���<UM�)�v���ţ�Sv���y�ޫ^��G�GK�Z�Jvem:92۷�Fۉ��U��u�j�gK� +Ā}U��[^:q6P�+��"d�pdv�55���.�C%�BY�f�'���hF ����|^s����/��N�V�n(��}3�U>9כ���>�D"wl�� �D4@�q��Ѫ��e�3~��eS��"������랮/��9&XR�z�+i+r��/�/�D �cS����<�XZҽ��do�^'�e���c�e��8�^S���D���ӝ���Y��lW��/�����8��=���xF�W��"�+ji\U�HC5̉BnL�f��@I��dQ���t������r|��sl׳k���T�JL�4W�F�k�7���W1-�$��~�-��4٭m��J���D*_�t"֋����p����K�5LY�NDX�;4�9�/�t)E]۰s��@Y��*c�{qP��IHE@�O2�l'3�dh���t6C�NO�	��n?w�}X��bmQ��b��m�~6��"O��;��8d�	�/B��H�5�̺lXp��n̕z�J��;g<�#;�(_�ѝ�e���W�i�����a:�������CH#I".9�s�g?��T)���t�Q�[&��ͮ�87x�V�t�& л ��^��%���
�+�aR�����P[��pda�>��a�X���A���͎D�&Լ�R��艙p�Npu�޷�}+�q����ތY��=�%���ȉa�>n6�N{�ꥣ�Vr2�PF�}u�x�Q�BYcu,���e�$��bb0��&F��#�d��IF���i�P��0�Y2�˷����^~�f?	�[_:JdX���j+,֝(�����-�XY�s2r�t�"6D���[hSc' ��N~(['�u��_��Ƒ��k5���n�{��8���@���*9�y��w~9�`��^���7����?�&��G�~o�C�}2=��)A �t�_�e{�X�@�[!���Z	:�ڌ��ׯ�H4�ӯ�L����x%`��4C�(n�FUT��jy��u�(%�&'[U#�����2���R5o���.�	i�������I��� z�޹�#�U���E��rH6�?��-�3�0q9���>����u��ٖ������!����Z�����
/��W���x��	�
���yj��Vk�n�X�Z��J�|5R��#��s �|G,G]4�v1ڊ�J����,Ǥ.����4�\nE�w��m?���ذ��ao�i�V~t6������k��l��4e"�j�	��kO5j�K���?-�'n�^x1hG�[�[�5i���Z�G%��������ˮ�N�&HL��"aO��1�ڂ�D:��&̧��	�0��������e���D���U6u�?ځt8z�O�(I�ĥ�ujO}Yx�sAI��mW]e�=^��.��6� �*i�b
`W���v�0m�g��Xe�C��P�W�pz_֗<�fe��(�\����x��NT}t�&�U�K;��l��fВ)�+�/�h*��˞o�J�^.cQ�b��%A^��w�?�Z��f��*����i���k=]3Y�Y�.$��eO'I�LG!'l�2�����"x��P�]�'ZG�.(�s�8��<wgk�j�t�D����
_7��{�>_���ie��n2+��N򺷖N���<�8���S�$�\�s��ı�Isϳe���<4�?���hF�i��OR���B0k�<b'ڄ}��VN��t.؏���%��
k�t���Bֈ��+��M)z-�Z޻�^�W�L���ͱ�f��	�Cx��e���V+��ձ��K���CN�v8��Gq��ԑ��5���k�֡��X�̆@M���O�n��V������턒�@=�����TVuO��15��Ӟ}W�Q�� �ʖ
 ��z��:�;)
XYی� �p�>\�E&�N,]W�C6-������wm���5��J(\�F
�i�/�	���!"�{l�� N��'յ�Eͤ�=8����C�Ec�{��C�Z=���썈k���c�0d�Y��E��ՔF�_%]f�b:�;���`f2]!�M��p���\N�؁���?|K�����7���w޶��>%&fM弆}�֙?�#U��5X��>2@&d�y;�=�x��خCΌ�U�\1�&Cv"wBc0x���e�z0�oˀ'[�b�C�D5�ͣ1���u�0]DE�A
�S�Te��ޯ�����'�[����f�|=����Ǆ�D�B%������+�3r�����|Sg4�?����g��q����b���#H�=}�nq"KJT�D:X|�F|o�'ځU�!ޚQ>W�`@���Xڸe�a�2�X��Z^^���l����+A�FX�K��r�?�Y�D [n	��j?�肚�
m�}�풗��0�Y��s��k'���P���IƱ�����
ni�ğ�~,
�-zKscy��z�4��� �����!u�X���d]��#I��D&˽��r3�����S�t�jo�3(H��#�C+>v������9>�,��'Yxy�b.&�o�q��;>���Ύ��6e�ls�$�-F4��;����s��r�^�1=aKY�B(����C�i��Fy��g��JŸ���Ϯ����U;`����u5�B��&b_�Ϝ��.�	tO��eB��s�^��ib��0a�����=��u�M���i��摆�A��{�#�o�-��3�- �Ea������u��/�U��3���H�H�`3��.?�05�v�����i�W؀���(j��[z^��5�Z���ӫ�p�|��s[$h��"y�32�<�G=��O/" H��2����ѪOٰ�� �\Y��9_�(�I�a�r�un��Va��	{=p�)�Ӳ+�����%߲+��	�z�g��7S��'�sz����{$���d�K�CU��V�����.��}�
T��'u�^�^Ӵ9���]��n{|N
�.����>�%�Ql�
~<7��y؎ uA�)^`1�q����o{���R��e\�

O�83;M���Œ����Y$)����ҵ�3(��F��ͻ�@ux�r5
�]�����Պg��&P�?�L})v��N��L�!����'��}��
<�c3�E�,?�b�����vR�N����Ѯ�WA�!�y7�|V'Ľ����m\��2�j�s@9��I����Q����èá�� ���"���zP?De���
�utz�
iNfH_�Џ������+��ֆ� EՕ]-���-���K
<xf��i���*�<�x�UǥqY�FS.fq�,</��
sZ��A����ɿ�q��;%~��ja�b�2_��L���A~� ��R����x��2�W����N �5rsj\���4
�V�۴^kC��V�.!��ux#�p��댉��j��Bsh)�������էv�y��{hX\ ��x���V�������<��K�����w��򻶷g���I�E1����Fü	k�c��g"��\ȉ���<=�h�:��j����ؤ>�*�/�zv�w����lצN�J�gH�=�������m�[ZGI�쐯}��;��sH':��2d��v��@�9̻�qp��Y	+>�ʫ֟[$�aj�]�%8��Y�����D��(W�Y/˃i!�l�Ԙ��e�E���킽ǁ _!�X��fz������FK\��?!pn5jf�!w���Q*��F�,�tJ���%w㊁�~��Ǳz��n<j`�9e�k+<g�"c�a��k�n�o��x-���'��ZK���#q�5�8W�(@��_!㫡��}|O�WT7��Jf��̦u�=�0kl�㯂Z� :�w/�>��e�#ֽ����o�[FXI��b�$���gE�|�:b���n-d������F8!D��ٙ����uCQЛ3�{r?B��bLikb�2���9�z����$�޶%0�lХ���.�2�o�4��n>؎黊���³�fi
K�z\�9��u�%���%("������uq�]F���^8A=>lY�XJ\��p=P7;��U+:��$v�V ��w���p�~�:�\����؇i������ϊ�O^���j�.�{�3b:]�|���z�����'N�_O�Y��������I@�j?��3K|�1��N��g�rN�%�}��n�Z'�3#v/?�3�_�PQՖ�ȋ��g)y#�bE��ӚP�V�b�<�Խ��7_U�(��&��='�?F�����Tn�>Od�Ƃ�����=����O�Pu1���+'.��O����\��f�l�!�gLنO=�]�Dg�S_eZ�*o��T��^Ø��>���7��,٤���&�@ɏ�~�q:�TW�@Rnmki)�3��:���-/9w��>Ú�>���Z	c��(:����Q�.�ЗÁ8�O��[�hOe����*��ط^TF���c5,�_�f���?@:�ǆ�?��v\k}^=ӌ��JT���-_�6�mw|)���D���i��d?��{�]��U|��|�QDM���^	����MVg�����!���B���4c|��3�1`�գ�@ޘ5	�c�7���1#�Q|���ohbE��懤6��j�#�����&��_�G݋��,wE.a�~�q4�L\����2�7&�U�xp1P������P�O�S�����t�mڡŚȫ[YT4^�-2h�����Y%��G<��K�&�\O��T�G���x��'f�n������$���g����>���C`h�����E���E'��Q9�U�E��XOb�"j�JOD��!u�A.e� �-�|��UX$��f����K��΅���}`陔+���(�0�cXip��yt?��b�?�*j�׹��:�5O�s�������ϗQ�=�,�9q0���}5R@�Azc�����^�^��4���҉����5����K�`N�{��)�hT�c<�`���j�>���yK�<���;��Snms�@Z�r�s����ckAm�)��oSH�;��}�L>)����KQ�S�ny���T����u'f�z#ŧx�<$��辳����[5�L�s��>��6{�ۖQ���O??5r���)��c90�`*��56T�P¯3�K�3t�<�W�
ߴ'�/T�U�
�{�IMi�y�Avn��U|d��\x ����'|h���-O����*U�J��G�'S25j���9��GC�_xt�N��RԈ?����gV��V�a]�q�u�ƠQGŐW_mׇ�S�i���|`Y�C����"x��=�\S��tZ�������N�R�<bV�k��s�H�1ZE�= {�����1Ԟ�u/'P�c�T�VR�vy&?�kʭ������d%���X9H=m�5��q2��JT�R=n�ƀy�v0��6�f��A�GE%O/yHW��+Z�.��d|��$���vɉ��T�~�L@�����(�x#sI��⟺�����h�;�31R�_<}��zIz��V��&߲��2����i�1��9�#/�w� ߎ_9��4�w���	O�KXU)���FBr��ۘ��)�g�8�Q�����"[��oXK�$6_�E���x��T���Z+�l���K��:�VT-�I��y�͚)��GW�*����Fe����y����<N.&�P���@#AWJ��=S���eiAVoi"F�v���t��ƾ� �M�Z������)���33ʲ�{�]��qϳB3��v��{ó\�F��|ĩA�ZC�i_:	�����lB��۽��B8^E1���oe_xO�"<�8�}�������MʔE��E>ɂp]�����z�������`��Φ7�+��:�/�@�2̬~�;����Bl	��9���I�����ÿ��<>V�1k�uʼB�2���^��<R_��yRג.�o�E�M8���V�bF�ĕ�'���~B
9r8d��xar�}�k�@���'"�P���j��ӛ̰΄�[� �b���\���E����Y��$����nC剛���-��%���C����C�1�7���G�_�[�e7}��[�K+~�U � ���)C5A߷�jִ�IB�c��)��-zkX����-I�|��E7�R�j�C�*�gA��yA��_ �u�f��O�y�|�s������#C+f��=�
}E7W&>o���~���f3�ޓV�8A��=�M=8Ŵ[i��r`�~�����Cb��!q�B-���-~��)�A�(�n�{T��j�C[X�f!O�7�)�U2=8)��J��}�T�͓�R�M��X��OT
�.jj���Z� ��K�5���9,�FY�{�������??�Vܞ����謭�V��&1řr�V3?o#}��F���:�g��U}?�eww�BY��pw~�_="�'-R�_\X�um��,����3��T�ܖҟ�r����F9���~�*4{~^�'��\���PZ�D�������a�0�tqq��VC�KTȹ�;^�x�g^T��n��x��^u��߉����5o���R��d(�&��K���|����닣��L5W��rJ�����P����Be�R/���8F�A+���H߹`�L}���XW��_<�Wh���wr�W���
PsK��l�ܙ��1,��3+�^M��IN�a�{�ٝkV�T�s���!H�M�b8����Z�����q�}¡\�Qs�Ĉ���0ʼ&ETa�SsT�"%� �V͈�,�|� }�&r�u���=�s����P��H�B���N]LQ��-]�⯌�R��G[Q`��we/��u���7�'�������7&����5i&���y��� �^�4��G[��Y�5����׸J�b���2{I�T���������c��"���F.�{)���8���g!g<�*!��d�f��HE�fQT�_F�޴���.3h�i$FSic���~Y�Aث� _�6�[��i}�E�9j 3[�*,]I|���TtIv�N| eʛ�P����Ɖ�A�8�{7�F+e���}�-�n<�$>�´_,LY�M05ɷ�<��>�M�h#o�&rH��x�R)���U�����	�͖�©���nxy��AJ��Y;K���j�%k�R7nx�(�l�u�K;&�n��D��r��5���B�n�fI�p?"�c�|��N�N�X��{o22�u�T*ұf��ia�I%�qV���&=���D�0O4�p���M'~��C������5m�'�@����y�W���?�~��J�)��z�҈!�W��o��_f�y��pf;N�������P������������זN(�n��ĺ;K&���MK<�O68a��T�S����i�n�6�w�l˙�wwm]r��[QBnp�g�9�Co�l�<�y��1���T�m����mC���x�ۯn��j��g����e�SB PK   t~�X�z��kW S� /   images/65d233e5-7445-4b75-a6a5-2d8c2ad1af28.pngl\	8������)�6S�BDe�ci!{�K��c��j�1C��%{IY���14�>���,������:��L����r?�s?�7s]�Tݹ��v�v�]Rց����u�V��֭ߦ��6�ϫ�m�϶�X��9]��� �
��J=]��׋W]u�\1�]nAF���my�閘��uܘ�A:�)�������~�M6%1hSq�}��z�����H8{�YK�3�;gWF��~�J��L�<<b���FĶ�7����=�90�kD'��޺	�󗾝�|���o�{>��|*�H�3���F�)�> �l������v���9o�����ퟭ�՘ (a�S�@����(Y޼x_�fϚ���h��Y�C��5"0CB\5�[6FGn�`�z'�!���)����!���P&��{=9�Ȅ��p�c֟���|b���Q���2Z���&�쵭c��\.�Z&E�vx%ڳi�V��&�ua�d�x4�p���x���V�$�T2�8���`�I������O;`c��2큈�Hp��G:��m/�s�D��1��ڔ]�Y��&(ƌ2ܔ�"ʿ� _s����g��+�r����[}l����ۮ|{�`���}SsN��Y��^o��ꭖ��[�T�O܊
e�ڽl|��Cm	�	!��t;Vf �Lu�η��1Y?���R�>V��D�1AӬ�LPr��@M�77_!~3�;Ś�㦚��Sm���p䛐~�s�ř���Ե��4�uP��H�/2���˅���L��RC����	CT�ڭ�}�/V���H+ɍ	�Z����Y��q�o�X�%p��-�=Q~�1R�J �y�,	A�	w��o9`��~��,�k7�j?�2�����7��߼�x Y��&�1�j+�Dӟ���%�e{�%؍��_h���3�~�����h�f߂[e��ţ᠝с}|@�ȱ�!�������H���h���aMi8��'͜X��]5�<�ܔ�JUÆ�f�a��//<l�Gb>�P왺�}��W����M�X��9����^O��)�0N���E��a�X��jճ���t�,��q9����� }��"VW�8�ɖ��wn��"�}n�(O�F�	��掤P^��~�Ee�XTu�3��Z�z�s``���u��)Q�\�����"�ڝ�C/qS2=�F���SyZP���
G,YYȳɺ ]�c��lW�k�m�0�q(��B�!���u��R06��K����ГP�l�������w9x��1���1�6)買�ʧ�a�B��v�[83VB[�_�D
��d�z��	�;m`1fWB0ְ�Zޚ|��[�G:�`�L�4�� �/ԍOr�+�4a��l�$� �VvD�V.٩�(8��NX�q�r[F�W𣣣�1:�[a$Bh�vm��wZ^���dاo��˚̌хh���߷oI�l� ��_��*וv.�yqn��Z���7'$_���We��ٿԕ"����c���n�L���{Q�N�sPhg�����ъ���7*Gw��N#���]����w �^��_��|<�a�>!�#���Ѭ��-ܙ&���p��gL�n$�O��tN/c��C6�f �u �,h!�"��c�6ha����V]��-����WK���=1�-T���mE|��֌����v��Љ��Uv݈�؅�.�� �Y���0�r˺��l����@&oIcti1Y��b	!��.qGc-�_3�h5{%��k��3�ru�ϣ/���n'_�7t������7:N�ڭ�[ 	9��(!8V;����Q26�;) �J�7JF��%�6�@��{IFzVق�� z#H*#�*U���3@�1{����Lf��C�%��V�@����	s�}^�C�,`�gřZ�d~/{��S!a�6aq��L�A�=zF�
���r9&o`�� �ֱ���� k��{Y�v��(��9V�7 �"�Eא���u�?�d�m�!c���U���7�Q_����x�p���?����Q�[ܱ5���7,Q"<��+�p癁;O\��[����2A���U!���n����5�bת�B����s޺(2�oK,��T��b�����s^���� ��d���fH��U����8�ZÃY�����W����V\�����U�&�Z�_�����5�=hE.�����N;��TC����;�=�? ̲cs9r�6
-;�J�3dHN�;S���_�������3h8���e
v��%B�HtCV9ޛW�k��ǰY#�%�
�w�6����Yiw�<O\����t����M�ν�7��+P���h����[�1D&��t&�{�A��f�4�+�16�O���tQZ�K+O�ii7[�#�d�3��Oe�f�oT� ��.V	�%��Uh'����=Wq�f�Ww�."
[8&.ʒ9����[�KtQ;8��-O���h�ٞ������-�X�z=�{�d�z,N�$��6�@q��r��R�ws�?�Y��0_)B`­$�8����}�o�no!��1�j���3GG�����s����(���9�/�6ǜA��9��5� g	ģ<�\v�By�:��,Kf���/OKcg��$�9yӴ�cNě���;�7"K��Ey��	���h��H胈Z����n]�����G5|��#�m�-�uQ���O�ޗP�p�UY߅釨�
�=�t�#޽�^��*B�j�-�7��!�R���R��to�\��8�;La6&y��@@�@��*!�U��p�S9��%N ����	-�8/�i�Ä���9�������Y^��	�V�.4g��E�\�0m.��X�W���w�=2����>�_���N ��(
A��RUϑ���	56vw�|��%�a�B,-?Q�'-��DD3�*�G��!�{M�g��g��Y� ��k���x����!N��#�*�1SZ_�ZM__[_��
�5>��M���`1y]T����O�Bz��?d]Kz����"=A/�rL�q8�?��uBǞ�G��,�*�̴�;v�{��bf�U+� c]�N�+p$-Ge���h񹀢d� �h
��]���&�B�(J-n�ĥ���"+.O����a�g��}��Ytt�!�h�s���3�\[!x3&�����&�<[�\�T����{���)N<�����uK��"E��̵�<��$�y��I�w �yԀ���f�z">�yJ'&R;�ptmf����*�:��c#�d�H�8mb�~~ϵV�*������=�666�(~6Pa7�������p(�����h�.�zJ�u����6��D�#�����/��S��8u:$���S�W��wq8ʢ��d=�{���5?����@�3�3����"D�Z׆��<��N(�^üu#��7��u�0�愸�9I��G��Y�+;�G~
7�"5�#{]G����y��+�xBuHJ�A/���J����!�	���"���������޻�7��.�͗�]��9Z�#��a��a�����O2.V�_���� �V�%�H���ח�ii#]�H�N��@����6_	~����y��_TQJ�������9������l�`�3:;����(5�mϟ
keF��
~x`G]]]�jUnjT���J����0�*-}}��T��rWVD��G{�����
,.YZ"���s���y�����S���C�cMX~�ݐ���+�᦯O���)peO!s�,�+��^��$��߶��	�;Ԧ��'|f�Br&����s}5�5��{���-,�����wT�
mVxz��͑p��N�f�8Mc�����"�70(��F��sJ"O,�$ڛ��2!hEl����z0�F���.e� o"��ҧ%%�i�r�3�W"/�a�{Ԣ)�ę����~A&r 쫗ݤ8�������˺2�-Mx�.;��������#&�j�Oo](�M���ɽ&����Sf�s�?䈷�;����W0���=�zy8��
hH���=����
�"�P����x���3ř!Lۥ�Mg�n�5�a���XG�@|rbFA=Trf��Q�+�D"<"n�����5��+�srHh��490H�*-0�HYn�}w4֕�ڧ�������f���Q!'�Y	��9B^��0[<�����m�]�%��%/��U�WxY�bǉ̜��lO��~1��;��h)/�`;L��M�s��hfV,���`���e�����Ak�o�	7Ŏ���c&�
���/&#M� ���"ZvE��L��!��?e��n�t\�<q�8�ۜ�ci�e��vFx��|��1�ʡ�}S.@0�(�<`��b��6+$�;�s�6��Pk��jQ:���e��61��dW���4S�t��f�`%fL|ˏʇ�f�3�ɑ�='E5Z�M۷R!����e`�UՒ��H!�N������uۀ����N��x�� ��U��@y�]xƊ�uk����~�1((��;�5�[#�YF���Ў�|�����������;���и���R����sӌ�׶$'&b�p�8�zJ�҆]���JKkV���3��N��/�4��~t@=X�3�c�xyP�+�bk�X�ױ(w(>��x��_,��q����ZU�;T�D'��,�[ǔ��:��R.<�6F��C�3`��L���C�����z|7�I��s�ʷ_����Q�B_g���u�"vI�ǆ����ol�(�?܋�'쥺{�T���|y.�(�s^v��g�:��A�,����b��h�Dw(��?���C��L�y1� }�@/��S|?ĺO����i��'����C(�IZ�M�W*��Ͳ��mP�+g�^S8-M��m�"�/�G͒v��!�u��*��Q�����$��i;t1g�y	��g����0�0x�E�y�\�"���(�}��6�J��vnE��: 雰�y�u�ף�בPpğm2*R��5���&i2Sc�+�Q%����y�Em`��r�YS��qX���Է�
d9� �?����(++�W-eT����x�� XZZ��EFr�:��BLb/<d[jMKŖ���*,�8���)"��WF��c�a)�8;$S>oB������A��:K�P⭟�C+,v����Hr��%�B:nP���Yx̠k���+S��Oz,?{��l?F��0���FKUg��77Y2��? �ܪ����;�T���Tai݀���� �������zIϲ0�>���g��\��,��_Tg�L<c�g$	H{�ª=@��Z7���we5�&�>561񹈢db���O4
��������K�؈T>4�:--��M��N����VP�^Ɣ]b��e׉_ ��ř�d���a����a~�`�?�~�8a/�"HX��p<�a�%��Be�� X�Z��~�562Z���b�>4�HȰ�M1�c	�����m��^��p��U�'����3%�\c�"B�m{�$��vԘgqq&��r�8~���UNs>�?e0Ն�rs`����?ղdwo�����N�\�T^�j>�e�������~��=�����/��uD�ꯂ�n#�����zOds �� �X,mTD����Dl��2Lj�Dj��T��iY�x���l���E���~��E_��̑T�dt횧#�7��c��x0�����Sü�Y���N%��b�ʣ⷏f�du\��1x<O�Koe��$��_����6?�����eW.Ã�3,��dd\\��?�MH%�Iu����>-敔��t�6�|�'Ӏ)���,vqL$��w6Kʒ�錦љW�� ���)��g)D]`r��"~��[���^⤡�|�'α���|%/˗��GbĢ��=+|�aܿZBO�}��zU��_����eR;�7�c��J|�����/_.�C�f�p`<$\�?����2bθm�ߕ�e��YH`��m�bq�O}lsE_�5�E��cBX�0ؒ��b@���
\%))8���ZJ ��ڃffܲ�%��F�\[' ��[=	]~�C�n|=*���8-5d�-�ie�|�'~�gwP��3�N$flњc�A�*A�j�n��{�O����Ihhx�[�!�������̒�� #yfa�z��K���t5�0��UNY��(T}�1Xm3�RR{D��eWg���T.c�o�n�t
:P� Q��5`:�O�>�A��yj �sDjY���ga�B= B�\?99Y@Ƒ�9JԻI��^�W���p�G�!�?��q��F�G��T+ ��4QЮ³O�`h�J�׮�gٔ��-s���~��@^ǣ��  �=B&K@����m.�e��^��Vr��d���e�̒�οbNn㲰�����Q"�𥳐�LkFF�8������r��Hl�����p<��M:L-��U��������\i�B^�f��J����7����ŵ�������7m'����N�*�1�;��nO�@�&}E��Zt�?K�u��ϧZ�^�F�ߴ�Y�z�e�x�Y���K�4�#'�޶�)�3L}��.v���,i]9f��ȴ]��MO?�)��Q����U@+�z�F�]8��f:�U33������C��Vp�'Nf�����" ��+�4 ��Ox�mX pÓT��gr�R�j�(d74���`;����䕒h�ߢ 	�?�9��9
<K��<E�y�Tb��l/��.B����Ɉ��4�^"X���#�i����Ȱ��"�Յף&O �j,$�♠8�0�����P*�e̶�x�JKC޻�(d?F�4Ѝ�<��fmڞ��f�jeΟV&���$$�>����q� �����@y�ׂEw(4��^������<����I���4��th�[�ŧnU�r����v�rl�Cv�}�Q9/���c��5�vq�AYrH�lzZ�W{E �c������-�z��X������*���b��Ye�G�D]��}~
��t��c��4Sr��:���h@����ZE\:y\L�OE��q�fw�����Y�R����bzT�vr�/<�<:�/�7��
� @�:=R�i�	�D'0�b�+�
�S*!],`d�*}=��͐��w'�ș�׮�>h�b�E >9 4R�(�N=0Z��}���z��y=�+���zZ;��6S�����C2gff�g��Ѽ3��D�*��U%�ޒ�=�A������	�_�a�"O�_�R�C��r�!��O�$��� 
����,,D6�prt�xj5���ȣm��:��z$����ֹ�O���Q��L����G�bۻ� q��Ro�[���߆Wf

*�ӟ�P6Q��=R�ڪ_��D�R���2�G�6��Fu� ����;�DibMC��(��3.+�ҩ]t�cǎ�+}�{��}>�9�lw`P��3�d�϶�ň�[�~���{�h��a<'��u�]����Y+�T���0��Gq�	���xeX����ҵ�'N��\���T�Td���n����BP�i$����Y�ӵ�q����y8�g � U��"�ٶ���?{�%��A���鍖666��~b�3Q� ��Mf&HWb�&h�fʞv3o��rԶu�$�亮Bd���%=����q�1f�����}�EJ��t���¹Ǒ͗j�`CC�|�1(@+=Mt�bm���_)!> e`�v�m��7~����u��ŪIC�A��Jv�E%�Z�[�3�`�o����!���
0�}4d�����=(a�٢S��SFI��S��^�Dt&�f�&BHyo�N�$ߔ:��;88X��Q���0d��(�D9^h���;������x~~�c�VX � !��pt�A�>��ISjZZ	h��C���u��:,��$�a���D:�I�SE�&&���2_o�����q	̫W��4�'0���ȧ�SGȠ�xa�n��ׁB�*��.� .�Ru�e���4������G�uhoT�E���c"$q�+{Ko���(�4w떸�K��I��x���	L/�>PQ};���Cl�J���w����pW\h
�~��x�/Ի��@���,�U�顴�(IG�8�(կ������g�^���
zh!t�Jz�����`Hw0�6�����A�%& \,���8�H��h��L^���iL�]�.<�Vv����ż�<�>�gBs�@O�د'd	l� �3Y0�����u�J؈���L�-=����E��.j����Z��ǣ��&]�Y?���̍���������"e��n@P*�A��a+�@��g��g��
�Wxg8��;��9~66F7g`{G������y|F���b�@��ü�}�hT]�<�%�q�܊C�c[���!��x=�۹�W�>;l+_�o�u�Aj�����{`�9�T��z�XO	}�[��k���쎎�6�á��qa�b+6�bz ����l�.�}����E���x��e�?G��?^��W?X����>ZE�bOT�d�^55�MI�m�����v�&��5��j�b;�������0��0z��i�O���
�����>g�}���,l���!&}%�泇3���z�7z�����>Pw��o!�T�l���*?��cϴP��� ���*�J8���D>֣I�����x
B����N۬�]���X��[=Wq���>�[�h_�2�+�z�H��>p����@;�?�/|>,���;��4���H�|;����X�VVɿ�;9�I(z8٢���M4v߇˜�=-���s��}e�k�a����-�2�Ehkߙ��y>UTTs��	J ��������MoRb�b��܏�$�/jj��V�ɡ$�E
N���<��K^;�����T	{�"�P�M_�GEE���^�G�!���1KMd)�����
]i��6�IW'�����Yp�d�����'hA�h4������8y�L�|=�,�B�G®�c���b���ހ;t�u��Ç{/C��F\�r��c05�1�&+�}�SQds* �q֩����t���oEig.�F�}�P��j�:-�8�]�j} ��S__�q�y�k��\�����3�]Kz4���cZ�������E���� �D���+�59��_�9�,�_�`g`�A�^�4�q��>DL�]F��\8�R���	O�o&f���m���I�f@��2�����a�����0740�=�v���[�f���	!�����s|4H�{���y��:�q���)N�d?P�|�)77L�RoA+��π���\E����z�F3rE+2� =���xv�8�k�{gA���/jK�ƭ5M�ڥ�>��?])����� �Rp�p�:��$���q
�G?�xX�覶������]�����<��#�{ە��w����U�}Pw�cţ��N/Y��F<X�v�������:*g�і���G40�zz Fe۔���4b��\5{L�VQ��4(�N__��� 	$��u��C�/'�n��ID&_Fە^�*��"3����;�y�����CJU���n����P5�_x={N� ���.$7��9n�Z!j�����܄���Hf:���b�]d�Հ��e�G����μc�̵Q��K��`���Y�K�������0���'��n�	]��M�M��ˑ̐�sX��Am�4.K!%F��18"���<�,�عj)�E���13�`̆b�؝��b%X$%@HJܩ�9%Z{KݎTV
X�2!�ݓ�\��B��c�[�[�Ѹ;}���X�f� L��Iu[�5�y��NM(O��h\�Q@��uLQ���
P�?�欄��/#:�K�X�}�Bq�r*�&�N��Fχ�?vw�X.2�x�lx0���_{���ԝ���o`1�O�+fʿ�#�k����!��%��y�f\�r���y��\%_�ڐ�k! �c
C�n���������i(y>Y�?�� P@IIl�,:8��i�FR�C͇�މ��n	x�fa0o�®��3��L��fD`����!�J"���b�%�F�;I������[��r/�9�<����Cӊ_���I�^�Lm�h�7��qn֭�,>�[�E�'Y�V�P�>�?����e	��Vd�����q�	���B4N�wA�A�);���o@-����B7��h�E6P/@��;�s��q���*�/y@x���t�rb�Ū�̟�@Á���E~P��x��M���s+�K�$j'��	$Y��Oo>w�f��?�q�omm��9Ùw^x�y��f;�s<W,x}�j#(�������P{��������K9q�y~o�:kIS׎2~C^���e^~������8�}��%����sU����Y��XW���nzy���/iG!(� ����?_�T������CqV---��3˯��ݼ�U_Z�~�ԃ���x4)e��$��t{8\�7݀���z��F|�U��t�c��O�ə�g5���J;�)�Z~�(�{�*���B��e�F�a�rZoKﭙ�ds֗�/ϘRw���~�>��6s�5�5J\�u�d	2TL���}}��5Ȟ:����VW�8���ɼ�1-?�.�g~P�޶�K�.�
_//92�q���!�,+��NP|��iW�/�2���pnj�Ƞ�,I^�A��N�5%DrʧO���?���7w��SW�����GԚ+����h���Y���^{��e��pb-��Nc\�)V'�̊j��*���;���NAX*��t�/�[=%8 �;��MK�쬍��g������M��N�y�8uܵ;��'�J�;�-~��0�_�e�}��<o<�UDa����70:��>"EБs�X�,C%�}A	�M�v+�͗�I�(���Y�Y��T��A>�=`�:��0�����+>IG䀥^V��*dq����YF᎕E���BJ�4A|�B��3�]6M��`-�<�j��x��=t!0̽�Q�!����$?�a�f��T�Nj���v%$��M-�VVw���D�Su��W�g�/�@Pcrr���
��"����}ư�6�1Z��&i��S�̄�='���~�5v5��HkMá}/+:�����_�q��bRۭ0���m!tD�*�w��{�V/3�êJ^�YRy�&g�"~�nj<�]GRҵX b��Ǒ�V`|�G~u�?��s���2�{^��y����5��i���U�ʳ+�m�@��f�Q'NW,U=�ӎ*N�c��2�0H����zuTG,z���!�"BP;�hf�Ң4S�joo�%�͵;.u�Y�y��LPivLr`���W�G���37&7]�ڵufl���Sa���$�_�Jd�Ȍ���>D�ĒK�[�h��V���v�Μ�-���17r7��;�ſ�?πa���E�,=��^�N��1.1s���S�g֬+�@�����S�:�5w�z~-|���_�+m�ś�(����<��%�-��d��S1Nlz��X¡˽*w��]�e�[b��� ���|���-K /�>c����8/��1����^^�5���M�~�t)��X_�D�����i�ׂjz��g�7s�tR51��Wñ�3;N���Ü�'w� I,���˫UW-o陭r^�-�[���X꟞�B���5�3ҏ�E��~ﯱȐ���*�ݢ�^k�u(|���E�VX����8c��iz�~y&�B�'�(�/}�L�)!>�L4t ��炒�<0��^�7|��mx+X��'�����cE�
Ki{��5K����r�l�����ռ����d,�Mk�����F��R���=&�5��̝n�>#���_B��B|����j.���"��Nȫ�ݚ��Ԭ=ݕ>�rGAlA1��Cj!*�4�k�2df��}��ǘ�>RZ��7��*����	�j��1�����T�-t1�V5ﮞ��r��>r�[��&��m
@����=�"0d� ��jg�����¡��Gy����S�2$U5�lo�����Tҝ�HA5�W�}�"�������t1��qݥO�S��ӮG)�TN7��/7��10�`����l����իJ�gz*��<)�]�o��ȼ�v�����m[p�m�w67�W-=��o�����?��ѴC��ƿL�B�s(���8`^��M����%���A�/��@4Ro=��ߝ�g�����M����^!��;y73콽m�\��
��8+]k�/�}X���ۉb��G�m��e@*gF��x��E$DEޱ�:%����Ö��?�
�,K`��a���:��Lj��{���MW��p��fs�&�Q�m<��3-.��/-h�z��K�ݭ���s�RK�+�����С���.>}��Z�	
W��$��c��P)-�����'��>˒��[G2��AlCm�;���g����2���U�a��B� �*y��M�{�.~��I�i$03��;�?�����Mp�����p%�L�ys��V�#K�a����� ��(5��~	�.��0�-���P��RO�����A�S�,ph%R�{��G8�6��r�A�~��h��vm`sb  U� �q^4j�g=���vϮ߀E!���Lu�Sգ��iY��SA�����ˎ@� 9.�o�d$�	t]~����]@�m����ʯ�n�5^wP-��2E}����S���c]��W ������0p�"�ĉ��ލ���/uL� �,��C�]+�'oԼ�Ez�:�ʢQ�wJ����]W�,ǡ�ns*X���Z��]�vIX k\�NMh�z7�%J5�|��Ӑ%�O�M,.���� ٟ�߃p�����,4����p~�F*^>��^C�P��ϔi5?��G�����@v�ךK#�NU㞺j6˒�-�cj�h���*�ߞZ^��3^*(�1�2Y�ZY0޵��Gk=�扈?.�ݺ"1�x�?�RT���sUO?6����@v���;�~��ʚ���/��֭�!*��5�r{:ְH��Vc��P,9�dK5"��X?
<��?I������ޡO���?�b��N�CC�RDf��e�����@�������\��Rw"�}J��YK��	��\��*f��KŪ���e{7W��[M�NMM��Th+�4-d_��!��>}�ܝ+�`�\��	t��.�(c����X$
_�{��i�ڮD>� �P� W��e�<.��eٝ�R����wD7�3�7�;�'(Bf~��}�gl�u�iA
�\��v@jyF��b��#��y��=�Z�3�j�w�@M�2ҒJ�%�L��?p���=�v%�h�x4����܌<%AJ����}N�O�俻]�2n��	@T<3A�_vb٪�ksg	&k����?p-���")�9��؂��"w�P�R��i	�M>���܇�f�Y:�i�s��A�S��V�u5Ev��^'�ǘ�(�]�5UP�A�x�4JV�x�P�l��}w�[�Ơ�����G-)ZJ?�_5�e]w5jF������0;�ڇ��1�+�z�a������W���D�=������۷��^'��㡖��je�[t�XT�'�ɒQ@�ڝV�RRR�Vw���+�m�u�<�Z�LU$2�t�$����͍����k��Z�V��u9p���-Ч���Js=�����PV�yaV<woP��qepnb�9r�y��
�hq��/��;�g��D�S[��>b~Q��uzX�eG��w�c����ǀ�Ů����GHZ�y���w��/�J��h����c��Zӆ"N.�P$9�ҍ���֩z�y��uF����^�D�M�s0���7����z;�[��E�H���;y�'0=n���e�N�;I��s�XkD	��Pf�6����zc�_�>Lq�5x�]���l��)�5�%���Ji�A6_�^T��X~e"�_�A�ð讪�Ҷ��Kzq5�Ѹz��}�wCG /��Roݐ+,_��]��H%QQ���"�%z�7�82�`�N����J��YNKII�t<�Y�������O��e�*�:�俲��)d<�m����!]x��� -S�s���9!Xr%Lr(�F'�y��r+���������Hϡ�{����^:�Wc�4��!\3�r��K�}�Fz��Pg��$����ч��ʆ�_�̝�J��˹��3a�[�C�;�-HEU1!���49y���{x�E��u*&��BP-R��(��O�J��KccM�δ�߿_T��he��?�>'jK�9�:^i�~&�@A�v�/!)t�����ۈ���F�!&5C�<��.�d\�l�,�K)%U��(�#��3MOtƈ�]5��Cf��1���g�¥�B�]a��˘>6�g���BSw ��W���>���5��a5{�x�f����D�//9��W��:e.�%�y�wTf���+�������_7ȳtAι�*�R,�NܙP��V9���b#��7;��q�M
�����)f�Q�ˈ�E��ϼ:�"���5��Q�rb�'>�K�4V���hm�X1�x���hy�m��AK? ���w�=�m���&k5����K��B���(�Se�Y~���S ���E���bQ�V.���*�"��Q˝����E�H�����O�O������u���]	�{,���._���I������f��E�Sd���6_���!��?!���)�q�%�o���e2)�J��-r�K��B~�����Gi�C�y��z�<V��
^��I�K^/iǉ�]�p	�.�xh�n;$������K����|��_G_�1��^�"�'-�v��3EQ0�v�!�|ya�:� 啘��&Vi����b:�@�_���[=y�G[t&�e��N�}ɢ�]-X[B&��f�u��K3⧫�_hF�Z3U�jn���ǯ49#���G�W�|�+4�R �B}�잵ʬk&����B������Hr��k=Q���1��W��Ay��E�����/ ��rg

�c,�3mZy���5�f�;�[LK�L�.�H�M��U.���B~�d?`i&BQ$yBﲮ_M����@&٣:@V�]��7r>m�!�6"�>�-^��b�����F+����T��d��N}3{#��۠23�,9�������S�xB�s��.��0��5�e�}�3�D}-n�,	�t|��'rW@Ơ�,|p��7�@B��Y��}�w���u�����$m�.S���̭T
�9��~���=O'U�gs��B�ZV�Q���A�k#�A5��;q��3U�ġǬ�nv�1�3�
���Q�{j&Z��~�����σ.�4��j�QT���-�6`�
����N�Oa���������}'�T6>��S#����!"c���\Y���: k���8�I�i	��Cɡ����W|�jز�Z� ��F��ދ��m����?�N1C�?�Uy�K�H.q�~JL�	0vN����k��.?�rQ�݀Z�7Uw^��*�����4ӮT���0�"w|�1��W��4�Q�<�^cc{�$ɿ�5�c��R��!��q�I�¶{)�^a�*>�ⷜ;[�e[�2KB�D�86��bY�,QI����r�9�<A�3�D�\�Y]���d���r�"i��ܞ����P���ѽ���~t���000����8`�l����s<�t���X_~�9� ��,��Sշ]\\��'!�v�m	$?7E@��,�O��'..6ׯ�ksP�<�k쬹Ob�)y��9G�	�~�[Η�"]�wX!�`.�q�z&�+�gvto蝧.%U���wz�K���Mz�z˝�)n5�1��P��Aw謖��S�1��.(`!!���\�|O��>Sm���stR#%��E�',oa}m_<X��jh�=�$1�a5��{���C�����5U7x��~wC�Cx�c�$6���~���l����>���[H��9G)3 �Q�.�Ĵa�^,���#� sz�]��9k�"�KVa�4�'��J�ti��GE���<��a�X�\�
�H��ĈK��w� &�@P���ͬ{�\��l;�-��.~��QhA�R_߃��1"Y.��؃�yjvy�M`����---Z�-��2,�!�˪)i�Ek1�6���lN�Ѥ���K��Td2���By��㫇ʀ5�V���!L�Uy��2899��IcvdLBN�e���( |�,�2̵�í�#��RԻF����zw҃�p�C�|�Ty;�O�8�T&���� �H�1���<�pjBԴ��aYɦ����`���J�K�و�G���[�w�E��RA[� ���ـ��:F1����s���{��s��Ӣ��w���sSw����0��cv����l(����oAl9���������s��h���,�?(�E$���B�7�m�R��W���!����C�T��vөCۊ�
�쵝���>��E�)9�U��Q��7I�G|�c�[Ā�Z��:e!����-5���k�c yA����:m��E:'��PBͿSd�,�f��2[��[��+c��ǵE�t���|�,���]��<p�]��`�j�,4%�6U�U�]=���zA<q3c�����$zt � �=5u�m>1�Y�ŢIB��#���\ș��Hc���բ!c��=0n7�����yY?Uo�ܗ�©pi��1E'�S}A
����F��I&hᆧ�w�4y�N��?� ��@L�<	��b��k*�D2b@�@��K�v�K~5ʨϪ�n+�ȭ)-t��I�
Q.F�?��ԁ�'��S��{�����{8Ĺ6�5�u=�/�eŞI�~p���NV,?�!�*����(��*�@Z���o�=���5~��_M�a@o�O�l�P�/%s�����&1|�9�z���Ʀ����u��v�"�� �u��d#��u��uD���%�^&�X:��O�bǜ��+.��i}�L.�P��\1���`?@�J��!$��k��YI�2�y￠���/7~`Qzh���l��-4�|�O��L�
��8�m� 9�rbפ�?�h�0��4����P�*G)Q��A&[���l���A����G�8���K6^�OwAe�b���'�^a���5�	��Α�`|<��R�e\c�Kwww4y_&� �+�X�sI�}s\���R㷽�33Y�ܽӺ7�8� �m��M�{�<�W�C��q[�ӏ{ �r���o'�?(6&f��!X����Y��.�sC�f ��k�#	��Ho���z��q��H��4avg�N�5������7�BO'�F�?2S��ߖ'���<u��� ���%���2��+�ٟ�r�bD������J�Dd��B>Y����։!��l � ������'2�cVF�,}-`"�=����F�[�O$�%6~|E|v���%g i����@��x�j hh�L7EӴɺ�?455��9�v��/o�}N�Sk��^Ώٱ�������	����RX�U���3Q���Ca�ӹ]�Ļ�>�؜���C��"@y �a~˛�����/ ��i�/�h�,6�>V�S�Ա	��3�ѥȧ�-8�����u�͈�������«{���T��scC0�y���jQ��+K������I���6x��Q?.c�wsž��e��B�� �Ţ��1l�)]%�����'�[:vj��U��c�:���չ������y���D�{��x�	:��zbќ>,@��������%�]��y$̼oC���Q�@s���{�D,GJ��_ю�UZ{������7o��y��ߧ��@�E�n�/���y�~����Q��d<���}��&ngiɫ?���HW�[&2ob��-8/A�FC	9X2k?)��>�����1�x46��������s�/�p�����'� R�m$����/$I�Ѱ�N�	���M|qR�_-'�u2�L%������/�1 �\_�s ������9�\]TTQ�iii���!$$iiP�c萖)%AZZ����v@��n���|���Yo��{��g����qG�G���L�A��������h����������U��Ȗ�C[�~�����Lw	i�i>O9<6Pw��qh�@q�{�ݸ���}#@��3�5��;`x���,,xy"�̿h�`��ź�M�����Z�1 ��W=�����PǺ�<�9"�6F�9]�f���a&
a�o^6�l�&�f����<�8���oj�ނ�y�T=�I�U@�^,����_�)p��PB���]rSC u�G��o�k��Q���/8,-<���e��kN��9ͥ�߆������		,���ee�'�o�Q�DbO�K�N�8U�"�(x'��%	,�y(��	�k����`��A��V��cj�)E���(ތ�t�E�l�z�������ټv-ۄ�)J^t� C�Ϲ6�����x�G���
��2,=G`S�8��#x^��N���i3X�Р�30<c(��r�_�o�ʠs�i�S�-�r?�*h���s���B<�s��گ�fi�֫œ��-{�(�	�r�4@�e#@���:�D���q7�e��9�{�Ü?ȅ�$h��M#��Yl��\��|�����uY����`���7�R<֚������e�cp�΋�ПEL� Ӯ�]���!�/<�%����޼�3���	Qo7�8���`����/��H"@<_w������8��cr�0�<��k���i�y������V�<LqV�����i�O��O��UP����lf���D����F긲��Y^_]�������G���Q%w���ݪT=�3�����j�s��d�?��;P���0��o �pD�KK��(�nRRR����ro�����sj��f�e����y0`�4�V-�c�θ�s�`6[r�s�~U�\�S0Lc�t���M�I���`�V:���$�yG$�-؎��J]����y%��ߏ?�Cޔ�������z�O���|����ޖ$u��Sh�߬���[���=��i�[C̆R!G]�u�5�來��uh��9����߶�i�8%D>���P�~K���r�����u|�~�f�:�e���˵�)��F�32Z�@�����'�1�&��EDDd- kn��3!?��1����:�\��_$�IWfb0�I#e�%��E��cIW�N�!xX� h?���/|����؇Q���d�������5b�R?N�rѧ3���={�+++fs��"�Si.���(:$�qG[����;f�s�� \�ZG�h�앞h�m+Y�A�U�$(����j�w�����Jv��_�@0q��@�����{e澏E��੏ߥA�a銅�e #��c�D"<����7i��,�Q��#0��x�\���ô����C#��,�tu������`S(�X\�(��S@��t
�owt�Y��7+Z8��x+ ��:s:!��ju|ŋ�]���. ] �6a��Ŭ�w�k�<���!~7o��r����3<��O��>J j����\HS�R �&��è��]2e�z>���hF���� -p�*Y�hc+ ��P2V\u��̜C��s��" ;U��lRB�����ّ�0�{���E���;�������������#�7)@�6���M����yͧ��/��};�N=��`:�I�
?8�G���3Z>qU�C�j�x�$�e����D�@�>���#����9�}�,���u-�/DA��k��Z��2/�r�[�b��`�Pfg�-��3�������e,���|�ja�����+�v�H�� 4��Z, ��[�s"����_�>6�ڢ��6�:圣�в'��=���T��v~~WN�_��\H0�
S��M;]����ͷ�`kە�ƧMIM=�-IШ����r�9�fd̑.�{F�Ps����O�ʂ6X�R�c1-���8���d+�OTU$�����;�W�q��y�(Εo�Vˆ�ّ�����J��>!��As��l�������� ���'a�5�9��'�qL_J�a<�$XE�+񱀠�ua��/�����V�sͭAQy0�\v�ӑ��._��liGM׌=�M{�7��8������\z^�� ���@c��hn�6�a��ܯ?ò1]/k���Cw�Z3��Fi_��x��x� #���/�P(��t9�� N� N#~rw)@�
m`]�8��׮�`��А(>rF@����������!��6j3�/?����f6Ld���@�&3�����fYIc�CL���2��
�	(�U8>��-7�����=��J3��k1�l�eE��2�!m�$��:m���.Q�����K>4�D�>�|�NƏ�E�x	=[G��l r�͠���g��to�@�5���|V¥���YE��V����J%s2�%ș0�����b�6d��=_����"|L�|ߘ�B"�N���<���g
�?6�����1�����7o��?۪�4۷!�a�ͦMs� �md�M��;����a�m�	�ww?�5��Z�7U��q?�Ā9/�$��9�5���_]+����+�.*�־n8���&G��[I{I��0D�̓�@Pz�k����]k4�	�~w�ԯ�W��>E�Y��?��y�����g�̠p��`����AN�|KS�fL+3���ȐE��ŪT�f�^��3���M�ZػE!�t�%'"�r���	P!Q�+iѡ��������kP��b�
:7�K�<�r�Wk}�x�"�>Ǜ!�$ }	�cB����e�Aˌ
Y<8���mԾ��gQ �e���@Ҭ��|��!��汽�6��`1�ʢ���c����tO�C_eY_ ���/���UZ���v�r� ��od����!�,BZ�w��_�4Bi]{a�QI����l����V��Ӓ:Ɇ���;[�,B1!8B1�@��
L&i�V�5�~yq�]?��Q�i|� �*�5W�5W�d�=���닧�?6�	�s����-�z��:�Am����>�S��(m�$?`�H�����b4�� ��R�e�@�y.!|O�fLP+�U�^��5?���t����:�	�%�Ķ��א9_�9߫�^3�A	j��+ε���(B���dU ��Gz�	��6[�">����0����Q���5Y+��Ţ�4��,l<En��<���,�2f].�Q:9��5�R�n�u�����GZV�#0M�E�+�(˿7��=�T���OU0΍��,�vu�	FPA� �pw���6��/.����ĩ� �����e/�
b$H�G��"��b��#�,Mܜ�}���:�����W����:��)��C���BB�H�Ж<�l���2�*��f=��.�@%��S}��}���o�Ɵ3�K ���6_7��2)d��e�W�2�	���?�H�9�۰r����o�r��8�(<�ZZZ H���l��Pv�j��l�c8Ŕ��:.L$r�{ �{���n�������Tb]U�Uԕp�dR��d��d8�������g�����X�5���l7G���Oۮ�^����bY�vr�9���#jdr ���0ό�'��vbds�]i��r�)`)�~��g�"��
�H�[�f��.�Ӷ�Ӷ� �j�l�}�C�k�7o[�ڜ������>��ZKꞩ��C\{��uA^��\��;��0N�ȣ���H�@Qx:�Y��!rc�M���b�朆s�bHz�A�C?TL�
y��.j����̊���)���s��f����s�@��8R'ͨJ���@H�� �{$6��Z�o��_�@��?z��Lu���ņ�:�kO�M�����KV<�'!)99�1�UW��\o譱�ɯ�.ɸ�	|�q���k.~*I0���K���,-��+y�\�O(��U���޷o�ހ9�6��%�.5�?��j $V��T�3�333�G�Qc��+�	~	nzA�����ypZ�pNs���d����y���P���"pؐtk�BCC��ۋE#��#��&&&v��"_K�MOp��A�OO�1x��y3��𓷮���u�x{���m@B	U������z/^䲭�	C2&�899�~��N܍�JLL,稡4���$�4;1'4-"��w|s�Di�}�V`����O%�m��_ǝ�JЦ;�s� �M/�"�ܓ��C�꣎�9���=ۿ�a��c��"��"�6�����t�$��h�L�9SGī�;�$F���)�ÎοA�������9c�1&���hS�o�P�>��"�5��*cO��G��B�'Y�<�B�=�j��sr-;c�K/�Rv��7�ɪ�d�ڏw:tj&�s�޽������m�����@�pr�X�� C|��x�C���A�ANs9F��J%�x+��f3�Nj�}Ԩ���1E�H8i�'���>�H��1-��y�$$����f�uϽ^�h��#���Pbq����y4���bc3�=�J�yxi�#�ڄ �i��6����zg�=�E��d�����W0�V<]��ASLz��~ERRqO��3=�r�J^�/էn+;�>�>1B]�o��#�f�b���#"n!�8�z	����hA�������gܓ��՝�Sl���7�9M79�uZǚi���X�S�7(�8�aȻ%ZEk�h���`�/���ʒ�$W��r�c8m�:�	y�r��=�.���}�G�T�+O�9���s�o��X������"�Ⳙ����+�ׄ�Łdb⑱������(B��fS̀���)���'�7�o������o�7��f���ntɕ�6�?<\���׎�~w��Ń� "D���i�zm��$b콘7�%��	��?!X���G��39q!=��9D�R��*��6�&���7��aT=2mԫzĲ��0*����s�J�� )�h�Ua�lz�bQ檅�1y��i�N�;�̔����U�.'�±l�*�&n'M�m�ZU�T�o�%��G��o��~�ج��߁r�g�O��Wh�����I��E�O�D����^|PKL<�n9�����jy�E}�Ӝ��Դ#6æ?	��8�����Z���܈��Ҩ�H�?EWg'����WH1�P�;���X�>��b���H�4}�xv�5�&y��o ��g�S0�C\(�9�zO{TP��р���")�sS'�rw|Í8Rv��Ɲ5�k+%WR����AG��j׵m��bK�~ttD��Z1����f(��e����q���[��*9�	�2	DjFo��8��	d|c�P0d���GY<���c�S;��\�,�j���GO��ku�娍��K��M@���	�#��ǚ���,�q��x��^j��i.�0�{Q�%=���V��J"k�����k�e���ݖ�p�2$Ff�ǝuՃ��Ez��=�;N]Ӎk�I8�$:�#Cj�b�0�T ,��l���𚯽���g9XM���Ǆ|���qky�xrZ���z
���SZI� �zpk�\6�����*���������3�MH�Y:���b��~�q �t�G
�g�sV��b�����bVE3:5��3��q��osoT ��?fSc%~R�����&��?y`�W��KY	��'���`��:�/�ih@�0dƒ*�q@�=��x���Ա�1��7g���C��4r�ȇ������r5x$�f�b��I.�*�qb;��h|�������NR�s�s]�{�%?��i�M4.L���>�][q���늌���u?���AoS�`�}��ڞ�Ƞ쵑�Ww.|p���o>k�80��p%KW��66Tg�����}! �z���_���d��5o0�fг��E��^@�����l簇4|)�G6��\��BZK����D����AxSȒ�n �;1���MT�c_欒��%�����B�Q�����X�V��;x �{�L��\�a��#(J���Yb%��@R�!�u�L�WjA>���.��$��<||�'u�+�����~	�(r2���T�lEV�n�k?;��C�&�����6u��לo
��\k��EG[Y���q���(?����9j!��#������0%f�~:�D��) �bo�>**d��G�
���t�fO�r5��h���q����_�5ߏ̅/�>��U>�4��
&03�y(s	���Ƹ���[��1=�O��^�_���yPݽ{7P% �F���u���ݛ���&����&
#=�L!=񌰬Ť�bsNV����&�>�K�Q�X���q�ˈ� �;o,>^l����%�jf	��F�}����-Z]�������Ӵ�^`�*��4Mo�.�m�uD�B�6����j+�X�*/C-'}�X_g�,�_n�� 1D�@0�Fyq�ؘ�g"��q��u| C(�?�ќa�o��X��1� ��q�tCL�U�����^�b!N��4��de�pV}��>I�(��fDq����7���ap�Av�zɤ0�E�T}ןfC�:b�½R�mI�\�3�A{o���N��wNfpÞ�|�K
&W1����ff�Mlإ�6=�K�|�����Њ��C)�襵���n`�bf�sc��0u��T[�j8C\/���aI�K�I7�Jݹ�B����[ElGw��g(Y�4K��K���h#��/]��/�5�z�z泙�Fnj�i�
�f��A������X��PX��8g/,?]�P�V�0l�xKCd��0y뛛K��ܷ%Tr�Oz.�)��t��Y��O�DOK}�է	)ٖ��b߮R� U� �5����)�=�AE�b0iB���`����	~��Z�G�j�F�ys��j�ʹ#�Ps�u%��]�n��e.����1i^m�25;�h��==�P���R�W_�f�"(���_@�X���O�ZK*,'Q��\t�[�wA�{��-�J��=K
1-7��[��U�83�X�����z\�}r�;Mg�äG�[&옷y�h$�.����NOV� Z�2d:h�z���u�����wX�r�v�j�{���
�IB���XVR�&�.��h�s���ޕ�a7�O�J��u�I
�b�zf���;^�]�zA���~��6Uz����v�vc���[C�=`z11�>>T2�{���lJ&�u������|w��#�a�l�g�q��,T�	L���p�><W%�	s\�]o��'Q�����eɺ��x�����$Z�ӝ��?�9@�>W�V�W�6��2iE��մ�����42<'�yy��������r��KN�
ƭ������z��^�L��.�"�ڵ��:���J	
'��d�S$�}��J	��s����!|�djk5�����T�ٝ� Ȭ�A��6'*��^H�;�̥�����1��܇L����3�qo��8>>	?����{S�"G5�������aītL/������*ʞ�V��@�r�.�@���mZ��ŝ�O��v��7ߓ��88�h`Eȴ'���R8&P������W�#+����.T7�M[E�0�DEp�����G��Y�N���v�"Za!�V���X����#��>$QBw*�av� �)��y�7��s��§��oWgˌ��eG��0���5��'��)��K���<�+��$�RL�H�؞gC�Ƌ�� �:8`� z`b2|�6�8����?4,
���p�ܳZ����|�r�.Y?4��9��;��T�~ػ��l�x�Wb�ԇ'�@��)�PCC5�Ǐi;8���PeՄ�^Z��TVWW_���L"jͨӴ<V�-�2��G����@�g�B\P�~���Ҙa��
l��Pt����y��$V���VzF0�I7joooА���og�Lh+�R�,�^󞪞�Q���J	��u�=@	"�����c//���Q_ᲜBv999c�P��c�����;��##���CM�Ӈ��_;A�,���:XlE�5biF�9&}&+�ǄhQ�]��	QdՌ���j;iE��S��F��[�˪Qtm��PS�%QS��VW�_IEEJ-!�%�B�~Z�]�Pjl���.�c#O��!����X��@���ЮP��8�[���l��(*|e��!\���1��'�>Pm`\VW-���\'�&���-�!���FN���\`�Pĺ*%Ov&�d��p���R$���۷�_��x�ܟӞ/�K��a��啕�5DH7՜_S{ڜY��}=���2�r�̯!�޳=�7{Q��j�l�V��-������l)�,A6�s��=��a0�V4.z:M�c�D 	������j��NJDD��XN�,�����M��\t�푑FA�DFLD�VP6�Uh��������;�h�>Ph|�y�����V3m+��nD�v���Ֆ��Z��ة��Ï��g5�[O��(���	b{>XQ@������yH���t�Aۧ�>��)4!�#_��x�EdA�Px�� �򲲀����X��ZIuM�=�Fޓ��6=�v�����mm����脑]�&s�a�N��<8( ����r���K��K%B��'�v�D3��˯�G.=<�<�p�[��a �g�^�U�s}�����ϯ_� ���/����������>��V����b�������[W�q�C���`��Ai-�(=?eݢyN�,ݖ�4�A��|<m��{����^"H�-=�V�>޲�t� �Ǆ�<������9�(}�#u?�a���)�a2�8�``KƳ�m����9������r';�}cb$��+�.%so����6��g�XX�����0U	榏}s�W�s]D#�aQv�W��{g˯Tn���c��efc&���!=��m kB��1 U�!�<�P�Q뼌U�_��C4��N���б���ۂ��o�o��k�P������4Y��%� ��,9��I�no��}���"�v*p�؉*��{�)��)]��S����ыB�:�P����G�*kj�uc�W5狐g���}L�'sz�XF�Q�@*1��i���{�.j����ۛ���������-�x��}d�y���M�\h��))�}7B�����U�i���x�E4��Ď�gn u�)c{x���6�`6����#���Ij�^q�;�١V�dySS�֖c�'����vI=VF�����qv~��W�2(��s��őZBs�Jkv_{?eQ�2f�=�g��f9�|����|�O��C:I��g2@� �\��>-'�ӢNQm���@?lⲴa$J�=�e�UG�S�$��N�ՠ (��"rPia~͉��$�iRSSuttZAx�s.0�l�?��%]�j����P��,/��,L�.;�>�x����Pe���[T�".�'`�In˝�E�hQGQ���^y�O�@��Ү{t���>�IIIy<X~��*c�A�=�����z��[�ĥ�E*�b�%H����L���}g�ݻ���)y
l.&RA9]a����u;��N��Ha�c��pC�L$ 7
�\+�t��7�
���Z� 
�İ���tB�p`���Tylr{d�}�P��$���O�WG�L���^eCNK�"U��8Ϫ�)D�	���n�?�=7/�UJ^�M�o��q�!Ҧ�mp�)G�k�?��#�mB�#^��	whl�ԗ\����8[�I��Z��oc�s�ޭ(?#5�,�%��w։��:��Y�X����i��<��h�Ҥ[zl g�u�m��*��l�U��_x��Z;�J��`�g�Q��]-y��hQ� �����%lz��.��yr�����d�˳Ci����]KK��:��K	�c{{�����ӛ1��ļIɸ}�4�{LOyJu�s�_�v�N��܈�&1*�{����ŵ�?\���]J�t����k���MvU�.����ۣҖ�[WQ8��|8�� ��:�!s��*B`��\079%����1^�P��
�0j|�RB)���Ŵ`ç�LEl���)��]�,mȰ�܉��΁3�VA�,�'��q*yb_�
�먺�=6��Gw4� ޡ6�k�>�o:/4&�h�R�ۯx˪�HH��3��j�ijj���ε2����i<�{aa�׊�olj��ͳ���)�x�<��BZ򱾓��>)F bґ��<�3C���TVYtO�X�u��,wMMʮ)�O��Q�-SB��uY_���z%�ax�X��dn��fd�ό�X%����4�����h<ӊba�vg�!k�m[�_51e�ñ����iwGZs  �ˀ�b{^�P���,�@n�Ӂg&��c

٧��µJoK��^���*�����·��Z9k�����'���|T��	?=��/|�#>7�`Y///oo>_ �o�^��#�+���H�YOo��C~lQiH����v�2��+1j���ڒ~`q[
!<�޽L���k��x�O�UVVacr����^��6S����R{}u��JC�X�7�w�4�\��!,}�Y/��J�О���&%��"�e��2�2�6f{mb��e��O�J�X����+g·rZ$:n�\4�;�G�k�K
ll�Hѣf���+����7����1P�%�IKK.,,�KM�.���!6&(�6 m���4�ޫ��
G����Z`��2�d�D��d��ɠꤻ�a�*=β���B�dJRuE�<�����v�4�f���R�B1A^M�f	cl0)E�Dk�ǰ��������A<�FwA*�Q!����+�1��hX7�DX:n��ߖ� �%�Us ��<�ܼD~��c�G
�Q`$/���Td�]}��w�!�%N��־xZ7���s�����r�� �a��O
5؁�y��ϊ���[�!��Y�C�޽��֤������~�����p������ϰ8%fߨm�bC�`!�Mr�Q��_t@,�Y�t�!��o�W����j����b�ԭE�|s:��
:��/�H���~���C�]��Ԥ~}M(�-�ua�a�aG��������� Qq��%�	�5�ITc@��ת��|rX��V��%�V��V6{�~��gQ�dhxᡛ�WL*����)��b�w:w����C;�"B}7F��n��Ο�u',t6���� ����ƼM�r�O������:"�S�;�+=��U����z̢�{T}愇^�k�g�;p8��� fww;��lm9,�O��*�ģZ�s�;%���x���t���	�����5���t���w�����G7���j�I_�	:���")�o��~�	���F= ��?��d��C�^}�a�r j�o�r���UO`�7j���.S��u�������̥�����QU��ڍ�Yd�>�-.�����t�ֳ����N-��c�g#�L����(�L��{V��ɍZǟȀ-~�\m�#�Wp�V�v���@JF�S�9<Z8���m���ލ~��g���kv�CC!��R$n�s�@��~$<H�=��g{H�t�)�����gN�߮,tI)�F����f眨���H���x6l�'VZ-! ��>%mB�D�����U˳,$S� �WμΡ@@ɐ�o%��S-�x�-H�wx�)ܽ]�����hl|��S�m�������b�G2+���d}6�ͭ�׊�F�XY�e�Z�oX���;f�8�����xq�:j���bo�thyA/��+u��bn��i����9Vz��?ML��ߋEjz�d/���!T.��j;��n=*B�ݿ?:r����r2�)��,B�NE�s]U����w��#�s�qx����;e��W�E��Ck�<�ct�έ��_2a1f��|�siT9o�0��P�*�h��e��H��9m�YW����VVV���a���Y�xAܺ�m?~0ʏ�[�ŸG4m���O>�D�}`�r58�|��,cWױJ�����D�R��Hyt�M���������3���:j�����T5.�3��.)|ۨ@�����ϟa���3���ʣ���m�<���pV��[F�z�&�5]cx�W��mU o����3�!䘸�(/>^���<)'8Dl��E����	]:G}����C�佅HnS3���w��2P~kkkra��ώ
�b���������c33JJ�@�:k�Q��E�!����������+T�닼�B�_��[�n>a��c\��A���0u~�Y�moG�����_Mےr�\�UWW�/ܧλWS��+Yw�?�v� 6������<��깿�xR�՘G�����#��m%6n����\�+[Ĝ�;K7�S"��ڞ����Bl$ka�#��8�!�kQ�:�@��*�$�Y�oͰ/ ;666i�)W�����~�计y��+�W֛�oƖ��7UmT[Y��^(	���ӡaO�T>�W�
��k}IX����pw3�DŪ�IP��>w��+�Y��4��<�HJ�a[N��fK�g�ߣ�2ݠ�3|P�p)�n�	��3��Үa��`A�|̷>�.tF���n�GV�,5,����.ZS+���"���� }g~�+��hhp���>��&�g9�����ŋܭ��?7�+=�r��p%��ڵ7l9��I�3/����K�����z�"����nwh� @�):��EX��%��Ǐɩ��J���\Vt�q�r���A�xlD�Č�r��Ub����vz����~_ȕ}і2s����)ޮa`Ca�N��.�����LS�u�WY�{܁N45�������L���|u��/N<~��=� �o�*1��0�g�������1J�a�}N�+�����Z��L�\�����<���c�t�9�th�q�E�2��84�#� :����Ʒ��:���bc�LL~��x�͉�ɚ�H�j�*#᭏�M��8�~ό�{���Q:������ַ�]Kd5�H�k��m/E��!�6����TR"�3����Ǔu�"���]�EН?��B,�V���)�����p���afn��k�NNx���<#��ꃄB�G��Hm��
�m�G�Q��0�o�a)��q~�1q�w�*_�f�/;;;Z���˕|�dgss3�(ub��}e0}�m�*?�ۊ�Lf��q����7���C�����2<��Hs$���?h�U7��]p=J[/OW2��zC)q?�q��+���	��{�: �����\]�q�j�^)l��@1"��{���H�JϮa��BT�����"+&��S���[~9그w��k:��o��ю=�{jht���:1���^K�9��6�YD��A��N�e�_��3���J��QJarpq���~�j�<��@�ĵCs�z-Fx�b��KQ��R���ݦ���f���1A�n�BO�κ�Co5j�_��G�F��Q2vm��+F!#*c�����²���uŘ##�~��+�e�H�8���'z��Rq@�O��A{biR�j�(-��w�+mD6��*�����5�հ�rc3���5Åm���=�I���������jh�����5o	=)�����,����S�zAY�Z��Vh��666�"}#�B�����ۗ�N��<!@�@?,92�z�A9A�2�e��w��ú�m�]Xr�0?n��PQ�l��?��& ��!nwӂ�y��JRq	hQ�\���к�7�J}�ț�����N�=��1q9\�l���q��K`Ao�c0��g��3|v����ֶ����_9(�cg*Ǵ|�\�,N�YR���a0rI�S&�%��;��@E¨��-F�����c	IrZ�V�'��ޱ��dK L��̡<J-��3c0��tk<�nc7W���\V[ۻAr��D5U��%�H�t~'40:7
�JX�NF�
Q�����@l�'��YQ�|�za�(��hl2��[��sx{b��1*b{�kk��m��'j�TǢ�F�Vp��Э�p���[����;�##.u�r2#y�6���|0A���󹠕���t���C]�{����GU�r�l�?)#�S�fKT�kh�
-,�2$���~�����Z�K/�%2Ad��y�Y
3@QbH-�Ņ�d×%H�G�:_*@�O������:���]5bw��'u���-QJ̣δ��o���$�l�I�M @�F�F���۔����+��2 6<�]���ſ?Ӊ\�e��[�	����5s+�p���H��Jo��Q�����]�ä�_!>��?���`�%�@�`ra	�8�������Z���3)9�3:�<���,�\Ge��m����-x��<���`��ҼHyAM�3����N�x�^de�]@��	+�NNI�qq������;�(�|V��XvϷ
�-��2������ �����Ez�vPw��PK���3�FZg�Ұ!B�/}F~~J�%X�y�*�*v8�!�b�H)��_΁=m;�.�UV�:_l���X2�~�����VC,���/ ��3y�����Cw��w�{뺊|U��b���]��
l�uu�s>�v?�679�{z��Q٘�zھ}S��r��R�6�cE�v�iO����>,'=�u[S�:,ӌ~~v楡x:G�9#����K��}�?�L��v]����H&T&y������J�E��j?���-�u�tC�t�?����e��vi"nX�Mκ��V1�?�?"T 1���<0�(�q�U��M�ZO��li[6�^�JT�����q�fA���]e�<����#�_�8̤�$ݰ>���h��qnn����b����R�0ȧ�_�04gd�s��D�V�y:��m�с�����Pw�`����?���ܱ�IS`�C-���'V�t�m�onn��y�����F��������
�z�NrU�9ץ�P���Δl�<a%�ێ�g|��������.���(� �n�I#v\i??'��9ꡮU'F���/��Ԝ.(����5\�9ȫ�k��d����#�hq�pϡ�=� ��㈭`�J**^��7-ƭÉJ�H�h�>�#�A�u�EA�9ߜ3��y�2�۾�7��ν��HQ%�L�@�]Z/:��p� FV�cf����]o� ���0Ă-J�cY��}�8�:ګ)XƹAI�+ǹ�eW��{�����u�=,z~U��#}��_S�o߭S̽�ҝO~(�,A�a��u9�~ǫ_y'=���Z�Ft'N��{�����mNH�O��x��>�P��p��]�F{w7�u��A��/2ׇYg�*�u'�ж$aS���{�4�.�>ȵ2uv&5������|��i�3`�#l��k@36-''��OIej���XN�ښ�G��qy8	�i��tli�;����s�p/��_o��kkV����Z��t~�Flcj̜<���v�1������X�єGE�q?�h R�K˧��C�orQ*�[C�R��jHxx�������c�W}6HI����� �A\~*
v�p��Z��xO��������_͎�bz g�1O6�
�b�He4�����A<���\J �ы�Rǌ����y ՗dk!6��C�Hr��m�u�L�0 �_��ƭIBMZ+8��(�B#��65E�Q?�5���5�mJ�u��~�y���o�! ��V����z�[�jB<JK�%��{�n��4!o�9�"��VA�\[s����
,�~��&�{pi��$,7�ϛ\�Ԟ:
N �YW��+F��~���p���87~Yu��^v�3::*-h8�T��%�׆p�	y���2�Ԭ�|��q�VJ��H;ͪ�qZ;��W�-ש-�G㙋�����C:"(����\oLLLo��9%@2���n��h��Rq�"��ߋP� ����9a`����%��?�wl�?$�'�����O������ڡ�;P��F9�b岁�"/,�ʵ \*�
��n��>k�ӫt��\�"�f[â���g�v���3�''B�2t�u�ǆ��=�����Z����[�a��������š_��3$�*BI#M�����瓞?؟�^�\_rl@Cub_szYwy)�١�˕#�O���+?� @ �b�:��s�}��0;x�\��9�4�f#�Uj�4���Z��
�֡6��A���]��OĠ%�}��t����L�C���2U��S�G�:q��_��,Yp��y �����{�i�F��L�/��܉�1h�$J�2h�th�%( ����B*��R�ƞN7���@Ø\n�ڪq�*���FE�)�C/�y"��3�J�Q��N�cl�-~beo�@�ϵ��B�aRj�&�c_B����{�����_�	o))+��85$ JDA�G��5K�Kz�0�~jn���x,���u�q�ş�Ks�����F�$Uz���葹Vͪ)��(�d�9�<2Nr���IvI-�#h ���(�)��_��QFm�u <�����;���|�t
R\��u��U��X���:��r¸<��#����j8l��9��ښ\@�$*�l,Z���:߉�Lׁ-`��~@i�M�����<���\W�Pr`�:{��n9wNpa!���n�4��#�x�"d�-BA-���~��;N���YU�6ŀ���a����q�'��3�#�����"�|/}�iK/u�dJ"�P6��
;JO��l�RA�6���lL�N�/;�n��X��KM\k�!��'��P씦o[��n��X˘@��XJ�S�T�09W󢢢���.�c�NU����m�?�0�닒��Q��q�-�ؿU|]^QA��P-q����:q˴_����5�Hkj�n5^�Y�ت��U��<�¨�í��{������(�ȩ�v����}��=�-�A}l��E���O�Z1�l��p�z����=Mt!p�v�f��=٘�E�B�����Zh-���	�V+�x��`u���'�.���T�<��nw�� ���*�O��t�:Q�E~����=������q3�.�h����{}�U��Ü�Q�A��Q-�[t��a"ژ{P?�B q�X�)`�b�3��>,�N1� �������A�o}�6u��5�\\R��O��;x(�.�:���6�
���~����1XM`�9��<�L�
t��Rt��n����R�z���]��.�uUJ銱���<�ޯT��g8��ed8lBY�ϯӗc��,�	.�@9<8���`'1�c^�X3<�L�HOϢr�S7��M���H3K��˦��F��$Q)҅au�W���f�*��oo� �d���_�0��{�ڑa��v�-��w "ם��t������ro����ʁ�bCH�$G [N���=.���ˁ��ǶZ����Z�4c�݂^ �PQ��}}�?6 �ĝ��v��Z�` �o� �\l)�"�����nnoW�Xxzzf:�U��D��ޯ1)�(9�������( z"d���&�qC���{ѥ��N��P��!#�ƶ^nnn��跱G�t�[�N�WzC�rt��2��v�<�ꅅq�I]�����T�5f�u�/��B�F�v�8��zq~�C�S�����~��O*E�3+��d�:����d���,��JV�&�X9Y!'����3��N�O����ݺ����^���?���y]�4gD$�S�S���;5/��!U�P��_���G�����tx/��Û��撒L��f�3!^Iu����w������1R�we3��L�����t�޸n
���t�ni�MMςQ�s�#S�U�U�
�B���S��7�9���"� ��#1�&&��7g�eˀ�9�iSg[�or�x4�]bΰ��]�\���_A63p���(=h����@~oTK�Ω��K�A����RWQ�ܳAI�5#���}�U?�G��0�ozr%���-%�ס���h�V/i�'�H@4�r�O�n���W�~ax(8��vm�e��{��!�䝝]��r�{�V~��s��!����N�- &��k!/>��(��#i�;Zzx�PSS?�oΘz������ڍ�0Y���(����^oc�,/�c-�$if�M~���9���I��O��)wo4�D�oXC�\<[�Si�ʒ�֣���L���ZYM�t��?�:5�(U��ca�~L�ߊuV���F�%������N�M3���&E���Ӟ�w��M{�����N2.�����ߵ�T�5��{B�r��51�X,��e�>+"{�4hnk[�"��SU[;�����fu$c��}�x�V7��,&tN����}~�jdÉ�[DW��r�,z*?q}Vm����"O�I=������r�E�jz��$��2�|�ϲ�T��p���NxW��e�����{2���z�\P�}�'#g��F�᪥��uJu�"U�7V�p�5��!��m��c���y�s������g�(�g�w���ش��N����̛�j���S��;������D������=��ߩ���'#x�����_}݁۷e�w����߷�rpϮ��G�9�t��,�\Cg9&�a��)�(�:��Pp�#h#�����
�,�TG���H~zT�U�f���c"�^i
JL�q����WyDI��3m�<�H����L	E1w�S��:���/[����kr�k�㔏NZ:������R׈�c�7��<���S��y�������V��n�3G�ܤZqb��㺝z-��?oƺ���T#�[�++ww�A60�
k����R��)�||�=/M�3����ƾK�Z�j��j����m`�ٜ���]H��sG�6b
*-u��Z��s����� �-zއ��-?�w
�>�4y��ڈ�O�C\�r9&�>���Q(��2��ޜZS��F5 �8����Ē�h�ν�>����������M�8(�	}���d�=~��ǿ��&��(Z����Փ���j��j�W�v������J����V�#���KJ ���=�鴏���~6��G��B�:���O��y���H���w%� >l��=�W{�+@K�į3T�ҟ���7=Lޘ3���hrPE��+�3���,(QT!z��f�<l�[�t��aFx��!nr.���\�؅�1;��y�(�B����e+Dh�U�Sn�sƐ,�u,�l64y�gk�g6L��r����ʔZ
H_
�ٹŝ��/P�8S(;���Q\������!M(_��}���Y+�7t234\-�C$R�un�tM��pt�8(z�Y)�ˊ$�`��H5��c���pk�ҫ���]M�%ݷ�KJ��� ���(S����R`[��D�eQUIb�ҍ���֝��-�����:J����ܠ�O��гe���!=]ݠ�%������,�Å���9��FC��:���m��l��`0��YxCo0? 2톎~!%B�i�QK���q./��_x�6+�*4�V�YS��*wGXPJ�QvVf0�6/^�H�Wo��V�m׍W@�Z>����&ϥ�ZH*1��_��6�gA�j����שA�܍�Z�z��LL�~�l �O�T��+l�����GAn�����=d	�����4��gv�r���)]�]��}.d?f��ż�+� z�Z�4ٚ�k8!Q3�t�7Ai ���ŭ! K�.l�26��]�)=�����~���/�
%�����ᎉ�|č�e`H��ݿ�
刿���_��쎴��#���\*ְ�5�4)goo���Orp�[ A��Y:8��$ߑxB���wo�5��z�tbnF|SGG��j����#70��$��I��i�\_���x�v0����i��'K
/KVyMX"�kt��m\��~
����(�:���e���4EΚC�A��L�yp�>��h��Ɏ
��7�!J�I�ַ"~=�.���$�Fyj�8>f�,
o}Q����_��:r�I����x�-96��k$���!�=����g%k�����\�XN{�uC�����Ov]b�p��ۻ���*�n������'�"BB�O�ހ����XPX�lcc�_���,��$nnn>�n=$upt�ep����p'��=�4���xj*c��+�?�����~£r�99U�\��LZ
l4�y��9��v�������*��o'/��0�|4Œ�F�窪Pp1��Y�ć�H���؍����i��������%��v�F�?]�E���hV��X�$�ag�\��p
y���uA��0�n7�	#}�o��.2��z�7g���8���a�ܝ�e�f^2 xc�6�Q41$�2��u�Zyf�zw��%��?�r�@~�6��A�9����A���K�NWRĆ]�LLL���s�J�Z�#77���I���!��������-pj�G�1�(^����((�o`�D�$sA�}�9Ec�e36��E��>�NP��\!��ѩ;�s�m� P�M��vǲ������C�k�� X�F�`�Ι/j��oL8�W�z_=��NI��)h/xq��;7A�ip�SA&���+E ��:�]��f�MA�U5�x�ￖc���A#���l��[oYp�u�U��v�Ks�昲^Եl���<�k�Q��*�����dU�4��F��6`{�p�����z��-�	����IPQ�Z4H��Rn� �J-AZ���4�	�U�A/z9/��!*���.�f��k'f�$V:�w�M~.��3{`{�'*#��_MY_����/�S�2��� ��Q��!r�||<�Y�񦂳���k��|?cu�II��Ys�G�o�b^�j��$�g}�Ζ2Q9L2���҄���E�/���I�!�/��/gəc�#�����W�o)���!w7�7'~�U�LU����!��}t�f>�7��CѺF��}�4�7 #� b��7��b��o>��R9��䝠d� Z����[�5���,e���	e�h΍�P�ߠ�����3�q���a��~�ю<|��	˭��H ���"��䇜����#W��}$�urŷo���Z�q;CAtf'��;�C��N�T}��� ��{1HMI&�O��ё!"<^��2Z�,��~��t[���;���M({�u矷�C*��x�8;WZ'�@9B}�G|�	�6p�����͉�<���%�e:z�4�R�>a��y"I�u�=����VQU�=JpG6�]�6w�i�v�8oP��/�D�����l��͠�Ԡ�:4��E)A��F�Ϻ�q�:	��ng$5�>?�a�f��g�dj��ai:$��ګ����]O��$�o��PGlV���J���ºb����ƿ�P�6���׫jj�z�$�'��Z��L��t�NA��Ҁ�D��l쫑Bubݺ>C�ZǶ���HsO�t,@�Û�ސJ�]rn��q�ҿT��w]�l�H�o�vthq��y��L6� ������7c@�3�	Ys����H��0���&uiF9>��[��]=�`�+;�̾|���O�#[��dāMɀ��!�6���P>eD# !엨��/����o���#���dJЇ��$�/̪�I����Օ��a��(>����p�y#�F�3J���|�����m�ad@r�ZDO�]>��km ���SPP�Z�\�HM~'���D�܈�����5��W)^o�WQ�����eGeD��₸��B��{F�i���_JG��'��w���@�#|0|���3ߊ�;Gѳ�uŜf_%pс�q������P�`�\��TG���n�)=C�5E.�}����WvYοxߴ�XJ���M��=D4�k�e����eb��P��ۤoNMM���*��-��e���N0�q���h�D�@��-��M���h���t��W�C��y�@ڹco����tKp5U�78x�ĝ�6Ո�0I�OP�~�;�g�v��-��绫�7(.�O?{w�o�Q:V���8���n�0o��fhZ���l�ߴP�ֹ��@f�>W?�~���&Whe����3St�H������)"���K#��K��BZ�������L�U>4:�)��;֧�#O�8Y�jz@����Ɔ�8���:Z�!{>�[��/�����l-�E?$BX�
�1V�k��w�k
g	<��,(���,Ҿ��ujjjR5�Qᜁ��{{�� _z;�����#Hy�������/}_E�7"�g|��)��Q��B��������Ǝ�.	�-�'a�0��ܱ�Nf�_�J�*�J(fɫBf�AZiͼ�ͦ����xc����q��`u��[��X�ζ�M��%��FR�,�z't	����-��������A3���+s�+G��Q��M�#�uE�{�&_>mk��o.�3�m�d!#��o{�߿g��WA[�<�UmM:��I�e���s0������ ?�a(������ʊƁWXEN�#�n���6�d��D�3�|�������K��R��9�[s&܌,,�^�{���'B��=yr�+�V?{|�� ����|��n�ЗČ�{ŕ;^g�(�ت�w��!"��;f�j��McY��<^��'{'�
e�6��� �������7.h6��Vn�X;�} ��7�������BY���`�,����z��P	M����s*�F�����Vnኴ�{GE@$��G~��ʳ����!MI�ss;~�(���?y�����uq m�z�j8;^���-&
h��Ð�o��䯍�۩�@�J�ӄ�˚�/����^��_�~��ߎ"9㟪e��T�?�{�;�I@yK��t��CF�BMǭa�O曕��Q3��eƍ���@���Ly*w1����U4t�4��*+&������_�w�ڵ i�h��
�!�bm�v�A�۷�7<�}�Iك~�G�.59�zsQE�����âj*� ����-��?�nL�`���@5Ry��;�EZ�?�2�u��YϿR��7�������g
"l�����ޭ�y�y����y}�T��2e�wyk��L�=����Z~�*�;���6���+�ӎ�w�� (��h���T'�j��C>1qq����9i�gll�c���T�N��+u��)v��p�?SV'�q� �zJ�N���H��[�~L��w�����|���ΨM��'=-	 a�}̗���p8FѤ�d� �G~��I*ŬA�;Y�n;�����-J�y�A;ۿ;>|�H������n{�6��1��5�c�Ӿ<AK�A��h/��:����.[-X�Ŝh�L�hSS�ܤ�=}�S�{	!))���Ь�y�|��sĎ��C��t��E6,@��p2�V����O�^���)�����w�ϝ����HM��U�q�/��0܃��p����g�j�\�|3�c'k���9���O��	���S�B��K<���{��R��:Qέ���޵PJWf�2h�t������~)�_�q�H3[+ʉ/�{�,,,J�~C�/�T�[-X[7VW�˗�omU3фq�o��� �f�4�h�y���7�EPt�xmL��W�>�|,(��#'�g}�)� �羅��\��%4�P�Pͼ+�����`iv��_)~{t��ܥ��z�]Ev�`���MY�}�������}�I���k(�3#D@c��
.&'W��CZ���:ؙ��T^"�9�4{�|�����:S��=����\G|�qG�2jz����!�6֊����$<vvM�ܠ��p�����!�21�^�I�A3A��)2�V����Xη����!�t��#
~�`�ُ�e��}�2q7�b�E{���]��S�Վω/������%�QίE�QK�����/
���|7����N�6ݳ��饌#G����8ۯt���Zn��VH�}aho�O��7m��om�%��S��hMjg�r��Ѭ�����W:I��ލ<�:���@���IWU�E����#-i�s�^x���rF7��2ߏ���#��'���ăa��M�q1��#\�1�>6�"\�xp�D���#�!va,g�i�b�`�mg�U�z;v;�.���.�*}Օ�Έ#��0�����t�{mj�|��Haފ�D������F�F��'���@M�&b��O�u��3�~���hcs�_�q/yV��/k��w��[�k��>�ja�M���h1-t���bSssLi��pJ�Z��'{8Х������zgD��`�ðZ����Μp�$1�M_`��8�h(XQATt	B�Q�]MXb��ܦ�����r�ӯL�0����k�H�z��O���~��k��w� #�C�x�Z�����^��{����P���_�����������r�ƟE����t��=V4O�+�e����N[�n��F�-�Hl���E�jL����#��g�YG+�Q\?�ۊ�7�l�F�@س�������0N�%	0�[�h�,�Կ��w�G�Cr��ozOzv�#w1�m�z�&��~��]����x��ܘR���Q�S���ׁ/��e�ɒb�F�Pe�Qn�!7Ĺϴ�^w��H������^}d���h��l1��{��7"���+[Ϛ�jof��)��h\��zy[���I&eǛ�v�!��/Uu+��݀�d�����D�!��3*5�FՋn2��j�'����l����n?�����M���I.���nכ�w�6ؖwV���w?��r����~#r�Pj�I�5Dt�i��c~C=>Rp��JM�^��/��a\�W7c6�>����"-4��z���j1�|c��@i|ì���w[���U�mA����Ѓ��
�f��/�p=V�a�&�(���q� K����`eV�B�&�U*[�D�!'ߎ�ר�����Ύ���[�I9;5���_l�#$ߛb_g�K'�ښ>m9:����Z��E�tlT^�%wl#��ן�ՆA�dP�N��'��}U:�aJm4 �O&�־Ξ�7�ė��)��>wR���8�49\�U*�V�-��p\3���aG�eA��-5���8i��������^��T<K����4| ���6�c���U\w���2�X�Ʒc�|��;2]�ğQ�F���wo�3��f�g:��D��)�P��=WItH$�I? Ĥ�\��fߥ�O"Eoͪ��z	��G8�K�\eY���[�. �n9��znũ�A�;?{��U�n%��\�_��A��fi)�(t^iY�/���l�<P�%�����B�++�_�z����ꍏ״�T�����_�%�t���o��pnk+�zf��$P�XB�Kgɲ���J=6�8����\���`��ܭ��;0Y=!�����Q�E���6,�J?�O�'��|M۠���T����9s�.��G� vTN��[���,���)x��W�5K<v#�	�^/����o� �^ZI#������.\l�<l��<Q��E�	�@ի�?д�[H�y��ړ�(u?���ޗ��/���Y��v�QX�A0�o�B��4=�_�-�}�~��鹒r�鹋�K�Z��v��ho�b]�%I�Q���(�r���9v�e��	[1�%O�Zt#�{�4��B�f^�'��oCNk���@|5|S�O�dAU�B}�����m�f���_��0%����1����_ט���I�ֈ��v�BQ��]� U��`��_��K�/��T�y������=:IG����y%�
�h<�399�cb�wp�=��wj������@|����:ڞ� )�mjjvU����q����@�efff��(3��Z�@�J˞�)f�;ڢ�΂j��߸U��q�k�W	���r�ڿ��=\��+K����� 66��yFHC�Z������WA�l�1��m����/�0���naE�c:�w|x����+&�Z�+��7{�Nq��+BS&���׹� �9Y�0�I?�|�R%�����P=1��-�[��~��2 �Gn�pw�$X��J��I�ʮ��O�I~i �>\�j�<�a�6a�U�F+Xwv�g��d���_'rꑲ��/�Mwz��; @�[YЕ�����r�ϝg1�?���tr�6�h@'Ѐ��ۚA{c2܍��Z�'��}y;W���/�� 8XI�y�6�^B�Y��x�Y\�p�5�
������컇�t_޿�q�_-��Њ
aA#x٢S�(ғ=��Mf'6�3��-���U�Y�+־���0p�7�w��0�ۓ*�}��ۗuv�G���6n���sL绳x���3 �Y��	��+�>kG@i�k��A�pa�2ئ��PS��O�%��;6�s@����H:|�*ň���i'f;A��^�������V$��������T�𓟪�$ ��*ɨ懐Z��Տ�H)!3�]�\q����
]�O��o=C]�4eo�z���7F�� �Gӑ[�8#�F�G͑М�yu>��#���&��j�x_�oƩS��=Ѥt�b\����$Ü�!����ðں���H���_y$s�E@P�>�`�p�$ ��G�4$�ҥ]/�o�9*�n��Y���/��(�`&(+�%���_��^�!Z�_�wDI�-��!P�h%�Ϻ�Fn�r&�z���X������Y�}~4�F	H�z�Ļ`�$R�\���Qd\A��C�>t�(2������y�^�=I6�Gִ�
\DL�z�C6��P�6 C~��G�S]�c`$�����3�ne�1�-� IMM�A�tρ���D
M�2�	:��l��
ea,,Q��ŉ�:=ԑ��fӷ��U���xQ���k�n-/��	4PK�����#{�\�o�(T�o?����������f���AlYzy����W�
薵@py"e>�Q��+�-ǁ��b�ew,�����=-xZ��ņ]�-���o0z��_I6�~����tX�j
|�o.FJ�C^����_���gB��?�������U�V���a;��`����R�'��-.�A�t�)Z��s��˗3�����A�l"��|
r%K��ԭ�C6]ʋ�&�nL�Bƒi��E���f3wH�C)�?w��bQ� ,Y�W���>X��7��M������jw=����?4WD�
��dxO��M���k�ˍ��M_V���������ysy������#F�#��PfcX��$j4R����a�O`'�<��������JgU�pz�/��@6 �nG�spǹ��[x�R��*@���ܷp{�*��WL���t%��)9�hBZc��0�Ai7�H<Bz�m�zy᧪S!�[��s�@Bis3nxee���񚯒MIR�Ȋ�էH���kM��@�Z�77�5�s������I`��4�D�+pi����uY������@�W;L[fw�������Y��ա�Aӝ�tѿ��`��6b�>��nD|Xk���k�ͤgI�8����� ���S/�oi�Z��v\�x,��K���@�7 E4��F�U:�CG\�PpOo�v�܄[�h��\~���>$�}S-C6��)�yf��3�q��C mႹ���uv:��7�W uo��~/a]��A�W��G����M��@E@̟�9�>į&�r�x�E�8�$1K�t���++�ՙR��ώ�*���]����N��_��i�F��2.��+)�0��k=���}58�Y�����*�Y�.m�Q�U��O�u}��o�l]gR�/(����$c�fB�&'�8��)Y�h,��)�����c;�!�9�����.	����+y��SSC=��5h��x�{4{�g��J'3����7�^��ɔ:1���ُ��*����>҈��M(����e����@qL\�)�@[�h�w�ܯ�+/�O������ؒ���5����p�����~��X���x��2�ߺL�
r��Aruc���X����K��ٙ<��ͣ����d�{���z�I"ef�A:z&�@Uyt$���ns`Z"����ۆ����3����ݍ�lv�ɕN�����,� d}�pC�������&��C�����N׻/.F�C�[�6Z��HS*��kF>��-�����������{M�gl����v�r�R�?55�{��b*���X"�]; ����1���p&:�o719�(����pm��:rȕ_�~2��ۯ�:__��ʴ甑O�ep����Q�#��$���h��U+ ������l�nWQq����H(ğ֚Z�^�j�5;S�f��7����?�+��:{䍺O66��߿�����+0��U��m�����}��s�`i@���X>�N�U�����ѡ�8�0���ƒ�����9��]�z�r��|I�͒�!���q�z���p63w	�`� �����9���Q�����F��:���<I3%tyrk�f�&��I?��<�
��_ؽ/����%}"�Z<�A�E�^��N#�h���ޘ��Ml���{�++/���OՅT�_Y�kH��(�(=dF<��Z�x�g������f�y�۸��M��WB���e-?��d`a��u���0�A�����$=��3j�_�_y���`�PŤ7����|C�k\w�����ǈ8p1��n�rW����C�CKbw�i�5D��V�|B�v%�ges����6{���[V����=��+��(7�pӅ�Kt�� �g؉ع�����#*-��U��c��k���|����[�d�[�IO��-�?��f'ʯ�����������J�3�#+����Ϡb��0��ǆ
��t�h1̮��'_�KP�Kh�/$W�]C�Y�O�'�+��$ӑtË���'NlLL�X�Zi��P�a b������G���>��7r6���]��u3��o,HWe��Sn�_]�2Vl%�@�~A�3��w�"3qv22�	���y/���ex}�֣L�hL��e��L $��Kc�u{�F���23U���@��)�K�鞪���P�G|xƃ�{}o:�v���)�X!W�6~��a�����l�R��_�L����3K&��ZkF�݁<�F��0(�K����������H��&�}#r�}Y�k�5��Չoa�0@�5.&�u����
w�
�OPs&&&����|Yn&X�;��
%��G#x�c��4�	�bz{{e�=�YJw����/A�Z����������F ��B�0I�˃���g_�"�y\�h��L��WB�X��b��K�DB��ȕ��7��~[-Xk����K�h�9�&�V�(٭6O8$�n\�ǿ��9��eR@䭧�L��������i�0��zǴ����D* ��K�I0e_}��	��ʁ�A�z&�����)��q�Yy,�J$~m�phO<�ĵ&�W��Uc����Հ����x=��{ʵ�>$b &���7V�#�l63-1%i*���� ޫ����n�@�T}�E�w�!C����zo�6�q�J�� ���S�8�`��7M����.؏��L�O$�/���3�]H¿l��F�No��A�Tƹ�����d�W|�/17Ͽ�Q�|=�����X�r�W0�`%%]s�V�S=�nQC���[�ã�[�k4V�u�6���w��	[GՋ���ä֚������Km����~�S�8t�453��H���������93����k��7�76�~��fZ������cn(�WW�Ժ��,B����ԷWݷ��������<�F���;#���q�pY[�f����g�N��������;���6��o-=�	$H��Bl��g||�r1A&���S`	�	��d׮�m�����.cs� �����&���+�^%��
Y�Ɖq�\�&��0Ծu�NglT=C���T�C�Z����S(@�g..?��ֿ<�����]�$ВL�¯���sQE��oZZZ����J�S��B8Eܵ���NM&�\Aw��I�w��yȖ��Ү���	���W�"�߬��L�H�����گ��r'�"���;V6;x�.A��J��倲I�z��!,ֆy�T��Zc�b���\�ߪ�R�+Ap���χ��S�����K�֘^��l�L�F		І��bP��n��>G�q�����{�æ���F��"w��g��o�]���#[�m��C��/|a>�a��+����\H�-�i�	�u�O����iHZ*�*� Ɨg�k��?�!�6g��"�"�����:e��'�����)rY�/��f�:�E��{������~������}����B:�S��y�~�+�,�2 ��2�Y��"��ӵ�ySl�|�-\z�����,I�V�0XV}x�')��˪p����,� o9@�y}jf������8&��u�+��ԧۗ�Ī/�mO��{*�u/�D��Z��2�G۞|��-�0��CF��!��%'?�u!#����+m��eg�65P�_U�F˗��������Q�Vc�P����5鑰6VII`b����XYY_��n��f2��ň��#�S)6�pe��,����EX��YA�f�2�0p5�'""�"P#���iN1��2�b6�e> �E��H�@"�	��)���d�K�/qw�>-�~��Ȟ�ma﨩u���^^p�}/��=�$�Ϙ/������5�b�60� ��l��ek?'_�fQ��G-��= 5��PuY�7V�?�m��͏ؒ`��EdM	�x����Dw�t� >�t�T{��$�E���;K,�>�-x���B�p=K{�����C{?0�8j�����6/q�����g�P�����H��?5ݗ8�)��~�2�,�=k#��q;�a���K�Pr��|Z������yf���7��c!�^��3�ךM����os;��zv�н�i#?���m?�A�'��������W�"P�j���%%�l2n�ۇ��u��;��@0J�k���$��E��op���@-�d�t�pk��~`�����/1<����^c���⠞��q@E+�Q���+�1Ar�����y7��O*��c6=�JB"�l��Y�S�@-H� ��!�[�P���w���z��(��Y�v������.��Si\�K�̅�8U�`bӌ�@��=v����yZ�~�ݰp��|}A/gk(###�v�蠲Յ��&��1~:*��LKr	�u�k�
*���`f\���y����\�͕b�X�ꃯ�bb��A���N΄c}�c7,U<H�2C�D},�u ��!���b�?���I֭�1��|n��*V
��a�k�]�Y�2�6q��A�/��@0J��
�������u�Fpr���`�K�T8�H��˘v� � m�q
���"!���5���8n��{ԯvY�?Rz��L�g�s�#J�Vo)>���r�]V�=�b���/<d{�YL�7I�W�7���Hā���A�b�����9n�žB 2�&H|���D��cC����)-�]�jJ��׺���X�W\�v�~ΰ�KȩyC2���6?��tK��V��%����M����1qq�����1��&z�o(�}Kd����/���ڣ*�:B���g�6��@`zu- ZP�H���k�\�z�<ގ�f�CN�z��Ý��ʕ��*��~#O��<^�9J���6`��c�N>}[�0�*��*����Ҹz~�o���o��YT��q�kiӶeVb/e>����@�v�� �u�1H��rD����[�3���h���߿PK�^�ZȌd�5󩱤5��V�f8&�=H�,!<�ɞ��;w3k���B��؆��`zh�;G�g�$�ذ�����D����I��������Nn�|�3i?������ʩ�R�Ɗ�:Y�|�{��K�s �@g�#{6i��{��f���[���^�������
���ȇS\������,@GQ1֤�K�������2���Hj�i���{S�/}2�h�YT����q�'��}�V@��g�ѯj5�5a��e"U�����%�D@mg!��%��^n�M{�D'�#	���Y���T�'կj��a����"sF�c:����"z����f�,%%���)�7�b��U2Cdbs���K��l���f�c��&�B�Ly�<9��F8Qz��m�oߊ2»~���>��I�6�*J�f�ky���p4Q,�h=q�!�r���&�(.��b\���yh ;"7�L��wZ�ڤ��5�E���٠��N��myu��q����[&�ZJ�Z�Wc�ZT ��cp�X�SӋ�l��pJ�Z�sVz:����o����}	Wց�QOI(*���UV��_�i-���n��x�nV��i�����ɤ�5322���:E]S�(�K��D[b��)���%xM��U0�do�lCX��|gdwOSm�O���U=�u�oy��]���/.�B���r�����ϵK�������F�du��Ӝ2�7�l�X�U�"��X�����o�������'���J�dK�ފ�YXG�-��ک�k&q���ԴO�p�bk��	�i�ڄ=�#�����������~V´H>��������69���x���ʠK��]��ec$6���wC?=��Ez9,���uvͬ�*��Q��NoJ�͌G�����
蒲o��U�q�O��f6��zH��3��H�.tr�ʅ�ޏ�Ԅ����٦���Q g�w�<�}fcc3��!��";i$�[��RNS�"���������yx�s<�a��1�0�rx��!��X����GvjcP,Hɰ����:�:�n�B�f��2���`��(�	Cn�
��.n ����[b��x7$B� ~��G��B]M�u��kȳ�\p�f��x����i�1f��D�:�u����oV�]�u����ݵ�{\�����y�J��>LUF����U:ؽ�u��2�ZZ9�����ks�����{M��Y�ҙ�_��)��r�	j7mC���4$��:��zOW[����7�܄C΍�"�8ȯ_o!�a�]ⶣ���!Y?�\t�۠A�"ԃ=ơ�>�+Q�>�+T�&��="��9W`�Y���*�6���nj��q�l�Ծt����-���/����&!w	I`L�A�E�iQ�6�o���x<����$!!����p��6JL��gK��3��H������B&Hk7.J������N+�PE��K��?~�0��ѭ�x\�=}҅������S����i3��]מ''�7��3����ӭ��ٳ��-�LC��X4]��GZ׮_��˓5��~��(&�f�!��tX�U�ș��[�!���<��>�f_�v �u�z�z���������lI�,z��KV��3�x֦�$���f��_����:e��	seW��&�,5����

No=ͦq]vD_�V�i���2#���A�Ѳ��M`	���7sҼI���֔�Q�$�g���K����ӍD{YYY���z��i�#>d��f=o���M�r���Q(&c�Kex3���h����|�5rs�g��o��_�]��f��ڮ���k�i�d'�Lq���Ϩ�o�,��p��۞���H�/]����5��3�3���h��p1{	8��	��v�V>>��:<�J{�y���a&�LЁ2�{e�����,>���|�{�<s)c���A��Hu���U���:�����tUYK�ߟ�U�E4�f�v+Og�t<C�Ҕ��Ѵ�!�~�Oo��Z`���x��<�}�2�����妊�ñ}�Y\f&ky`�BҴ��Q��dE����im-fdD��ib"�z�߾,���1%�&s�B�c�p��W\�1��#%G�c�R���B=Y��?���z �8�����Fi�)oiɣ�d�GR\���öp�����p�RǓ�p:���|�ȸ^F��n4�[�����.����T����^%���955�^�(@�1�ۻ�j�w�Nd���1ռ�9&�*K���4.q�/JIr�C+�ݴS?|�"�\����͆/Kq��{�q����.>4�
o\.�)�����]���~uӶJP�g�q�-�&i/�X��F�%A���=�ா����B�4� �6t&��䓞3�uP��u{)�3�>��so?���@C�O\i�s�Fd]Պ'�7��	S�B���B099ycվ���ߎoو�rT��>P:�TQQ��~uMW8exz���56&��n���3�[�φ�8����V���/:e�7	Q���;������́���㑴�3���y�,��@���Dih���i��+D�蘾3��yG��2]96��y��VB�6gQ�R0wu��G�Hb�b�N��w�Y��ل���Yz��o
�Iժd"^���oB��,��%�WיB��.j��� l�k^X���J�8#�O3�BMN�t\���Ƿ��}jf���8`������輟1��y���y;y�	�Xݐ���u��ϧρ�6�?��trQ4��a� � ��Y|������&	c�� GB�s����	�����*����%���۵!"$⭖�Ω��RÀ�[y��N�xT�=��[G�jL�iW5�CVϓ�㒯-�e�r������˹��ma��ӦBW75�������9�dl�o���!�>қ$����Ǉ�;S��<�"g�m��?뼔���H��Q������7����6����'���sk|�n�o����6E?�(?�:<��TK)	'n"q���(����;�↖��`����v&怹�ݸ����@��f�U�͛G��z�F���~F{��O�RUo4^Z[^�e��!���|:/q��1�v�}ė�
��,`�H�_#��h�I�aU�����P<&�����I:M�o��_x�����By� x�Bd�&R.�?$K��9h��v�����Q<M�kg�\r�.�g_�m*��V�_���+b��p�b�bP?��{��N���Nն��&?��շd���X(,J����i�!,���X�[�8.]6�?#5��.?��@V� b���+0���&&&�ݯ�}肍��Ӆ�/L'/�,����j�{k���-�h������|
�?�����s����������98�Y��q��E{g�F��2{\�wD��ޖ�a�L}w<�����(!�ޛBR���;�W���3R!�؇�ñ�&��X!�����w�}�?�(��u^�9����`�3*2�@��S��6}��U�1SR�#?^\W��8ꖨ���~��yk8�����K�~nk����J$�*+�ӧH$�",q��v`af��ϟ?��E����6l�*B~Z�_Ý(�dez%p����*�ȇ	�k�C����1E�Ά7Ȥ�@���y�����_�����GN�7y�<��IQ��z���_���w�/�OZԎ�$U��(�%%#���K~��E��Dh�������ʦp*�b�c�t�W%J\F�y6��pO����Z�ڔ��J ����_�����)�� ��]vwt��ƥ6蠒_+Rp'���Gt��)���/c6H�N�a��`6��W

���3��[=߿��x������_���d���]��a�|1�G�ٓwg�q���C���"�z@�xMeE2�&x��K�(�`z�x��P��kt�5�l&~==�N���ź�����gƾZ�y�J~ڢ�g���h�
c�9S��W�6�8�7&A��g����<�?R��'cUWf�w�S����U�YxyѢ<6F�?� �G/�}�����R9�}��Ѳ����(@��]�Й"��TI̍��7�P��0}V�T�~8��C�����a����d~�]���YY���y��y���`}�����M�|��gcQJV-��='�yP�����j��;Z��>�a����	R�[�;4Y���%/M~�����dKxf�����wcD��`���E)��^��-�C.��S�ȷ����<E@):-�����V
G\U-�;�'�=��Z��D!,����QN	iizI�����S,��?,�mZs^�(���aS)*���~��i���?��3.�E\碟�u����
����0MV��+�؅�SU�f���?��6��V�{�RO�4��A���]7��L����������8;kiV�p�,;A�-�F�rp���!6��oibS��1�23�����ʓ�bF9^����Vn���ƍ9/Jf;XI�@QQq�/ �Po3>*�0��`�=n�777�ߣ٭H{�{JڔW�r�aװ1J�J]�6��1GG�I�Fru�J���1�S��c!��� =I�Wr*�x����SNhr�.���7l�^<jpY�9ށ�ևþ�I{?�^��Z�=���^o�0V�?��1���ݭ89��o�x��_;��rQ��ݵ�V3A<��x֌*aƆE=��7X���{���0OqG������g���+�?U��U����Z�z\^.s�݋T�x�\`
�[�#��J/��C�d�>���޻܀,�������C��-�����.5I��,����5����5���W���r��.ЋC�w�>��Sq�ϡ�-�;Z����z��>'<	ʖ����ߔh��&���̿B_C��.�.�v�žt=L����(0UU�U|ޫ��c�b���ﶗ��P~�ɲ).��mCG憄�4f���QNVۣs���Ɗ�nn��3�P��Y;�Y?!����9��J�&�0e[��}�C%�Fô�+� ��,.�OD&���@�nh����x�~(���m��4��'�(����s�h�%���z��3ظ�_�a��/�P����2gIn7���L�8�L�;R�`W1D8��Ow^�B�^ܥ{�������m��9�r7���]F�^�k[�������kRѩ'>���}t?=ݵ����������#rӖ��҄����˴U�#Q�Yg��ir��
B��5nLT�ޝ:�3��{C^�BAA���H�~�75��^���f'�Q_O���82�Tcp�ѣG���nS�R��5��c+�GY�����_���
�4��u�iK�i�5>�./���',��η��g<�y��x��#[�F03Li�Ԛ�q�i��SCv�#�IP�vx©���H�X>K�V���������~��H�fw�6��B�"nߩR-�]4"�u�s�&W>�!�z濶���%x��N��p�O㧑b$���$�Nuv�I����˅֗�/}zF�?�֍���#ٜ��q�k��u��]8�2�612�9=y%�R�EM�U�KM����#9 X�U��n����������D���FI�ذ����O���͍zO@A0��!E���JA\�W�5 8(X}�����v�V�Z�`�����l��Y��}cܭ�K����S5��HOƛ7��^3&l�Չ#�z<C��v"X	<�F���ng�{M�מr �����,��{��r����e�SL����C���8��)K�Ɋ[��N�h���q�r�U��������NʇG#U���O6����%�=����g ���g��2f���b:]���:e�,��˹�m�
k/�"b�D+�$�QL�������Ш2�_A4}g#d�0�=��uo�ex�����(9�A �c��c\Kۭ�����zᗝ��ve�%vޮM��ݬ���Iy�w#�����1aA��:!�3�Mu����#^mv�WV�jR�=�ْby�y�����JzŰ`����i�:l�'��
{ӓ��u�M�R(����׻�ύ�2b��g���,�3�`�m����p�7;�!�.5G�ns>m�H��1s�߳�J��&~C����{���3}�1Guаz)!T!
τ�gr������!��1���܀��@1�B����&)	����ܲ��~���=jN�YFo���c�V]��-�y�f*�.Ѹc�F�q�Q�S�G�I�����elj�=�}q�!IS�ݤ2@Y��M~	_��&]kn�mg1�O���$����d~��2�ޜ���J�Zi�js_-~4TZ�U�-?1]�{���{L���ü�a#��f\����;��o�*���CQ�F�8��:a��E Y�gAK���J���4�����Pw�z�NM�/��q�%\gD�^�I���=����\�_�`�n,�&�*>�HpΓc�ݰ!?2�{�����~�ߡǄ����	�#�v��/桉qwr�}S�>��J�G�cb��V���qT�P���|�`��"�%C�2{�d~c���'O�p>���\嫴�UE�����QI(�M�?�n�ɢ'���WV0O���S�c9	7�%���=��/n��̒��b�;��qrw/��Ö�3x�N�ñ8@�F�?H����T��F[�n�FW_w�v�]:${���Ku���'��8�dc�+��5�9h�w���e5BeUF>[�zS�������Um�0��/��n)6D��>��k�M��݅����r@���ʕ ��\ȠNj,q�Hś&���NU���W��RP�hǶ�{��6ez}�?��gC1���X��	���:~���"reI�K��(⒒��X�řъCZ����&�\Y8:^���9�8O�K���Ki�##�^�7��1��۰�Za�p��`9f�%dx�_�9��%��BP�@-��fZ�7��::ư���[H��>��gz�70z�Uk�:k;ɨ��۝�>�˿�u���1�fD3[�v8�ǋ�}����6�=M�|T
(���/���(M���E?p�{C��azQ����I��iM7+�i�c��/S�������~�:"��=ӋXl>RA��K+O�b-]�� �j�l�=Zl����b��n(`�	�1��t��ߧ蔘�����ﺯ�<I����-���U:�I�]KX+��ǿ�6��PA'���r�Ҡ1�a�����Y�O|v};-\~8�!c�1�,�U<�5�
۷	H3V�D��+����!!�&3`���ww��7ǭ)�%�zeN}���{���9�(��� �	��O.]-�9䖔�z���gg����/�QH��a]ӑH��a{�:�Oָjz�/ZS��5���D/ϣ��ͣ��"�p��PI�G�5��[����8�*x=�%f�:�Ъ�_sT n�!�Js��e�O��Ki�IJ&V�<��w4��m����^���7��N��"�d�m�����V___�2�塈V�$D"zK�xN��ꎳRk-[z��y�ԟ�ȁ1�=4�K|$�����.웳������W<�Ս�	���i�^��ؚNδ�aEV�ơ��6��u�#�\���T�d�S����BBB�#�x�S7����Z�Ѽ�f͞ �$7B�.���Y0k�a�������bm��rB����@�.4��h�=�/�?��k,�V;H@���U�����
�7�N���ro%��%oX��Ic"7�_��%�}s_
wLY_n'�ޘ���w�*����"��|��*lw6�����K2�s��$V�^g���{z�#��UtvN��a�����JN�I���'�<��rf���.Q{{��
��&<�W9��9kl�]K��@�|�MM����h,��Z����*�:!-��T:�]�^�����S:[u����%Pe��b_}-,Z*yV]!lnX�|�aC¸C��N3���u��89>�c�G��D�4A�Ͻ���YV�GSk�D�2Wq�3�֥���W�/�QGH8Ͻ)ؙ̧ۢ�A9�#��j��+�s��::�p33G�i��G4�S�,��|��qMбw�V��=ƍ������}�FshfGo�x�8ϣh����ll���
�k1+�8$���Q�w��B���!��� �D�H��y�}i�����������g�bn��I��dHg�G_���XEE��s]%8��C����*�:�ЦJ����K76�o�ݗ��qt|v0��E;rK��As�������X�õ�4�tpQ�\��H�2 _�8���ks�gr0���u��˛:���O�}� �Ǉ�h;�_��*&�|/r�?x��J��f�[�H�-�����]��J�s�9-ͪ��x�~aq�+�U�j*�ң�,H��Y�o�H��|��d�R /K��C��53��x�P�y�h�Ac\i��� 2GԹGp����G�ʺ��-�O8 ��h5�FFF"k%)��:& ��=�m�4�z��ٵ/���K�����w	8??*y�5g�d�6�@!�?ܒ`��a�¢������{k�r)B#|m���T��G>`���������X3��'~�͂�o½���I���lg��2h%��g�9J.zm%'�ĉ�.��A8G��ڿ,~��Ȋ�iMի�{̕s�^^��(�e]b���l؊�-l�M���q�ϟ?��<�Uxg�Bpǋe >�gr��O���cn�ݬ�Y���_����+~��<6ovg���}���y�`g�j�D�j2�Q�x�NN]�y��uZ,NAu���x��\ʎ7y��$(���L4.n���邺+̵l\��)���&��.b�D��p��W/,�I�
B�}b�e�˯��87�!7r>?7�K7i��dC>���鎙aE��_����q�!�]�a�֌��J��̜�_R
�k���]Jqn^e�q�ew�k�;��9��]�5�3p��a�%��ݐ�:^�s��꧖0���e�g�4:�afJ��.��^�0\k^�H�l�h3�H7�����y6h�y��6�m�6�����i��r�VGK褉bY��7�ꧣ�|��u.Bp?��	�~�m���<F���;L*!�$h�Wa�.BLXz<PS�)���|-o�R��OM�U����l�[	�<`c�J�}�~%=:�I���			�#�:#!�>ZP���Uڨ^���Y��=�#:d�9�~|��5�d��M�et�N/�|���spp���?T���bJ̼9�.Ƈ@�'������T%C����Iߏ��xg��7����Q)7X>_^����}��mKqv�߫]�e�+���-�m�ܪ�u��	|쩒�ߠ;=2�#�ڀUڇaT���at-S�IQ/&k]k���t���5�~߱)�OS?��������v���4c/B{�͝<'��ͷ��͙�q����Y��,�@��7��+��iZ�A�$m�����$��}.��(����4���ƎWYEE�o�@�A(��#%b�hl����\�����h?z�P����ߝab���B�br����G�h:yrN���"��r>��
L��s)�%3�]2�l�#q��[��7��u�C@
-a+2{�7�oF��F�T7[�(�J�*���^�D��&��w�[���98����F:7��'e�p�ʱ�Ҫ/�N|��&ʄ��$�Je�9�a%����|W~��%C4��j���Ŏ��,��}p�
��I�7�n���˜�G@�y��l� ��<��ߚ;����
昲M�^ڡϯWX�ήP�����e1m!�Bl¶?>����_ΰw����[M��5��#�qy�븷r\bY�t(�E6��}��Kh��tb�Cܼ�l�T�Q�S�l=E]ϽK�#Cv@�غ�վ�-ed�-wPy�)�\3{�l�C����	��������~ۚ��AGl����,�B�_oh�i�Mr�&+:���=9s++q��p_ޕ�>v��~rZv�&��Wܲ��'&&�k:z�5�[�f��v�������k\�9pYݑ)3�b.	Z2z�H�ol?
�8��M�9&�d�R-/E"�/�,�;1eB}���b����7����$�2֧ty�����^dY�Yo�_:�W5��XA�:*�|����T�M�V���i�%�1��H��&�AP_������ijxA��wG\�?0lns%>�N�H�G���^��X��چѓ|�T�H>�x�}�(��4߷�tX���F:U��=���X;���J"���?���qЉw���p�[<��o~!�n���+C~��t��ҟ�� =o���U騕�ö6�v=cc�5� U���ls"l��h��"1LK�)$�`��g���lGw��v0W��g�xP�4l�B�l�Z6��1�5���`��u���l�����|�yT�p�|&hZ�K����}���,�7�����m��$��A�<*o�8��P�N���L���y�_N�W�.�	pq�w�[ɾ��ҽ��u.��������ۯ�ڑ�V�����fsK7����و�s���+�[���5��|w+�Ȯ��0j5@�Mf��)����9�Q�<&M�D?>�-�'���{@Rb�	\s�ɺ0�ģC�c���	�R�A�o!.*د||�a��k&�F�������]�� %L�E ��˅��;�{q:�/~{�������Q\G �>�|��v�=9y�[�2c4mH!g^"�Z��y��q{?�1����R���}���o饒�0S ����?�97�g|j��0 �)6�PY���A0x�J��1�P��{=3s�^��Q�s�[b|�����7ox&ȼE.
Ժ�tB)"���m,rѯ])t�!	Pk;���o*��8���CCl<��"�r���,�tb�%�����ښ�QYU6�+�\��f��\J�pAh B�m�Ep�+3Ff���ww8���U6�@Q�x�&EF�)�+E���ս����b�o#Y��:�E �F!Gz���[��3��{����'U����;�Ahww���>o:F � r�5�A�JFK��X"h�6����Kl2-� �˛R�{w��T���ܦ4��pO�1k�SZ�y@[��
�6C���@�|�څ��ì
�����߫9�/P���/�GF�C���EFs1ՙ�����e�nvuuM�����9�#mc�����4�|	0�$��W��~�p�t+�;���.�cq �uʒ��r���6�^h**�hBSL�'g��ɦ�_*������4oTx6Z�Լ�~t�Ձ��1b���d�W�s'�ܪW�)r�렚̱4|(��m I0���zҠp
�oB����d�a0q�����}1�ۋ�����=	�,�S�Ճ���G�c��"h����M'���?k]{��E�T�۹>�Q�Or~�薔�e������� 7��"7��bȂ'���f@��k�e��p���DT�c��y����鮾���Uz��=\ ۄgqT�W"g��".֏�B2!L�@/e�)(R�n2�B��y�j���������,禧U>f�mx�ż�G����?7]e@�)�ߏ�"��r�'ռ�p�b���H:u09�'�Q�/�ң�m斘����+Ę�:'�~����k\���"G8)x7δ��k��r2R�*ҡ��2�?K[��byӯ0T2����pαC��<�&���H]EX�� ��Q j��N�ڨ���T���Ϸ7�ﵵ�Z+uP�`"��-�����M��t��U8<��c���ښ�w��1	�#2��u������?�F���!$@k�Oy�#��v�c�h�ƍ�����fR��Aǎ�}	���SvG����V?�X>L�,�����<Ah?ޖj6`�7�8[9��ǯ�%`|�vƀ��{�`$^5�����H��p*"�j����M��9����b�Ҵ������q۴%_9���P���*�"� �;^ai`l��xx:<��KK�LD<�h��%ݽ�˖DA9�en�G�@^R�F�T�ik�>���;�O�eX8ER0�fM��JR�k@9qD���1{Æ���2�5���?��yu��p���zW]X�x 3l#Z����#�[N�����`S	�;=
��H�#�dqVI�e��09G�,�/�r���k��Ɲ��ό�9�Zێ񘔣�u<���g.�J<4ֵ4kJM��a����6��V�trN�HJ�?}�pp�|?���E_�T�H�'��F� =^_���LMM��z�����K�6W0�����iK��/�
�)dF?_q@�|�*27k���E{��5*z���c!5*�e�͜hR�Q��,[{��ϸ���I�#:�<�)�0�I�����d���?C;(!}�H�SzZ�t)��w�����n&�=>���n�G��b�,����Mh�`h�O���x�"�[Y&t��[�����U���WJj�
���؀	a�(e�Y"H�`��)͉����iM�W�G�Q��ʓ�_#� Q�{DnsQ s��ډ�''%e���Y�qRL{��U?��L��E18YY�d�.����Q���Ãs0gՈ{�S�ޙ~<��~��O&V��w�Oz%???���P����h�Jr��O��� Gb`�"FJ"��8��0�9���U$Z'xh������W���<��Khk[��G;�J��I�Y��׀s]�s��~�֝�{�щ׏+�a�LJ�Vz'���u-�*{�6��a R�lڅ��ׁЏ��m��sp�����IM'�o)z�(!�����rS_�/�/�Zk@uoJ�uo��l���F��	\���lw^X��(Y���	���i�m����Yt�@��ˏ�1E�MU7����ͧ���i�=ĂIS��n[���iσ�F��Zzd՛&m��Uo@��n7���6��q���h-����������$%��e������(���o�#{�a�LT����%$��3ٗ���uE�q+����y�����[6� �5�S6-?�#��N�N�FFF��rH�:�tb}�qꖽ��2��ξN���$̮��y��F2N^�\L�2҄֫����S�Eykˀ�q�{�7vW��u��6���G7�yyuk��M�҉w��痋�>i�;��"0���pң@��4�ouu�����oS��m�ngg�},L���k0ZI19�/]7�E>�}h��h@��ÀHn��x���8���;�Z��[�7��拾�A�p
G��x9��7@�m)�O��aV�ƭԍ���\Gɦ�22�f�M�AL_ƢP�y	P�&���@�I]Z��@��1�O��mti��]�V_7����� �7��b�q�C�M1�[�5��.�(&=p�0)aȕx_H\��(u[ ����0�MO����49�I/�[Z�줻���Wۉޮ�?����o���3�6�^�|F@��%Ի�������Ζ����	�sg�1�pr~�F� ����箮�Q�>��h~�:�z�^��
�m�DX)7#�,�/��;^e?Z���p�C��,��g�G��'�ɇ��o�fӮ����[U���Y7�@:"�J%��[��y�4�JV�ݣ���a�I�M�������(z��Ǐonv��\���ꍰ�m�4��u�ro��~n��s>��lTxlL���iQ��5����R;�V��녺��Uܬwl��8"LtҖnz��~�3��P�2�nL|מ��F�X92��|�`c�5�����y�/�0��wKG�fB;d�;`dݠ�����0l[�D�9�Q�NЭX���b�oT��^RR�B�ɠ?W���{��?��;�F%��^|��x����J��a��-�Q
����ȋ��-�)��oc^~���zo�Kt����%r?[�J��A��:���k�!�[�G��]N���,C�ӵ��&�O��.M�N�L�Ǚ���y�!�������z�*	���~n+�]��_J�~�wX�߰��\�0�L��kp��Β��q�b��MX�c[�?�l��环�髴44L�C�-�@-������
@B����W�����ă��{9���}@�T�L�_��fh��芿hV�M}Eٱ%����D������O?s^$�9l����J?�4�N����o��KBL{��k���*?#��\���~���R|L�^����{�?g����ׯ_1?zz+;$��#Yq/�^���߿���j�T�+�ܷ0�o��_s��^�$"4�@����|N3���y�^������q�r�9~F19�>���N�ؾ@ګ-S7�]=�Zd���R<��= ��$�JI�����R����b��"���L2N8�~�lJ9�.V��a񉮶8TO�SG�%����8/1B�t���1����jU�7�bV/��q�r��پ�kZ����аR����u���80b�&?~��~Ex����Cd�r4�Q8�zZ���h��N�k�%n�R=��q<�/S��$�~af��`x%7�����&�0�|�2�&z�@��=�h,f���B�N>�����F��f1xؓ���c��MX5L��~��a�쵖�r��>�uP�|�p��đ��?�F���&M���Ԁ�ո�'I�_���8
}�T�Y�}}Md^��>�\C����Ι��ݗ�(,��=ϫ�~�"*߉<xr����c}��5�������1�~��6�1M�����s;�!��o~!�wBv��8���4N�Ԇ%��=@�uP�[��Q5���N9%N����9��\X\�����1�Y�V�'���t���F�OBz�gP��k�AE��E�$�?�K6&d�+�._2�Ӎa�c'�8���։��R��?�}�h�i?�v�3��跳�=�w���3+��=�	�؋iKW&E�Z��8�3��)���4oW�h��:���zg�k�e� )Rw�t�;����AZ�L셇ICl�ư��n�e�d��2�P~�je+7M���w��Ҁ�?�XE���
��fV�Υ�?� u���8�4A��g{�S���!r��V��)����
���j�]��c��\����ALJ_(�q�B"�<���8I�S�D��	sQ���[�^]��=�2Ģ,����I8��C!�n%��i��xt�qQ�ǡ��dU�)G�hR�{6pGPC#���O��\�?H�"���eH$�~&�)�i>3����'*�˂�����ᆝ�vz�a��/��^@Yl�����_}�GX��D���#�л���>��k�O���r��-�A�h$2�[��8������Xeg�9�yۨɇL�?�S�ޒ0�Α-���:_�,�> �s�CbE�fb�CP���[�,���3�.�I��T&���:��Y�0���j�Fc#��QwA�pC�BK����%�����+g�&��L�P���O���G�۰�Oe֐���h�WUQ���J��ҹ����I���v8����RRRƨ;N"M�_]�d �1W����l����
)���$�)��bDF�dT�c��M�G�HnR�
M�)���K��YW���V����}	1��mQt��2o�.NwYz�6K�E�0�]��׌����\���āz�TH{ﮍM/�,��b���F����PN]=��)���
;�4
�f�B�Ȏ�g���"��&�k�􄓮��yޘ�3ov3S0C�.�Z��Xu:yte<
1�}^n-�ʸG�d��T�a�Rm����'�ƾ�>JY���A��:�]�Ã��ģ�<#�U��fߙd`��D��߁�:������j33�_i�S���b��R� ���v�nܦ	ӕ���Ȱ��׿AuJ���O���C��5�t�g� �S��a������A+����n����Z0���1���q�a��ͯ_�m�¯m_h!jZy���h��>�v�Z���{S ���H������{���������h+�A"]j�����5����A����D_�Q�&WX�#|�y���e�)�?=9V`xxs�V�{%�YTL�9A�J�j�T���Щt���&�gU`0�6"ufK��y�-z�a�����W3����,,TŇ������h�ʐ4�9��E�)��,�T�$�A����(̈́Uf����&Ok0�܄ʼD������0\�ၡppF%�mn�����%ɉ���X�B־;N}���Ӊ�S<]������d��ZV2<L��NmI�@����^�'����Dܺ��u�	�)L8�'׭0$�@�^���}h�yTA�bA�5�c�U[
;qa��>3������:����Jz����ſ�f�%</e��ޭ�[�-N?9�t���7��FWN�v7L�%|������p��kɨ~�gϩkx!"��H���$V�ۅ��8��ʊ����4ܔ (��)�:��!n*M�	<*L}����l�,�Q&mb߽{�%!@��;�����,1���iv�l⿰HFݢ������
)����T�A�7Y7�ipΰ�.����!C�D1�Гk=v$k#�@z:@����s��E���PSni��*�I�d�"�_b����NH k�~p�����0J��:`0N�C�T
�����o�T<���/õ����É*�^_����aP�I$9��X�_ːUL�7���2 Rjjj���ޤ�$pe*�h��P#9����l�xk�>�FP��c�@�X�������)E�֎P� &�����<#+�ɕ�,�#�K�P'�c��a�_��������0�Bѽ~}}}ɪg�Z��V1o�7[[�b�%0�I�?�xhn��&������Im�`5@��P)spkO�	���?W�n.t�����hkLҷ��Jh޼�O���l�!��5/�6`��"d�\�Ŋ�"Ѯ@e��I�*��0W[�4!9���7d8��g]�Z� �2j�K�܂B"l%2T��A �o�y�
��W���j�P�V��MĎ<��"�p!��{��wT��p�C��Li=z�ͯ�ŕX4cQᦎ��L}��	pW4��*aCP�|��\�R!�Y?�����,Es��Ǟ�BO�Q7Pa��R�^�Oc+++�ѯ�b���g|��FZ�c3@�Mi��� ����z����&)���b�	��K��T������R�j�"~"���罃��������o�ңa.�XڻK�e.5�Eύ�B4H�����W�Y�1m'G��Ɉ�(+����]	�������A�鋸�Wd��}�l�N�|h�t�L���������;n؏�C�����J��Q
�*jj����v�!G��n�@L�����D����o�;���l�w�����������$矇8*vO_��g�M�7ȕ�s{h���B�*�Q,m`��s:��	$�͑�u���?��I��K�	&�����������N�P�@��P�Hl����ױ����6��5�k0P�/w���h��F��L"}���KB� "Yi��j�<��eAn��d?�A���d���	Pnؠ#֬��od=�1�B�����4��հ�Ka��a���	��ޛ&}���>�y�B�3i3H�Zh	n�M��o��%�ݿ{�h��RC[{���(u���cS�_���[�6�fՌ���;�6�Ҳ���,@��!�LiP�F��=�g �eR��6U]V�"*	�'uDU7�"7����"����Q;��q4��eF�����$�%H����Vҙ�"�l�Cf������Q ^+y�iw�>&;[ZZ���8�#YY��4��h.7����$�K�
��o���:zv�c�������v��%@�R��D*�Hc')��jkm��\V��d�iDu��p�jz�6 UA�S�L�	�d�������@#U��U Dz`�jA�34��J��KO߃8}�Œ��u��,:=1C6�@J�����S��	�y����ۇ_gf���zsN��y�['������ȉA���y��V�˴JPmm�KA>�,F��}���u�7�2ϣ�7��e��g ˌ�UIr����ך4�6��ԁ�Ӳ�M=*KoÇ0�	��`�8o����93���f�Px��P@�fᰊ����az�t�p����NpmW3�y�^%O,��I��cvcU��5�����d�J��]b^�[� z�Q1ۻS�;LZԘ��=�~���F�6^`�U�o�h���Ei��p�V�u�����x�!	�|�!��f��3O*��?��WT$�-�/"%������T#���)���X:T����c�+�ʣ᫪�Y�ձU� ���
)*	
W!�ydcgvVS�dEh�����c#	n-�M��9���.U�O�^ ^��e;�N�ڂ�ː6�� ү���V���!vs�r�aTGx�+c�=���ʬC���ݻw)�~ P7S�
ȗg��'w��
�|�#Ľ����m�� k�WىP� `Fԁ^�zk3���BJ�?�"�L�4�׎�Z��F�񭐿YSB;7߽=��@ZB��*�ъӲv7��ұa���� k��GW��5p���C�L����us��|`��k��j6p��Y�Q�����eƦud�ǔ�a � �J���{^�"����rk��K��<�:����r7���E���2;�X'���B���gV��w��7F݄�2@ �e�c'N�5Yg���f<�(��]�?���{؊�0 s"�f�K&�．DҞ��q/��$�_)���!A	Җ�Ux���]��3�-,,��C��˻RO��&9TaE�"̽eB=~��>����wi�?�&8������6����D�l3J�87Pz�4r���R����J�\l��?�&�| <*s�5���
|�G���p$7|!#�!|��˗k(�B�tگ���
ܽ�V��5���юX#�o���t&�Ҭx�}�6��"�P�D��>u�o`�%�P�xڡ"3��i��t�ߗ�ߛTd`�1G�2���
��/N�1�wi�=@��2��[��vgy\oD�j7+�-r���O���{c��̰�(w^�nB���"����z���wҖ:��|��
EYLǶwR�m{�/sd���=��S��ӧ`��0(�u=K/�k}��9�i��Ä���,�k�Q��.3�X�<�F�b��5��Bh��3h* /aҪ;��{�X����*�� �q�N�� i
0}Ǭ�{P�p�׊���k�^s$w��5��BC;ZZ�,��^��ajv�T����@��T��mwm��6��
@��U�(DK`OO����ӟ�0p�	��M�\�>l���+�s[�/��8���)��x����������
��b��R�k
d�K�%��C@X�����wwUH@���W*M5�s5�vs����kD5i��M�aQ�᭙ ��3�d2<���n|�B��\!�肿�[��z��ˮ����-Zy�����K�wp��������=���������)� U0�/�/ y�|�`:;n�nX���qU ��<hO~��9W��o��M��%���o���X=�@��������w��EU㹵�����l�(�]�G���sp��h�aK��*m�yܗ�H����"Y��-M��y%�\A��J�
{ޙ�Gw~�TT\����㡤�Lٯy��:rϵ���nacå!�����*���/�[!R=(ӕ@γ�	�c�Td�0\�uo��&*)�}@vh�����8��� ���J%4i��Ѣ#&Ϡ���ⱶ���Ťk,��b�\T��\Uݯ"��RzguoIy����Ѫz�Nv�9�(��V��.��v��-���.)(�?�%�W&1�9l���ێ�tYUQU�����n��4Z,.�ĕ}�<񎞟�~�Aqb/	���@ݵ�����'��!��K7d 2S�x������3a��g-d�%n몍�����=h"��u �6
��Io��ә�>���gk����@,ŧiFs�Q�]�38c� �Sh9f0�xtU!hߙj�.}�1�bP����l���j@����3�ۋ}Ċ�F5⎞�Q�$�n��=E����vKc���N���Y�S���@��೘.%U��*��
'�w`pVtb}�c}Bg_��,1ȁ^jw����r�1�5l��ָ�����	�PT*j�������/$PN���)e��3Z�=�O��Y���5<�^l�ȧ����?΅��0�gψr!�����7._�����Q7O���K��L��g*�}z�}vS�̓7J4��oM���QS��P7�HSS�!s�E8�{�1�K����_I��%�LE��!�j~���JJ����6H��j���dX������94��M�'�z�sN"��=7h��Ӟc�j��*��? 4]^^V�Z�����������������a�w:9$ ��H���ď8�S�`t�Ϡ�AݫR���&� ��z�$(c%������?����bׯ�u! �
�zƻ>Uѐ�o���� ;��4io��u���rm��L����۾� ������������0���L�%����xp�zV��Wl�����lm1�Z���'�:	���Gr�\��&�@9��Ĺ"�����
'���O�y
�pT_+mG^����~��3�d���J�z�$W"t�,������Q�ͼ�_S|8��sp���VIÁ�.�FpW�I1�΍7�{���z���F���P��m��TUU[�Zִs'xj�Ҽ،|�{��2P� s�����p&�1+�_+5?G:��߿W�;�>N��u��k�N��뭅�8�M��a�n�W��g;�]�_]�/+-%Gm ���i�1�sNZ� �?�9���$^"n�»*���̇@��F�F���H��Ƹ63]j�df%�y�'M`HW����B�7a|'�!�#�fl)��uw}��E�ϠʲהPSԈ�u��G�#��M_cjjj��_.�i>��Yd�*�����@�Q��I�� q+eB�j\�K�4M������o�g*��X�8y_�.|���0#v��g�KgF3��)�0��d����:lH���b��$!��i����z%�����+�ߝx�l�v�l����������ޒ�hx	����fy�<��+9~ ܜo9ݨ~o+Fda	gv��w3��.,�iװa%������{�p���xZ�)���HBY�,-��!�!K���(�=!�p!iȖ})�d;c��������}��z�{�����\g�8�j�|��~���k�?��0��3ݞ���:M�c1�ͪ�W�5U�`s�\'���Ó��� �L���N`V�Q��x�׿�93|'��,9��n�*@+���	���A��#��拞��FY�y����UȺ$%�Nf���>_{:�A���ؒ[�LBD�p�Z���ԝ�ԗސi�E�ۨm�)(�*qJb����IY'96�Ho��I���*�%U��U�WN�x�ϊ�~����L�^����[���,a?7������׆���}	%��9U��̬)�I+]��gzz:� ?C��+���vI[�A�_3��uzG��e����؟Ir!߃�/?����)K����e\sI�7�77]--��g��5s��pQ/?͆�՗���m�����>$�thg�˃���x��h��ǩ��������o�(/���m�m{���;Ix��֫]��!����?o����F.Kp骈5�[�cx/\�6#�^`���񫛟>���R���O�v,�
d	7+�=�Ƨ_�XL��P�Y��v�����	ξ�Q�=��͉B�q���מ��ݲa^	2j�ǉbT��f�tP����5S{���e�y�@���Q�]��}̸�{_]��y���n���'����|����'w<��c{u�yx�iYD_���***FS�0E�����ֻ�+ٌ��8I��ғ<��}�c><�7_"��%3d&=��t�"Ҏ�Z:lǒ���ʤ���%x�|�Bt�gwh=�h��v�i�Sj�n �E��]]U����I��f��>9�<OL�V���o=8� �]׺��>������Y������F�����J**�E�%YY�&''?�_�v��Bbu��=��¿�<���/_�������4�T�ͭBۛ���-Ky-w������u�M�eq���KmD=�>:��:�O�|f{Mi{ˎ8	L���wz|�|�1�h�$o
�N����k<ZW�8�����x�k���tͤ��"��x�O$%��)��/�\?T����<�ȝ@6H�̗�~���h��i�g�K��r
W�'� 
�Q�� uhl��@��w}mޣ�J:~�����~����$��%>j�䉎����y�P! [������K�OҮ[�tq't��z�������=d���}�0>����fj����A��B�z#a�ħ��3T�8�������M���%	$��yo��M�Ŭ��
��>�ΰ���{�(��i,��~bD �J�Vɢ/\�1�{7�S(E�f��q��H��M��W��Ǔ�EX�$��p5x�-�/�(�ο�hO�N"��|Q�/�.3в��Y-��ć��i�x6wS�j�.�7	���~¿���:�$�@�'DLd���q���x����V�����kegOz?�]�5����Pk�$O綳��b�[�N_�}�,��%(S�4�����I�������Uފ�92_�l3Ց_T����u����OO"�L#�b/j�512�z��0�iN'8�2�dO�tR�ߨu��N`���;^ �4+#E8��ą--9�ܽ۝E�hK�_kQ"E��#��Ρ������KR�V��d�g��� ���޿�cs}�ky��/v�b*bL�W�׎�����ʸ9:YwnS�*/z"�~5��u���^��Z�բ\`����-������<K�oPZߌ�jN�ˋ��R&����UPo9�ӽD���G�s-�$��_;�C�����E�p��2eh����`�We��x���L���h�5��pV��e�CI��d���'_�.*�Y�Ծ_������I롣�܋��/$��kdX,J�=�5��/boE�г�"�<�ku�Rb4�׬O���O�ꘋٔ�̵oB<���d�vp�3ag��}r�g�H�:::��U�� �y�+�b�3z�?BO�ٷ6 ���������ϯ�z�'Z�u�mc|�ܕ�N��xX�fq0��Ys|Ul���������rs�r���{(�)��\_h�ِ(�8�K��$��cy �&�-�cN\��ٳ�s���z�	גw�Ђ�*|a[�J͝�<]�.2�����|�un��c���v��U���^���z���w��+��$_�������l#��޹s�Ϳ�(�G]]c�2u�g�ڣ,<��BG�u���寖��*�/�a�a�puO�z���.f��Ƒ�m�'�ђ3�#&P�/���G�-[��B{���O`��!�/�=r	�
`)^��xf�/@+aX0`�.�z1º�Ƥ����f�lIX���GF`->���a�OB?9��� i
۽�~d�}s�`���<nɘc���g}&��@��(��b��O�����ώ|�౔n8���\����m�.,<�h�z�)C�=�:�<��E���D�|��مcm�Ш@92��A)�&�R?��ֺ�|"TJc��`V�⾄��6mÈ@&���Q�����-���ڔ(� D����-����G(�ǓJj\��Ɯ��٬Ah�"�?����.Nz]����W��'�����$��gP���>��+���gQ*%��t_�k�;�Z��\}f﹯�d�����2ɟś�e�����	+��+s�5���	�U�|� �p�ٟ8,YP]��i`sw7���u-��to^.LMI	���l����������P�'|i ��;�?h��o_���㗖��p./o���'̩<�'�6��굍]:.-,!�h}��6g̘���A����ui�Yqb��e1l��;����.�9�������n��?�^�����GW�Ǩ�3�;������R\�L�-�X�.���?��Z�~�#K����
+�w�5A�[���s�b�ѹ������e�TF���Cs�C-��'�F�[E����Ҳ��_}W���ằ:j��*��i�[�Ť�%���|����6=���sd2a�kJ2�u	��(¶rIE)%�=>�;��O��]i���]����׺Ҵs�����m��	O.Υ�z~/Ӡ��SYr�u.�?����9�suN{{UH���G�{y��M�̀3t�^]�/g-�o�9Ñ��h�[�9x�B+�¥>��J[�ku��u����˨q�l�
����oѭ龖$�|���M.NE�)A��\k�՜u]]��R�#��Nt�H���ȸ2?[IW��]3X$||�CD�e��lO��C�y�IE��@{�7a���'t��)�#���*T�#bԟ� 'q_�v
�R���o�p(�#��R"�u?G+��gt��'P�����o�n9��w.�bB��,����?ݵP(n��W����];\E����UOv�=�jL�ŝ5�W�����E�)�M;x/�_���Oy�D�7�W˰f`��y�:\�O:|pw� �s��L~�Z�y�"f$����<~����θ/Oɟ� �{��^wR&��&n�1�g��DQ��?އ8�%�����w��R4����_���0ʄ�N�q��<P?��C7*B�La��]&�7���Z��=��3+ncD�+�2/~��C�����p�7�+�V����}}^Fa�j*t�� ̬����&!�2X�B��G;��q/�U������\ƃ��ˉ�K����ɶ�3�2���a��ʈ��<DU�M��.xn���9I�����i��)
�vگ���k���v�d�{E�%3n��E����%��JJ<>�Z�c��սI8*�s��{� �~Ww2E�B�\^���i'Y�\��L�k��6ٞ�J��g�S�<�۽�z��f �BR�?n=X��dX򈡦%I.��:U=P��@���2д���9�%�C��D�ob$P�$W��q&x���a��rDM���{O��i��y4��r���6���P|s+]l � Ag�ROptvt�z�$w rE��pɥ�ta���%&��bg�?L<ѣ$츢ᕨ���0�R掁������~��ؚ��ռ�o��ٯ�̕���ޒS>�������dB]��h�������t7��Ç7;y��{�i�f+v��w.lxstik����öy����Hx�����Z������Ǐ��1 �y���V�;����8��~!B!��Z�i�X��7,�tO�ۮC������r��Z��2Ȩm?�����r�ps�Lވ�8Y�x{��hG]�D�@����|�'�
���9�955դ9^���c���KRRR3���gb'��[<w�D^_����ZO�o�;n{9I�}0D��D���������M�_lV���u�G�} ;N�&0z���}Λ�+�_hؕ������Epy�F���N��O��8-� I��K�$��ꪫ��w?=��?�����`�pn��kg���ov�k$?�V���?�סП�aE�]�r��ٚ�9-�� �XFg�3Ort��Fdd�l����aFY+��a��JO��{�,�˟<Y
� U��mDք���_��]f�Q;�ɰ�qaO���66(��z��F1G�0#P�Q�9b�79��!$*)+Slm��p�w_��^W�IF��OO��]�|�q_6x�6�L�)잷_�^��U���Pb�|wkZ�O�ٞTztwO#��+���_oy^��L��b��f`]��zo�V
���Fi����d��aP��TjwЉ�2�L�>Q���������C��MV���eB�v%N�"x�槮`�6��Q�51�!��Qg9���m��AQu�y��u�Ľ�ս`��m��P��q��:���0à�'N�˩|k���p�.Nڋ��C��[g��:�mٗ�q*���P�A멮3��F�^km>�2^�6ִ����;�]��bzۉ���wV���o��)V�1�)P|�A:�Yo)/�o�C��U��kP�S��{K�?��~O3gK�pZi[����&ҁֽ��h�%y�޽�������>�|kk��H��?�3�㛶��A�x�{��N�������?��Ν�*]p���:?y��7�:������ֳ�ޗ��?�D��/�[k���w��># ؑehy!�O?�җN1���y[�U��"��2�Y�X��r�|H��{��M�A�|r����d~i�B�]JQ̸�%����b��m��Z���.�X�e,^a^�Ҙy{���O�Y��/Dh��*JN/8=����+�Z�频�9o�����:E� �mF�/=�����~հ�bA�䞧��L����J���]f�q̕�֗�'4�By���n��m�~?�Wj�oM(cE�*����x���A����5��[i�O����1c����ʭ�Q��1�a�v��i��4���p�aS.��÷��ټ B�)��(��ǔ��nJv	ey'�6W�6WT�7{�	�FFLߙ����� ��ļ�:~�k��B������m+3�DOB����e$%�#�%R�w`^��8>/����2?TwWJ+�՟S���SVn.c��0� z6��݌���c� =N&^���Չ�(��!�3/�5�ׁ�>i������O�ś3��6xeԪ����'������ޘ. U����**��0�-y�,ll1^O"L�z����\.��n������ ���1p�̬,���(�?,�t!���\�LiZ�[iA<$ac1U���MS���:NKp}7��re���t᧼��0��ʊKJc�G%��� X�̒��Nk�+��,#�d���l^C7��(M��a"���̐fa��}x���C�1/�wuɕ��@���%�TR&�ccc�r(V)4~I��rs��ByS�24i�bG\r�s�4�9*EW��)�/v&��ǌ6'Դ���3 �H�N�)	28j^Dy��e?V�ɾf���VZ�0ڔ��_Y_h6+j\�pMY1&�	l���aaL���t&�}r���hPRRw���rg"� :� ���m���1#i�7йϕ�J\��K����B9�e蝉}�I!�w��n��r��˗g��4���,����W�ǔfӋ��aU�	^'��$��݄�y���K��%�*��(&�0�����/|��."���̥��7~��zT���V�i��v����L�b�?h&E�Tʏ60i�{�������$�w[KK�9Ȗ|�{�)�����:���x,�-�L�x�:pA}%q������6����1�1񥘖w)����O�u/�!�����"�pUrp�
x�ƨ���?���v[e+'�S�̏���D�c7C�:�?���w+�Z_d�tނ�	���*�}q�һ���>5�ʖWVƆ]K�Z4Iҥ|[t�xK���<�D����
n.镻N�ࣉ�W��i��V)�T	�H�du�aZ�7~Ah�9Xv}}T**�򻁕���d��@��7�4�̔�4W�c��a�׸𡻧'�<�&CMM�>h���BF��K?-]:�w6/BbV� ��qd�����"/$p���	70��:�Y�ٗB�j�:G�;��Q��0���@���7�ď�����vhH�˳�DA��|��i=�,��Y�7e-�$�'���o�^����9��쐀���;t�AN89;��O57�Y�L��x���H:��pY�mF!��ڎqQ�=�5�,�f)T��~����`蹤�1���̀��ŧ�������6�G��:�T�8%)��+���e��,�---UZ�232���f�7 �"m�ي����p.�Crs}�e�BR-5����� `F$dE�ɇ��J��ܠ@+W���J�P� ��h����<a�V��0��S1k��1GH���:� >�)��i6צm(��j���9~$ޤ���!���l���|��_�~���,��b�\l9��~�Gx7ת�N*/�����\J�d$u*��V��W �Z�]���sc-I��C����	�˜�u=(K��:��'�Rܼ�FO�b0��li0.7aR�5�\�T'�a��)�E�4������K�̞��M��l���#dE�,����Oh�DDD�\�	��1�����s�PK�yhJ��&�����ƕ��̦��� Ω������V�$2 N5�J1_��
�"�H	z?�5�zR�f����P��o�v��U.������|��$y*G���k����/]�g�M\����2�l����	G����,vc+�#E��S=��>;����_�����|X����0Na�� ��2��M�k/���_���;U�c�[ǫz���=�Z�P/�܉�ǵj�[����G?��]�����je_-~s�������	HU�L��15@���?�F��O �RȤA��f����K����̂fL�i�G]�@�Jڠ�U�Ӎ[{�@�g�K���qRk}�D���L��TR�~���2�y�??%�_�`k+����g �VC�)�	~�O=�$��L2��g�6�I��t܅��x��F���]ggg���O7�>�p~���+�Ƣ�%rxU�(B^s���8���X�cfgm-�e�ga�����Ds��q�xC,+`��A~^���Ƚ��bi�S���u@�ц�mU�Z�J��jx�ԯ9���
&|̖�0|R��0J� �e�����67i�y�Ns�r�I$�|�TH3�hⴒ����3��B|w%�|-}e,)dDd�C�X
I��v��#��Wi����к��������v{`�Y*84�8�����ec������㮏��8�_7ӹ{7�p}�)++�b҄�r~w�� ���[��R-���P]����r_��u�����j��\	�\	�
w����r����H�c�ۨ��2��JXⲃ|9~۩*����;��1_�Q�0]����pi}I���b�u_	Z�C�pnq�U#�x�C�UR��h*��@��X�&2�����B�y��?b}�6��/���/��v`
nq��>������p�\��3Q���=_�@B������@ ql08�8�i�14tl�1)���s��?��P@ZҪP��ϓԻ2��<��	?�U�$�S��u��KŮ�Q��&ǁ�4�k�ڽ���0 ����V�m��R���W㥰l�i����B8� ���d���9Z�x�m��J�ˇI'�����`���#����m�*
q_!�oe���e����7&��|,9_oN��:n �5�)/D��o6e���Q\�t;(��?�r�{�UZ���۟Q���{��zF��u�#�H��a��ؔSDf i&���$=��UW��L?Ǒ���2����+>xd�B�,PN��_.L,�iP����cR4Ji0&�@��	��/�.�e�1v-�;�V���ճ�j��o��C6כ7���	!0����
�W��#g3��E(m@C�{�������EYdS[��jL�f�D���Q:��
�0O�--m�S�/�c�����]�2�+5R/Q���4yl��J�d�)��bY��l^c3�Q�/�Bʃ ��~���=�z��w�J��N�� �rp����E���\uc�ڋ���y"
_�s��I���&d3hV�B���@_�;�a+++%�o�9�&���9�Z����q��d��ef8�Y��	�I�JW��H�58�se-���}�؝���l�J`�J`�;ɚ�Q��,�b�p ��sQ�y�����.�c-����� 2�g�&%�9/Ĕr:�Nv�a*d7��b*δ[��Vn�W�s1I�-�ׂ�qI������VGb���q��������	`;���%�0N`+�t�N��L�\W�Ҭ;innN�����RNjyX���t��
%�����VR�)? !���-� |�q��Ѻ��M�@�)�"y0)���A�IՓK���C�R�Xm>�'�)o?�����afc��|4�@D�/\���:`Y���Y�ٝV��؍���N��r��Ŕ$@]��+ ��I�_E��py�V�*/�f��s��؝F�y�R�B�ǥ���t.��)l�!@c�����B�/⿘�&�; �&� �cG_��u>3��o������O���Z� ��=�ih(A`�@����:�kU�������J$Ջ�]/�o78`�[4�K�������0)�2j�?}Az��X������3�$��LMO3o���L�]�m�
		ܠ�3����VR]\;�y�����ʀ�{x��%�t��J�2���{�{*�\�ҏ�V��Be����^��5�rv44?�n%˼�*kO*?��8H��j^(p]0-��
��>�u"�E&�Q�s+#.���&���=���i'�9i�@�]\]��@fwtu �b��Z���>�,����]��n�P1t&� �S �=X�\��H��?b�b�G��㳒�g���p�PӉ�)5���I�K�O�Ĥ�on�L3z�����M�~|����Ni��!���nyг.���u4n�߇n1���:��W��7�GHL�G����\v��a��!Prrrj�&�̯d�x�=�<Zש���#���I�D�ۜ�Gq/�j��d& =K��>]��ϒ��J:(-����/;��}�d�*��[�ϐ��l�¦0�䶦�TV�=����n��T��Ӣϟ�n%4 �lliy~�Dj��~3_���e�zX9��ұg�M�V��`�^��� M�h0�����ׯ��M
m-���D "�!
��-�s�J�8]--��6�¿Lo@�|_�z9�h�8���w���o�Mt�9d<�(������F(��	O��E2�6���=d�1L��#Z=��ׯ���	��'m��ǩ�}ț�͑�=��ߟ��'W���*�naD���~�����,ڄ�������ʂ���H:��egg��RHζ�8���)���HT��;m Ē y�/�'��Ԝm�^ȟh�  ���,�ײS����=w��q�x�F+�E�]��l�4��D?���3����@!e�����-���|zzy��'1	Y��P�����;�n��ipVSUN���l��8�>��ͳ���`��y��~�m�53�J6U���-�WŶ�ذ�V�4�� k�,5'H�\u���Fҽ>�� ��W�$���;­U�y�d
�c����p���c���Ebg<�F���v��;��G��P�@�M��P!A�HOu^w!ȿ���5Q��GKA� v�qFw��~�>�va=��4==N�|v�R�4����=��	���%�7�ίF9m�܀����L����6s�s���5Rvhs���0��s*F+FsD�e�.o��,4�����L��L����Wz����ꑑ����Vއ���Ģŏ�dT�e���{��$�Af��JE��$z��^Q�%�auxW����蠤+�;�a�z{�����m�����������ZY[W_%�����x�Z�磸ϐ��ڃ>��s��p'��|�?��߿�@E >^iD�MVN����uq9����/������6(����1�m[k��$!+��W�׋Q��L"N�fq����e��هg� ��r��]��0��]���S/)�a��7��t����h�G��A.1�@���FZZ��$pl���?�2�$�Oog�5���ww2NdT$�х��<�.�������4�i���y��t�
���v�]h�	\�y󏭅H���Y]�A�p%x0$x��#���!��6�.�xIϵ��?Ӝ� i�`
4����s�՘�qO��@�Ij�?���MQ��ޗ5:���K|�d�7�$kYHV�t�q�7 tP
*wz&��J���}]�}�X���M���T�%��ѹ����)�1������I5F�E�3�/c��}�xӦO��|z�ɝ�L�����&ϘƔ�N�0��O�@�1�&Hƭ�T��) �ׅH�1��ԅvʘ@3L@@M{�ݻ§!��ff���lE2�IZ������i��_�ڊ���+�!�t<�;Ԥs%KN8��r�
Z4�n>�*��ֆ,�%����ַ]ls�y@@2jJ�sH-�@Y��E�%�����)�; �s���"7�!�;�!g�����<
�=}"�Z�G�t�Y�y݂GIݟ��o�E0��C��;::� 'cJFϖķ������=��JcO�n� �A�L?�z��n;���}چ;MtqZ� [���[S�3n.�+s���Id�F%1�eђ:����M�d�<a�0��6�	t�4�}�˖}��4�i9����� �&:*���<I��Di$���I�H��Vvtw�ұS=$�T0���u�Jz[@6o�M}ٛzPa=�ĤC�a��=k��H$���d�s��ZyTϘ�Gd�V����r5���+�~ ]�}:�/[���O�l�bY�ģ���G�X�=�e���M��JL���!j�m�����^/A�#��Y�b����A1�w�����6�6��#��q���K�"�- -��3#۲�h�%�vvc��f�9"�ǒ%y�<f�(��@�fg�T�qs�4�lb���g����1㕙�W�ܱ1^ G�����DdT�P��L�&���F��}7��=@J�%�G���4\�96Ɲ�˜y���lk/h��O�ʕ ���o��N�o333?��r(����Jz�g��T����ʣ3ʭ�r������ڊ�٥���J#Cn��y%}"#
DK����Pp�����?I��ʭv	��m��[h�Z��EcC��?5m-�N JI¯�7�ݖ�u!�4,�s�E�xt�0�R
��@�|ݥ+�&:/�� �;�d�ۊ^��%�;�j-����]����Ro��[��T(�}y"�'��t"�}��{*++A��D7��*�����%rmQ�������^k�7C�J���2a�h�H�%*$Yl��:n��M�+ze�9xm2�Ɔ�T���݅������ѥ�����B�����N'㙃���7K�SI�r��c���a_6�M��n��K�>��^]�ƿW���s��xq_q����%q�5 0D��=�?��~�q�j4��m;���(�#;��m�|�.ݽ{Wc�:�o%�?��:"d� ?2os��U�-ζL$^�S�U�
������/�f�x30�K���ޮMj�S���J�"���!�ӊ�@�z1%Cpz��r��?��p�31݄8�@���J�DZ�c�G��Vve���p:<7���[S�cCu����=�ۚA�ȣ���S�&��~V� ����7E��5��O�r񇭕�3R��Kś�������$
;�GL#~+�a"�32;+ |P}WI.ӹ�7��?0����������f8�O����(x��p�m=MTLl��M����3���?k�;We����>�i�&J�^�fT%�^�z�Y��U)I�m�x�Ʃ�ӂJ�wk|��n�3���j�^@�We�yLYn��Pw@�˰bg�ڨ�� ��� ;y��1JѨ�v�[�C��;
�/�`p+E�r
2����Z��/
§��>�#8��d�Y���SCM嘆��?�������/k
��چ�X�u�l&�c�֩e2ET\<hpp0:���<��cAΞ|.j����l����1�ʶ�ķ���ȅ�oS���Lo�x��wB<���[��D>𿆔�g�F]�uw�^�􇎴���Ȱ���8\�Ӊ_�{2��1
�o�� �&�kdD����5�:�蹹�S��9������������6�z����tH����������@n�xeR��kY�M��w�a0�.R�cHy��}��򎀇;Kb����?V�5���=9X<���2����P�:V ��}�m(����w�ɽ�r�&���J�(�du������+���:,(�P@S󘦡>�_�	H�~;�$|��pZ�)$t+ʛȼ��s~�ُ	�:���q�JHC�0�b���� ����F���*ٲ�7��o�6
si����	�|(g � ꡧ�O�g?� )N>�{�)��'<�c# ��e�MI;0�thm!���Bh����X�'�1@��2\8�L�hH���V*�w��..��	>���,�=_��owo΅��{/�}�maA�����n:\�qG&��;[�pLP�e�>���]���o�" ��=�0�J��֪a�P�o�aBQ�i��qa-l`���i|��:7U�r��O��Ĭ��BF��YRO��5�v�
�NH�%M���ځq����v��qߎ��Y�#+6jJ�r���nT��T9�%�����[Ȃ+y(**�S��V���ϟM�m���T����9m`��%Xʅ�`T���� � n���:������3 5*M�g@6C�_
��HE���.wY�<2�=n|ٰfsc�BFh_~���D]��N
LP\½m?*�033�?�8ĥ�b9QJ�+�_R��V4>^j_LK�r"��>5m����2vvv6%��>9��z �Ҵ8��7��c+�v�\�W������I@���]V��)Ny�6s�{�RV?̐���Ve�#�4?��O�٣� >2`�Hl����rϔ�����S��۽�{O�F�Y��m7v��6b�))����XJ���i�����[^/�h㴌���?�M�ފ��r���}�+�l�!D���o�3�(�h��$�|���b�8��"��3�/z���a�P�Cr��I]a��S@��8-�+�A1u/M�V����a�NyHŨ((/ר�
�-�މ	4+(,,��
ݭO��v	XO��2:�J?�~�]��/��^- �vM�n��V���7kz� Sp \�P�#��c^���Vut�����Ɇ���<;�p����˹Y�K{�?�	G_J��m�L�X��j�f����<H����4SG�A'`iS���a��ɊD�X`�Q�ݿ��C�����jc��ذ�|�Ky��9�0�9�Ey ���P�(qPuu@��/ܡ�������n:�N�~�����zi3�g{6nď�Q���D�,�QO�=�	h��V-�1��g���bH|/o�0���QW�\���=��]���JP�і�贊��&�/� $�sr�2�	܇l�i)��`�Y@�	�jD�i3��}&���C�C=���s����)M����W���`�^�E#�P�=�i
�B��r���Hd;[�C 0AƏ�8,�/�h����֣z���h}š+�($s��bl����Dp˜i�=@KK����Sz���6z�3�S�0�Pκ�m�~�[I�]��FŽl��hu~eE�E寒��g�����!��l�ν�H�/�P/�v��[`ER��$*�kF'���W�<��A�u�Ng�&�7uw��Д�E_��i-��8�cRh0Aj���1�8ф[���#�j��N�M.�����Z����sT4�.+H?{u�BlO����U��-N���1=!�������
[ѷL��BGWW�wµ�{B��Y�}ֳ��#��s4 �sG1�� ����7��14��  k�&_d˦N���^jO*�i@����=�:���+ i2O-���By]�MS%�3�+�CC֏q���,�����?M���5��X,�I�{,"��L'�㽗z��aXf$���u@?������ُ=���H��Q�����O^�:������aU�"a���O;�E�d��d�����g�A�@�!`�t�/��>��B+j)C(t&:�u^w��OQ�~'O7�S���̬/�l;�y
�=�8���TH�}b��Rk�?�P{���]E=&eV�{v���N����p�H�\�f|���	��yK�㽋o?'#�ٟ��Vn.#�(D�)"�R>T�h'���Cי=��s_o��
�ޮ�?�S�f��g��yO �lll��F�x�zS���㷇����<�#��������G��Ӥ��V u1q�ۨ� 
'�?��1vр�qp 
C�F-0��*hO����T����u�+�s�S�f3���H���P�u:u���wh�����~M}(�I=&E���V����EYd�o*$_�Ny���j.M��8!ZHdP�(�
n ����[?��u����FS�y��� ��vEP@��MĈ[�_�+?�l�o�ֳG���1�R��Q1o��o�0N�񻴱��2�����=kԏ�ɁJ��m��������!@`��+��v��o�nr���0ۆ:� �|�k���oXh�2�+�a���hG�H�du�EX�Kn�0��e�V�����S�}=_o�w�`�����z^��}��]:<
0k�;]9��s�~���`ȧ�#�����0~L�.uwnɨ��g�a����zT%�3%���G8��r���������?����Y���j�5
�?�����k���r�����;��;{�cd��Տ�[��A��][�z�}5�P�����%j
*�q���_���(�A3r�D���l��p��'t��B���w¼m�\��������ͻ"�h�+p�_��N��o���-�'(dm^d��$q���N��R�a��g�^L��ټ��n�kj���0�F|t��hwK�[�������O�6�m6�m�"D�w���z��u�:�^O�����ީ=;�矟����w���>�+�>�@	��
����B��h'��M�u������M����hgzKQ���ݘ��.h[��HXWs�_�;���(���y�ȩ�c�߹�$���ѧ�W������iJ}y??��5{�f�k��x����5�Nm�Y^l:�6Hz��x��T�c�C���uW�~s����kѺ�u�Lյ�5��0���]㏬�T���X��ŝO�ݝ����W������V��[S˶����1���9�=}O�Rc�x�͍ᚐфg[�˗/��\z_J��y�����~>k�f/��8�a�<?ߛ�^ӷSћ��;p� �9m+5��]��jt'��Y�.������e�m�R��v�֫N#Q��!�����E��nR��f���������@0����C�����=מ�o���8X���૓�5�_��5�_��5�_��o�yʏ�칆����������������x�>�{sH���C[Wk(|ˆ�gj�ѿ���# ���*��g�)4{m�����m�fd%��z9
�T�����ݢ۬�?E{��w3�)4�z?��[����Ƿ�n�y��~��:Ro�QԖ_Vqc��r�"��ջ�}�/X���sU��O�S[�}3H���L�w��uUY�!T�4��������
�O%���2*�7�=�� PK   yX�%��7 �; /   images/67e1ca3e-4bd4-4ce2-a74c-9273116ca70d.png�vUS��A'����܃�;��HpI��5��ݝ��.����?qu]3�5�0U3S��"��J�
  0��Kk  �<��?��]��� o#�,��G{5C������ ���0�^ ���i	-�̳��T�Ewz/j�ŕ2���XJ�`�/�x_�Hh5�������ަn_�@7SJ���s���H.`G�z�h�(!q\� XԆ�l"����Η+��\�������B��o���UI$��A��xj�&`&���æar��GG
���� X2d�\:��]�����A�������B��̫H�8��\>�%Ɓ;'<=�|����'x�:��������kLn�<oP����l��脤���:49�ޤ�Vm��x���(�c�t��P���M��5
Gج��Ag+�E�<o:}�,ۆ_�7o�/�<�ƥ8�&^h��L�\�+﷭1\���F�����.���d�߯n����/x�wS�Rx��[p���Q�<�:m�#�۫
�ݜP~9r��(2XA�AN��>lhզ6PSzov,3��9`o
В^9>���h�Qf�������,�����޻63���;k����so�V�)�t��O1�wλj<��<d����rH��n*p'�@xm��z�Y���Vԋ�u�(�ڿ>DM��N>iVC1��Pc��[�5�P�AL��{:���G�Ɖ/Y��4�fOjq�=�CE�f���\bo��;���w��4^��VZ�S���B���2��(T3Ԟ���8�))�ca�Mv�G�p^����Q�_�q�mS��M�#˷(��ĕ>[ށ��:p3l\sȠWA�]�#��u�����㟞��v,���6|�8@��'u��k#�S�Z�X����A�K����U�ڋ��(�����D]���Mm	�c�a�:y��%��`cKN={n�x�LQא��@��OT��Ǆ�;��*h�,�"�) �N��]�tN���(�����4V���/�)������|{� ȾԄ��*h>��I���c�k�&Kb������>_/���!jz=��i�@i��y�;n��!c��-0p�-s0>��t5h'E�85���C}k���Hx�ڸ�'�J��fmv���tY7��@OsV��&m�Y�\%�bW���b��$)��J�z��1"�rw/,�C����G��]�N�{�{�!�M| ������K�?���5[4r�78j��Z�,��>��1U>h��H�o�ܯE��V���,���*��aL�`E(*���:[W�h��v��r��$+D>��_|9o�yE�5z��r���y��u������(�����hS^w^m�S�P	o=�"����).9�K����IkƑ�*ǛR����Tm�Q���:U��4�֢�;���+.�l�p�àE�gb�E�e��Q��~����ERc��F�ԥ�����xV���ި��~���3ֹg����zU���ΰQ| '�-(���T��Q��c�3�J]��3�E�g�Jy���q��}XC����5J�o�̞0���� r�f�#��5"�`�	ݿˉmN��]Φ��1��^R}w�x����X���#^�7���:=fV��<.>C�������C�˧R���R#K��y�m��T��o�����"�lſZ�[�d|V����������C�����+A����v��X���KI���B��s�6����)����z����\l�>v��+�ֲq��1���C��C$���~}o6Y������u~H���e����n/F��	�Bl�2�uV0>A�@0H�d��M^�ɩ��͟�ˏ^j)G�P��6W�¦C0��+�"K%��S:�.ƣ.���ʽ���3��񧫬�я���6�I�_�Þ»wN���)-����-����,/*�v������.C�8�f+"���~��W�g�T��6�����Q�%X/-�QK�^J�oek���/WA�0Df�hf�-� `FZ�9e�Mdɏ�b�HHI�}s�.���گ]l��]��
��.�YM�� ����!V��gԜ�?��wP��o�s�Z~�6�J�J�ƩL(H�P��V�"�o`T`]�E����q
�+�����^j���'����o�����)}�#�����OLN
@<Go���.�w���b�.���|�I��?I�u@�MN2�qW�q�(���6/��y�Řm��7y<���`��`ʃP��1���\�3�@��,ڜ���n=��Xv�;Q�`���VI<��P\u�W�Y�=jw�RB4$��P�V=�Y?���k�VGFZbLsa�a�f�URJ='�˟팴S���%6�tX]�:<(q0@h��`h��ܚ$��-b���Lzk!�̈́�\�d������e����JV1,@��t�痢� ���?��Xe$����
�O�T3�݀֎N�$K�h�:���U�	X���,"�H����D��X����%9�����l?�s	Y�vK+N�	"��� ��ح�~�k�5�E�R�(e�Yv�E<0�����9,�F�T��(�PQx��F{��]�ލ������R�a[�����,�+2�9��8�
q�,p�k;�8ȿ;5�<y�03ߢ*���5n�t���K�"HJ������A����;"
W�P\�w9� �A���i��>4��(���msXlʶ�u����D����l]u�p��oү�m}�fg�x�^�=�wX�n$5#�ߔ��
�Y��n���XX\,���2��G�BU�8~��@��u׵ѭ����Hb���1�����s���1�N*�g����� w�l�z���P��M���ߺ�]cOLMe<�d�4L�����>>qe׊�ѧw]c�>XF�"��복���<�qr�P���pBx�mXpЅ'�ı��(�X�[N�k�k��mkT�Ę�K!�V;d5�A�����N^� I�3Z]	�,�c��1����Pэ&�=���.��М-��Ui���C����+�m��\�a�?�)N ���d�Յ�B�?�v�
�n�w-��	�zR���Y��S�5��`�A�k$�d�'�ߒ~0�G�J�_�	���3�^h����B.)GD�W�l��K߮bdZ����RA�rLh�9�@(�Bz W?v�_p�9۩o�4S�����`&Vҫ��Ȉ�GB˾�YW��WЕ�K�3֣��	FJ�9�,.�����(GD�(�/<����Rb��y�NK���}�j��2jhě!��O��T�vԍ�D/���4!�2���?Hbo\�>.�yA�L���B���n����O}>������Pu�{_f��|��T��F�ଳ��0-E�wb|�=YL�L����mBi�c � �u���$a��*�ED~�"�cCT���,�����Q��V�_��r�F�mGs�Ʊ?�ITI�mJ��}�_��Vq'�>�A<W{��,��9th�A�;� 8x�� uO�Y�Ndr�O-�/���M�Q�s��l;qf�X��_��{�t4���� l�4�����M�1׎Y�0�i%-l�ՙ���QO��<[�`������Ym�C�G+a����pb����
9����9�I��@����˺V�Y�_�Z��KXFT������eW���z �DG��X�:�� B�4�R�����N��&^T���X��������[o��a0��� �r�
�j�M����C�zK�J:���ty�����������k�nz�M�}nNm�h�/T�6���7]ܟ�K��'�uc�k�˞�7;b	4f�g]�^���?���Ba��`�A��~g��d����1j$���"(��Jff�!�Pb���S��s�R6��XCY��y����D;�܁�f�%Y�E�d�0�_��IA�<��;��qو�RJ���P%��:�Ɓ-��H�+�uj_U-����%N��Z5�l����7J�|�A�h��6Q�To���J�%�+٫]�H�������Ș@�SϹB����7�Yom�'sM@A�
�[�^�����31;<v(��Z��gHw�U�uBu^"<+0)�"d�;�m�b�E}y��5o��Σ\ww(��[��D{�� J�?W�
��p�L�}��Y��c6�&����������
zpv&���io�z�3&��i�4�`Za�i�El&���T!����X�QA����;)5?B�]�Hd�꬏C�J�'D�H�t��$��U�vr�֢��)�=��`OG]��p@�&�O�}o5�z�9��g}@�R���	b/��uGP�L��i�ך�⠿Zc��z��󷡾��5�)#iAZ��$t-�i�]Ad�Ƌ�kz�����76��9�i��Q���n�vY��W4��i�	I jvl��.�9��ȁ���P?�r�AI�&b��5��i�����C_�M� �7��IӤ�A���T1d(�l�<�vr�˫���;���]\]�ç��?���x=�M^���@��vDe���W��Gr˧V����$U ���OC����D:PXӬy1sq�ҕ�	�#�����*�C�0�D��d����?[�[n��6���Av��/�PL���o�Z�>XrjP%%���´T�o�5$t����z�$p�PV\�.e  �|�v�be���VE���<ǀ�_pZ���9rd��#�o�A�n���U���1��Q���i��o��Į������MJ9m��9&�`�ڛd�����n/�g����j�O\���cP�jjWE�-br-�T�M6����\�K����v�9n��T#��o�U�3d~`�oB0ڻjL��<���u"�}$�0�2c{j~}f��ڱ�S=�����8��`Gα���ޔ�
H�^	��,�;�szV���>'=��oO�]FD$	�����&+�:Ǟ V�p^�D��
��d��Ζ.� �*�E{���%���֟�@�OI��O�*q)<<p)7%D�s�!��u�?&2Gt�|BS�X��c�]�([����ƝQ)ݔD+u�����	"r���<.�`�Z0��=R��=<��q��)f�,}�*���F�/v�oH�������!���j��	zw=����
��)��.����A�s��n��0Gp���HWN�'�&����A�����x+%qIi0�*��i�k�w�6���q:;��kC����q���}#]iu��7P>j��I���f�PX~�D�IX�@��-�1_��w�¼���z�8$'���\&rM���nqP����z#/�� ��\h
��U�,����D^���TV�`��3�����hU9 ��
}�x��� |E|�`d�W�m��kL�~
;��� ��p�[>4^�9;a��_��ʨL�N�wJ��W�~:ԯ��
��<u�='9H�	��#���k�sV@̂e�E8��MY˔�´�t"��j��w^�&G�J�u�R:\�[&汌7{FlH�����!����;���_���G����=㺨�VR�7,蚡�\x#��p�r�1��?��߮��F�!>*�Ի�`�8=k�-t<����>g7 �va��ٰm���5���Y�J�Z�e���]��h<��C'�ÑFH�	oj\����z�$�
r������]�.b+�?G�~a�l��_!�[�g���ُ^��[)��ؘK��"6��X�Q���+�7��'YF���j���ʷ����p0�T�.?'Y��s�����,��/�GxS:[Oe�����o}��w���ሱ�rF��I玢N2�ט6��xԱB���27�P�d�뺢���-��%(��Q_��:����L�۷ǧV�ɲ�J?JP<�8UG���Y��q�j�i�gm��[��L���fŁ���_4ᗟ�7�g��jL)@B3���|��%��� ��>(�����=g0T:&��`;�$! ��PI����`"�����9�;(`�ou��P+l����$g(�@�|>�c�Գ�7D��J&F�P�k�;j�-.�iE�<tp���K���)�ć%��8��:m �	�b�FJx~�u��D�<(���H���8ѿ��	r��zF0C
���m>v�� �}9i���F�����}�=�K��=iDn;�8�ȝr]Qв�VZ�C�YN|q��l�~`�&Qq��T�T���ۯ՞֖�7�������0ӯ��TM�^��i�_'#��&���2���.�"�H��z�k2C?�)7$�-Nb;��ܰ,Xiv����j��$J�/��mW#>�0������������h�23�z�a�D�9��"]�f��lȏT�a���7Y�Y-[p�]��K>kC{�$i��gHGpl4ʁ��y\Z��X��|�� ��祉���~��~��0�0~�&`�E�l2�m6V	�t�B� L���%YG�#�`�ͨ%�0�����Z�MJ Cփ_�5=��*Z�Ղ�J�T'����i����aF��q�����\���A��~%:�ժ����-�q=�aZ:�Lao$x��_�\p�R���Yjh��/��6`4&LN�_�l��\��g�ڂ��~�����ΝF�ZY����L�"�s�����5�\)���O��~�'���tB�Ꮌ���XX�1���fi��nn#PΉ��E�䔗h'�0�Z���܀����d~F�t��=˳���(w�aW�ԫ2�?Vqx�?^���l��ܡ~�����[M�Zx#eZ���&~��t_
w&&&�2s^����%�,�<<(*��MPV1�1a*B$�"�/����`�U�5��\##�$���������aNܷNpYDc:g]+3
��u"0�"��c4q��ܷ^D�Ռ����0N7��m�L�~S�������SL�u� ���R�\	F-(u�G�򅈓!����gI���.�3xU�%���Ds/�<3=$<��)�7�R,����r�j��_z�P�h��AY̝p3��k�_t��	w�����i��R,��?�>��7a����˼��@�fP������#�__p�	ē2��ovMe0�ț����d����ӭ���G��"�ٴ����ޓ�܌ׅ=-ƞޞ��`�Nk3�<zL��0��a���vY�	���Vl�Cwi̙)-_��1tW�vp\��Q�|�ӑ���4��A�ߓ\E�p+�?�3�G|��9��Hp���.�W@SQh1���P�qkC�R���qSzo�V�'v-�ׯ_��-�u�����[�E���d�ؔ��8� �0��W��P��j�Dk{��DAkU�#��,q#���l�z7*�bY�=�sg�+��G���%}K���9��-C(Z�2�A���˺;c%�;���פE7�Zv���� Ba�q����*��\T���ck_��}���u<l�~�w�$�Dד��L*	M��3f�T�� �{�+�u��J�3�V�Z 0fi8Wb��n��Gu��D�mMQ�ب�Ls@���&mqO� ����b�Խ���|�8�V�b����P�;�D�A�ˇ��,9�\�;A
�s��-�-��a�Aj�H��]�{�L�
��x��&Z�c��t����Q8z����4�x�^�@��7}�lŘ����޴����c9N;��`D�QC���܂�R+0���>�A!�1ϱS׾\iآp���ɣ��(�d����$&����x_����2sf^%[x2㥣��q�2?K�nhP� ,r�hh�/��i"'S��	-B�# ��E�YRC�� Z��8��7���&/0��^�+'5�,ɷ���2"%�R�`~�D�1�z�y�f �ޜ� ��b�nJ��C���tw=�.�74
���}�k�>K� d
N{Ym�/k�+���o����},�)��F�[�i]�?��q���N�9Pn�]��ڣ�i@�Y�Wdx������Uٛ�/��1��&��Ym߭��8���[�i����Uh�.I��[ޓ�{����I�>�x�5��������7�K{��+�Z�"N�m�$@ҥ�ZMy�s�;\�����؟ �JxI���+��Y��V�B���Q�҉VߩYR�芣L�_aU��șүl���jP6,���.w��A�~�� R��G��1�cR��)zŨ��z�!@R]�-�TK��%�6R����(`5W[E�9�q�>M#����Ⓠ��q�a��H	2��B�F��$��?�涃��cH��0�s �f�O�4EH(֦���i0v/Xt�1ѡ�G
&� 8�1� U�Z����ۓ���6KK�(#�I~�c���2�`���N4�n�
�v�6��8�`�	k XS1X��*����VgZ��"R�Z��&�N����A�N��R��v�3���_�M)ݽ)X�F|�E�f��蠕�]�=�|��[���&E=�����z����_��Q��;'Z�4G�D%����֓�m�XAR�Ւ�Lb�)�*�AϢ�2y?a����Y�[f�7���+���DK\��J�v��s�����:5�Et+n�)-m���#a��k_nP���e��۾}�s^d���$V�Q1	�:n 뚲aͶi�ݦ�R|3���I�kD�<�3�vm{-��H�b�1?�X���5J��.0~��P�RjjzXy�?�Np��v5�[��4��@�"v;��lڍ������A�2c��ܿB����K@|+buNqAr���,+©n�^�ƿ��d��2!U���y�+�E�ݐC)��{����J<жIp��0"�}��_��ʩ�]�����e������K�)�qe���Y�a�}�p^{F=���l_�W�׍��Xn�<{�5��(x�-
�'TO���t2&1;���Jh�k����g�����ޥ�?��e>#�Kmw��jUC�:�(ކ�"2��[��8�[�U�+�����J ��{�v��N<�Aa�Yy�%���C�ksޟ�������9�k����4���16����R'����� 8�	�w����?���n�;�@�����~��n�V��C�<�X]=�l�@I#�V䌓�����S�����{���t풥jئ�6�d��I.����<Ud����/х��o�LL<3��7��u�]��ҥ�qyF��wL3Z�w�n[�!�Z��U��<�o 1#��ݨt�׵������a����މ�ĕ�?<��ԝT�t�����@˔��.Ų�qy�\�e�Rs-J#Q=�����ǐ/���5C�����'$#���*����l\�S��Th���i�T�E�D��
}������~@qL�z�V�֗#���Ш�Z�Ҟ�c� ����Fh�"�w<]̷!�ĕo����B.nc�Q����/��ClDA���
�D=�ޗ�ľ ���rcxh$O�'����J{�Zm63�KEo�U�̫�dZ5T�|��NH*w�C�%��QK��0��D��n�Um���fv~��)�L����1X"*��Õ��o��W��$�e>��:#Jy�w"��e��c��kUo��DI\���{�;����_�ô��Edf?ւ��L��%����"���|��	����ȓ�Ú�������ņi�-�������"�!�Ŝ#�x�{q|�V�nO�1p��G�7����C���<_0��h2���).W��
T��g��qt;e�b��^]s����h�6K�~����Z�i��{o�BZ@d2�s|�!�T�٣7C�ϳ���Z���5�֬"��R<p���6�D��,n��@���8�m��/�Z4|�w���PTM�Ro�.ޢ8?Y�3K�ʸ�g��ҕ�y���~�[�4sK���̱���O ����>��؉r����n_j,�0pQ�'3q,��{u���_;��u��#վ&�����'	����\��[��>D�����?)��+$,�V�_�G�:5;�$�|��e\N����9�]!�!7�^����͍��������rFa���7K�c�cI%�0,�.��r͎u�_[��(�PX�N�fx%_.�����0���Eq���c�曀��l�f�D4��~��*�le9��8�����TY���	 .���h�t�]r@����}+-���WDSZ�H���n��������)�����B��XYZ7=��S���%�"�����Al�\�J� �WI� ���Ow�����mnN�G�e��\;̬���ƪ�ڗ_��$	|��D�>��c��e��](����r��4u-ս����IǿPS����Է��X��Nr��k����{���ݵ��1<��mȦF�R�q8��F�@��u	����"kfY��P�pb{nAǓ���i�񻘽�� )r�}�������˜��	g��L,��ׂf�K��ca[l��y�#�E� �B��������ϤC2��g����a���x���E�7IIS7�c��̨ {���CN��>���>\����v�W�"c(w�=c3(쀍����ﴳ;�oI>%-�r"��Џ9��Pƃ� y��s��Oo��%���a2|��ZM��L?�9{,��v��^~>���������8����[�������+��_DSj�x����g*c7�Ċ�*��0��77�°�<�P��#�=BT��s��
�֎���V)âߊV:i��ko+��ְ�F:�l[KָF���OK�)q�|�,�jb�LH���m�uA��NH�?S&�e1`��q��$�iD�o���")�`�sKI�̉�������k>���.s<69�Z&7<��c�a�P�?�B�ᾟ�ә��׵xiwm���~0��?2�� �x]��b�F���;�.|�]o�&��m|�9�?0lq�c$z��dy�n��E=`2hJ�/�ɐn�g
j�ǳ-U�?C'���2m�B��WsL��k����У�/�[�<�-�hrY/�K�ce]��w�:vpg9p��OP�݋�kd*�«��?�"�q`�@<A�&p���~�I�R|dnWշ6����i�ItJ}��;~dɠ�n�ƿ���<�	T�|�V<�i�5��-R�[��]V���uH��T9�7�9������<���/}t�V�lc��ϱ�-ԉ��咪�NM�������b����ñ�~Q����}сZ�����'7\-�#�����u�L�=|q��KY����%Z�J�q��+ǲ?{2�V���mz�֧{��s#�ۼ�����vv�b[�jUc����Fvl<�ev�r��9j�c��*��ѵ����Y��K {Ƃk��ΐt�?s4KuI��v�:��G:�Y�ۋ�J���z�U�,���l�U��4ߒ�>��� �Z�Lt�#��8���Ƙ�M~���[�]lZ����I��o亄!^�^�Ƴ��op��U����+߬��{0(!:s����xf�m�|�O7��m(���j�{�QR�ȉ9�֐QkP#�Pv�����v��efեK����8%aE�~������Ѕr/G��#��R��=BH܉C��L�oּ�
��o�T�n�D\t\����d_��O6�ʍ/�l|���C}Y?�/lO�]�	j̭Y@�pL�L�e*3����#�Tg�r|���^`x�hx֬��	4k�b�4~�:���Џ�5��qo��g{/�����A,w�$0������&��Y��J�~
��U��um#�>�~� {i��:������2#��9�����s��ZWn:�9-ܓ��_v��(��Oyi�#�"�mo�ţ-CΊ�m	���u�ȋ#0��.��@�o˾�{�'���,�4z�`N���G��d�`���H?��&.���x~�;��m��#X�Z��4�GE4?�ҁn>���d#��/Mka�_���7��$�,�<1Wp����Cu�uO�~�O��42���L�.צ��ӗ�'�q!
gi�o�m+�T�k>-�R��ҏi��-7�`���>,�GH�{]�o������'�*"�N<��gmP�StM�"C�I�-TA}��bH��J̥�x��3_���
�Xle�y�a#�# \�9�h���d;\uf.�Si�����vF��j��-qWW*�B��yF�)�/z�AƑQ?M�0�Ջ���o
d�J����L�ڛ�Y5+�6'6�p%5	d�_5��A�Q'���������zo`�����&�g���PX#�_�����E�V&�^�'�Y���vC�$���Ȏ�Ͽ#z?|��ފ�LK~�|��_p�`�Ј�6��*�gN,힑)�E�0�.z�u�����T��hR���q���̈́ɦ3;1*��:�w�$D�f����n��h[�֜�s
�H#�/p��#߃��x��23��/@ߟ�Ǿ��GI�hLr�8V��ԥ����ç���I�h�ϒ*e*����Em��{�|����b�G�7�G?6��6�f�P|@�_�O����.��(d�u%��ü��J�@z/�6�*%�����Kg��KH�|�� �Y�w�vēKEB�+E��:d�q�Q��hzR�F�MH�g���?w�?��ӫ<��m{K�s������U���ܵ�xz�g��_*J����e�]�����YK&ȭjC!*��w�������3�X�K}��Pu�riw���q�Gl͸�[�@��ʼC�zN�����A����������:D��f���?b��R\�� R��]��F��4BŢbl{��4E�8{i-<�>��;���c��D���i��?�9u��!��ki���c��<Y�%?�*�x��B��5�P�ZQ�x��{Qxó��xx�Ǐon�4S������oz4�ޮ�l��,2�W�@7�k=Zb҉p�K��J�|I��ǢG�~�]3������m<#�3ҷ����Ԝ�{�	�B�_�O���� ������V���q��ᆉB�m�8G�(/V��.+�f��M��&lEnoK:i5�
>l����&�ȱe�>���3�zh}<B�+ӊ�s�8̟p�`�R��E�J�E#��If��b,H�D!.+7��Պm̗P�2"��/;j��c �X:{��~<K�������(A���Û�r�{-ao�$� �?+�3cwziW�c۱;��0`=1�]��������L_����x���}W_�T�k�_l)R�#�|n�*3��ꑦE�m����C߻��z�踗�"!ݚ͕�����%�v�-|��4�5f8������'�?Gv6�}12PpL�v2љ�ޖ�MW4˛}w��6�}�]� �9[צM�~U���j�bu��������=n#�",�6�h��)h�ʍϗ�j�I��E7$k^G�/1I��A�t{w�^���՗�/�w��kԅ��7Ĺ�������1؏og`�9��̂!�6�������=��7�}P߅��%���z��z|)?l����ugC���WU�!�2�S�w��i�
��qX�<��P��7���T��C�\���R�Mv3\�����?�,ᙤ��D�G�F�}�V�V��E��k6�V��q�)�W�:�����$�,�/�S�yu6\�G�oW�b����6�n�mu��g؎��Ctф*�f�	�w9��t
��|����p�����v$
_�{B]�=�g �n4�вt�[H�d�wy������!WY�>�%eѳH�	 ~���P��"Nw�d����V^��C�^��h�C-`T����gs.;�Tή�d�y�PX���׈)����;NX��Ҭ�Y�O�,TD9�h�ɖ#"�Oh��6�RM�#U��%HNOo����x�	�C͚�~(<.L��d��!���wA��\��4?(RRF�mz���\)��y�o!F
*!|�T�ο�}�o�@9E]/��bO�bEe�C�uD��^�xT�FC;�`ߎ �"�Io1Vɏ��sê���[�A���Nkju�)��OrGe��?��=��D��/ׅ4��'0U�=K���J�m�R�\���U̕��I����2�1����&�0�q�񃝳�c���UU�4sZ�UE�"�u�9by��H����5��e�T,w����i}�g/���+�;��GH���8Hu��A��6��1w#���Jn�m�iiV#��#A���7P\Zs7tF]̮X�ƚ�2�To�5�k.R��|���ɫ^���n���})��|�hy��T�.��G�n��4*4h��_��1�[ƈ����%��ӥu����n/�}7���ة>�Ogt��]�9D��q<�r�f��a��g�ގ#q�b��r$�h����A���s��)����G���oZuɣ����*]���Mˢ��m�x�"�:Wbq���GC��K��湣�v��A����ԣ����®ױ��Ŧ���|#N�(�)r��"��<���U���$�Ξ�+�^o�f/��/��v='��~�w(�hZ��ms�w���՝��$ͻ@5M-��MUB|ZcW��[�Y��%a����p��Q��qv�����j�^��H[}cP��SzZZ�M�wB�q�M|f����f��b%8��t�zY���v��V0��$�Mؗ;�a�d���?*յu�Z�O�:Y�Z�A 6�CZ��ڞ%���2�%��('?g�l��)W3��ѷ����{����?�������[�+���;�q���2`��}�ƉЏv��q���m<H�$�O�~�ъ�X-�cE�E���kq�"�d�K&'��5����c_�qLF���/��kL7���>�e*GL�=`��v�% +�L���X�m�L}�8<8}[2�kרlϽ��̎	ڍ�"�,�c�fL���.�8X|��]�{�.=^̠210�OBWEtD(�Z��eg�Oϱ�{ ��rb�����§�	�������C�3d�俯)���x<����m�v��fn:�j�SYހ��z�
޺dM�ij�R��4��;AArf#xs}�%�.}}����P~m��mj���#��}�둁u��ۭU]8Ӽ�.K3"`W>��E@.u��WC-�۾ ��L��};��r�>ߺ�� �'�F֖��Ri���v/F�����sC������������`�W������M����j�B�IlPl@���}�Ŏ���)�X������h2�#?�$&m�������0!*a�X IeG��7�2$]k��s�Kfzb�du���y���|I�u.�K��L�B�6a���ش��ϋ1g:�MU��������uz��G�����NE;M�/��b���M���P3*
�D-Ň����{H�⋪�}�g�?T䑊����=_���O*�0-�q|�Y���/^$�W���۝��~$�J�r7F0���`�Q��ج��y����c�<U��a����}�5ӵ݆�-Ɏ-�^�T�oL�k_�S����'L��1ZR�fQC2�����^��_D��l�)�Tc¢k�A�!U��.~����O����Y�N��CV
-L^4�n�Js$���;�kl)m��`e'�u�U!Ι
�N��7����ۘ�w��7@A�%�a��~�e[$̊����I�m�O���XSH��6���b����=�Q������
�+}tۥ��7��F����$�t��ǹ��S��\��&WBv���JP���wԉ���V��-�vl���uU�b�.M�J�4���dlT������a]tx|�K�yeq";���#'`��7�FcF�Nj�����g��G]`�~| ��O��Q<��4$Ӻ����[_Vz.&mk;_�`�AB����Un�~��|���j!�Cq*�/�2"�񆗿*�f�3�qX�q:�D.�G9����I��P�E5' 4 �����g���dg�l�B:I�>D��|1��B5-=L���V)�lE��K���k���L��ƆE�Q%��C�0�ax�N�֊t�
��3tu��=`�V8�Ko�����/�iE��-Y��Iݚ�����oY�g����o�j��]�6G���/5=��
M�[[P���� ]���z(nzf |	㯭��p�G�3��z���Ը�f��4G�!�#++���������8�����t�v�!���ǥ3�yUA�YS�+7�ZCތh�}������˷F����2`q�y��gW���Н?�Y�!������53c�������es+����	��c�U��RAa����9l���u$7a)�Bq��3��=�� �?�o��(�W���,f��֎.s��2�_�8��3�����5� C�2<JMR@m��܀[S�2�F�6urgח�s[����,���"8MX����a"�����Q��܊oz��z��G��#K�����s���<_�����P��/��韪�e���j!�,��-���.]ml�͹�/|� ,@ӿ��+��@`� ���壩�l��@�ϔ�s��5�ư��D���Z�a[��: 2�X[�O8@�SO=�_7��{p�����k�Ή+�o�1k?�oF����*�+�F�'��Tݭ��C���;�D<��;	R�͞H��S'O���޿��~�Y����BZ�S@�1h5q�D��M(�M��2�\/���V�c���9@�ռ)�Tj� 0�ە��rb���EM�Oʧ��2��رc�����->-����������">�@��*���z�N�휝��o뛔v3�ؼ������B��R<�xo�[��vV��@ɨ;s�{�[{�J�(J�`�O[Yuv���v?ݓ���u1�c� {E��}��_��^�
������ǏP���=�t�BE6E;�ڻ�A{@i�gC�]�CL]�S���nx���p8# ٍ՚�F_�&���������
W�6_��̞�3�k��f�d�I���r�
�M��V>��<���ӡ�#���?�������?�{��.+vw�3�L��h,������(�W)�7_�J����3 �ٳg���}��)>���l�Zkz�R��T^Ĩ�r�T�G������$&�u���q�5z��15��꧘�EF�c����3�G�J��g�K����duu��Q7ϹsH~������m9 3 >�y뭷�w��*�� C_��#P�e�k�S��a�u��+�"e�	¢�䒆��u�%��w��%�'�!�Ge��=~���ߤ_|��jJ�5Y�$����m3��::}��Z�c��*}!�ˊY�5�?�ׯ�(��A�<�i�����nJ�033-1V�*31\s��m>N�O��.2He|��M�G�;�dm����?�W_�%MO� :�o`f/���(�Q����-h�k�~
���v����X�|04�M�u�6|���O.������7
�Q��4�r0pе�K4q��t�A\XeJ�
����i��u>� �u���a���8���n᧜L 4=;C=dC�=%3�v@wn���-I��uz���Dp$���K���Z�nx�<=��?��O����қo��
�f�d\^�8��ׅحd�Yk�q|�Mf�]\\�'�x�A>�5P�(N�>�ՠ��dܫ��ʕ�5�X׼Z���y�Ցu��(!���κ�ؤ��V3���*~�&K�n��X�سN�>>�	���K��+��N�Ϳ/M����l1�v��.^�H��ԧX��d��	c@���	������?�yF�?�я��?�PN���"��ï6_�f넪3�u��F�ǵۈU�H��h��k �NR�+�S�����_�2}�K_�J� �~��L�0 ��n޸a K��.�Ç�Q��5�-ъ58M;����.>���a� �tUm-!��^�z������p��a�1��föz-[�?�2���0�R�(�bb_|�̸����[os�R���`�.��d{�X���[��qY7vK�*�u��G|�v4:���z4���O�<H�$�7�@��^�2���.�3��a�@�ڝ6� 	�M,����}�ņ7��jth��*�d7���:����y.��S�Q�2"��xNF�f������4E\�Ȁnn���J��d�[����MV�TB��UrՕ/�$�nڥJR�w�t���=Oא��_�+]�r���Yv����t�-�,'�;"�`�:�Z�XNMN����Ӆ�;��CE~Xl�w<`��XS|~��eV�_�u�կ~�mj"���l�dsp����˹� �r��I(#��s��Q�|��b��915 ��o�G���Yi�3ũv����[�`�d���`2��ca�� Fp0��}L>#I$����7���/~��Ł�bh!.x@'�]�����4w�,�8�a����J��ݻ��M�D⺋"��� 4s3���x��b����9ÀV1T2��ly��ךt��I:q��s�_�J�F��Xop�4+<O����͏����ڠ��Ԃt��^�!a�[�f��0s4�ul45�pؔ�V�n�������(��[pP���0����y��?����V��y�Ԝ-g�l�F���ܣ�a����������ힻ�x�{�݂���2�wN�,3ܷ8[=o7����I;�öWf��Y�q��SO_����ߦ���;��Y����8�8jHpL�2��ll��k��o�Ҥ�Z�ӓ�` ͑�t�����F�A�ɸ"xR�9�A�ȪBY�n����O�4�?���e#���i�ǊJ��fElv2�q� �͸(�`9l	��Z�������u�h"��
���rF޸m7{�����ɉI�g���L�/���;�~@��<<Uy4�৐{ࡸnȼ����l��w�r;y��Z'��8>H]���!5� (�'�k<i���}5:P
X���
C-��^��#u?�F�
��	 &�{��y3h�6 <�n80��ѣ|?�8x����51Ѱ��_L�o��k���� (�G�c��;.S+������Tn��;N���]��&���[^�K=i@���:w�m4֌��s,/qW�YYY���Ct��iB����M�{�-4�VGR�m����������P0�.(��u��d������Dlu)�6�qʀ����liY����!e|~~��D�:递v��?L_}�%��t�����>�q�ko�Ƒ7b��؟�{~;Y��v���O�m'H�	[��|K�^7���ߋ1T��
�{`�n-_�d^���q.��Z/��w}�F�Ξ��|�[��s��R�D+p�g=v9q�#�Gʮ�(�5.#�)E0p�K�o�ҵ�o�p�&�5�էi�>Au�;�g>��R\U�(v�j.A�I�	$�t�r� V$j\{�+O��Ɗy���%���R�`58^��� >b�S&�W����tj��h�*��9��o���8�1��c��qւ�z�5�^��z. c ^ T�9�p;�BҴa��u�#�w�<�[f }�Ps��m3ww8�a >�ѣ�о���}��N��	y�1�����-@�J���1��@�jt�����P�&�҄�;� �ψ�Έ�N$!K����M���k|���=O���7����<� )��[������FXx ^Xh��+��x�N�sQ�,-��G//*��|F���r��M���$�-����E�җ�D��ː��9�u���2�Z�E��$�?��C��y�]��k�2��f�������0�C���!��7�֪ԁXw��(��t�(�Q+�d�Y!���g�y�lJ�{��Q����cG���������l�n�h
�apj�[0t��Q�w�]>��o��o���Q?�۸�a09�������\;	��Z^v�*�>ϟK�Y�?eT�vu/<�������І�-Йی�Q7���ƹ��P�qw��\���-rt%>CVṇ��7��5��
,� � z�lƅ�
EQ*n�4�J��n��o����� � *� j&��m��-��J��6���3�DZ7�l5�ЭTl񵘏?��`�+Qc��V���X�{֟���f��f�#'�������
��l���(���,�ˏ?J�����������*�:,���w~��nH=hc��O�N�:E׍l�L����P $��3�4|���+u���iVх�.�7�|�]��g�
*ڂ���-�ǅ�컡]|/�,��Q^c�$O-�G�k�#,>��:5h+���sWx)�[���k�6��NA*6��:� �!����iԥ���>G/���^\��`�!��p
|��`L8&�	���YZ�`H����gm��BA5TIq.��V�e ��ߡ�$kO��^y�>��s45;I�+wX�8���B7��bk͑C���wȵM��z�d)���@�g�zz�4�u�pӍ�\S��|3� 	�A��^r#Z��n�ǧt��⮚6�8���Uds�Q^�TO�I���}�[��������W_}�*�l�!�i\��F�H�;%��Ҡo��!|�ǝ�*T6�?�'h�
��R���xh�j6�2�g�e�s�\�F�}���I�q�i�9H !s`erz�N�<F�����/~��f������G��T.G�Zh�-1[��l�A?�v� ��u΄,��J�g�5��8hS��S�d�!���W7���B�`����赥�M����W�f�+%���~��UA�/��Ck@�F	C�2R�Q��"E8����{eQ��Vg�-,ғO_�o~�����s�CpJْ��4 剐SP�/��(m��	5�`�i4b��|�]N����Գ��a�ao��Ǐ1�<CH�C��g���_|��S���=YVK�a�Éq�p_�a���~`4ch�-5������T��'hc���~�:O�ޏ�ty���!������(��W^�{�At��K/��	��\�6 J�͡�%��H �>,
,4��5SF��X�{TS��ڸ�Z�V��b���o@��yČ��4�0�~Y�g� ��{��l��o��ƻ��A�KK�8s]�TK̔VW�9YgK��h`20H%��1A�9ku�v�F�	�@5*j2((*�3���_��m�A#"	%�''��t��l�e3G(�U5B5a�`ʙ�4f & �8;3O?���\�̓d�4s{`�V��ƹ&@{]+�u{��U6�����>��
��7V��;� �d?���Q#N�������G�ڦƹ��!������~���?���I$����2>07c0p�(u�/;u�8�9w�N�9Ů&d�(�I��͐+q'�<׃`a� N�^_m�9�s������(�=�bP���~��?�E��47=A��	��	2l���fy��������@�S]L����2����H��D��(��`k.��	��(v�EIlZ��'��/��|�
����ϴ��bEH�6�O�O���	!p�U��/|��w�0�M 8��;!�C U: ��
^f�2I5��Ȅ�<{��ez��X��|��B-�z�S�eHN%�W�Y������S�Y�-��}���l�_5k���G��:T��t�{~T_S�"��_��\ ԅ�UR��zn`�^�`�;S��Q���$�� Y0fL(�>�
������?J����]`qv��"��M�}֞�z��!��+/ӅGf�'4����u�;�1��1L�F�J�,�6�Z��.'�!�P���3�7���?u�9���=ͥ�d� fdD\14�+<��W���O����u�Y�K6�;76ۙ�'`
7̪�nQs�E�M^#r,^�PG�\8(s�0�s�f�:��x�-k�+���>�e+���
��������s�? �`�_����_���Ѫ���k'�5�Ώ�c��b��ٓO>I�����nc(#
pe��x�MOM3�Ef"����QQ�E)����o�>�J��t��)�Ξ9s��;�}���Ǟp5`p j4�H�q�`�l�>5׻���T�3[o&���̳K��*W���Õ��V��q�ocEP4/�w�M1@��g������<�n)�֞���xI�9u;}�o�Z�X����"��X7%��O�<n��o�;o]��ƻ4@�@;0G���*����B �� �G9��6��;q��9a��r����B��W�;��-���S��	b~������u7n�(�Q�T)�c��H��LX��z}6B�����f����m$ 5w�&�sS�h�|�hkMW[��Č���T0��I���QL�X
��VϛҊ�x�0�'r�A�=�(��,�͛7�"&3Lk��k��z0�����r�ŏ/�������<�֤�0Ν;M_z�sT���?��rPٺ�Z�nܢ~όeM�.@�;�+\����I�
�G`h4>�3��0��O�'E@�X��1 )�/�GF�}(=� ahj�J�[
�h`h)�52�3L2�md}��~�ɩ
��Viڄ�
����9��i��7����͡�����v�`b��ɒr�{\�w�ָX��AY�&�} �l)�Ch�{njj�-9���޽v�f�������>���E�njf# �2���t�҂	��m���5wӇ�x�\'O���I� Tc:�,�>��
�3Vt]���
?پ�mؽ�E�z���ؕA�� �X���ZL�"�@�1�K��b߁WgE%Q���R%6m�̷�*�
����;���åV�GB)�#�Då�8��P��>-nꢯ"�t�YA�#L��1�p��h��.�]Q���Q1���g�϶��ڭ�0zmdy�z�}{���Fi��ri�+ԧN�f��'c�����������-,��-p�(.���e��/~ᬰZ�ï��b'mӘO`O�DE�B��ĉܜ~���5���}w?����l���j��sh�B�Bm�E4�N"���A\H�������ɓ���K"x�p�D?&�l���9�ҏ�A�-$��nKKKV@�n��>��go��&��
��~��(�O��9�A�`X���v��ن1�,~�������:t��#�ԧ���N37��U�ct3Z�ݤ���ш&��Es��hL�
�cm�	��8G	��u~ԍT��++�?V���J�;�;�V�H
t���XT��*���'�&Jd5�F�o6�K7�UÅ��F�Ra&ʌ��'<��G����n�u������/�^5�:*ļW�n\!����8+ɽ�����~\A�q�V5U�zD|��i�1����qp�^���r�*����%�_�+Æ�܏�IXx�������me��k���M:7�+{;�#mN�Q�8����S�_��/�����B���"�	תMQЖ9�V���R��q"vʵ��gd��Kp"��]5�#6��<��U��l�X���|9����$Y,V��~vYO�� ��ǃ+ER��>�9C��+�l'�p!;��֚�<#�;����b�=G��O?I�^�b��0�9	%�@��T滥�qۜ!�na�^��`�C�F���d��;B�F��Eԗ# iL�|	>CQFd�޸���9s�}�<����L}ĲSc"�M�Qw�!��]�mbe�R���)Ïn�˃�pJ�j��s�DV ��I08���,"��4@;���۷o�3��=r�[5q�h.�g���#��d�݊yFd�̠�\�{�9~�[o�e�uF�r ��Z:�Pr9
~;M\A����m%��QdA�9�^����$�� ,Ҍ���0 ŌMb��T*���,� iqZ'~�!�j��l%����^�Όl�I�-S��}t�����q��
D�c3xj�Xp�u�Ynwf�D5�Ls}��g38��Mj5|z�`a�K��F��WFC����E#��~���hnU�O�j�����@�~�:���N[�|�w�����\�V�ӧNs ?J(����a�)��ŋ�ȑ�f����s������@�w��]ke-�4RM7݊~]�K�K6�u��	Y�k���t���4k�t�(p�Ξ������GÀ�yQn+�fH�[a�<�����}Ɋ�4�À��juXe&��_-qi�RR���9㍢��$)�5R���LL�3 ��T8��ft��&ʴ�~��78,̥��h)����D- .���CJ��8�&�3Ĺ�'��&�eh�.?y�^�W�����X��RT�^'��.�	Y/ ���q�'�
�i�nx��La���h`��_*{�\ ��#|J&����,S�@��R2���۠\�J��O�	��X��p�*���1��L��}5 �z��e��h(X[$��9Q����l�E��f��!�b��}V�^�0_��RԜ����-E ;8N�Qo��6*<�@�Mm�Y1������f�`¥����?�6�� ����A���
 !��x,C� ���=�u���Rz,X>SP��r/�B�0�n��A�
@��G�L�t�<�NSF��s�M��ӕ�v�`H3E`#R���߬Z�:�����OA����l�U����t��1�я~L8/�䜒����`��֙?�~��󫓯�X������{�1�n���J@)�Q��`>���a{r(-4S��~�����Uz���'�"�&ɼ�D�	�Â�(�����	�������st��i�����<�띃�΅�v �p�!Ď���m��81:�R5JCŀ=�7��K�ĥ"k�c�"��%����~�$��b<+N���k�-�M���4�ϵ����qSd�&��ƿ B�α���4|��Ir��X ���R�?\�G/=Fo�s�~������Y��{8����ݛY7������
�؈n�Z"�Ҳ.���:ד߇����nPb9V�\e��^������ uJ�h�Pe��^��>M��3�����@:2
�<���:@��ں2N�o�ZZ�7#5�� T5*[���v}(�m/��sS4~k5��j�3Խ�]��"v�8�+�7(�=R�jS�����O�܀�K���Y�#��l�� �<�xqK�t�	�h��>�J��hP�@6a�����*R-_���y����`A�Q�86@i�ANo��l���)��i~f��CLԳF�����3�v��%Z[Ye�<4�ڜMe�+�?z�(�^��;,s�s�ݻ(o���@�G�c��=�~�z���k�w?���7�1x�%�����K\�MF��ͿG�L�K�.1 �߿앁P� ~����~����{hrz����*�i��_j͕� cQ�x���sѦ�rw����A�y���ޢ|�6k%c�k����D�o��I�% �3��l��%#k�fw5O�A� �q�i�b�!VX`]E�>�}�w����D�kM.�ϡ2x_(A0�D�:#�$��(h�)gG��_U,6�����r�N?o@�F�̞�}�6���Z��~�n�'����$<
�<��pc���CW޽��Y�T]�n�w�| 幸��]����l��w�(wH}ǿ���Q�,k��Ak�xV�	S f'�t�L����̌͘��Ǡ� $��M����W�!E,��&m��2L��H<Ʒ{S�����>�v�_͔R���%͆���s��bdJ>@P��._h�l|p����˗�N��!)�iu��\�s.fU�0��l4}G�*�c���!��k�
q'
3�S�an�l/���1FQ�_�"̢��K������koPv|�l�y��ň�(��Bݴ9�s�h}�v�煵?���%V
c@���|ی��:�� (��M{p�em����^����G����Z��o]��<����Bf[c37�Ga�9y�g�&P�̹�6�B��Ι�^ݝ~����}��G2C2�j;�biP�ڲ��_����R�<�мf#��b9B�s��=�nFh#�G�0��l����ь�XRr.Rg�Ynd!W.G�L<�d� ȈHΑ�)�Y�`�,<�?T��\,�e��g'8�ٯ-J{��B���r-�&1~HHS��Wy$�D�j��2u������W�"��.�R��CY��68^)�F�<i,t���[���}x�Z�2:}��:s��&�l�3�����%��(o��[F����C/�-\�X��]��6s�VG�J�T| ْ(�H�8~���ʩ�> ��J��4S��^�\j�X�E����鲀GS4�L�˶~���ve�I'�<S������eaڰ�����+�j ����׹��ڔ���̥��_~�G�ֆ��)��f+P���t��t��a�:|j��{.҅�t��,>�c��
} �@S�	��i�zԅ�RT�'A׵�:%`���U'qY3��!�zB���r�q90Sc�����UFM��8��\�hj����x���Fh �l�i��#�.]x���λ�чK���'Y�������=�C[{�w/���=���|�0:73G��Xx_��8��o�>-~�NGR���������5��w�Ɖ�k�g��Ck-��|D��d��_��LL�L�YjX������Vi}W�S���>ҴG�=q��=�L�+�&�����%e� �s�'�*��"�[I��5D���}�m�P &=$����o��Xj])Љ���'r8���dU���f�S�9И�kDFp}�\)�Pr�<K�d���P|X'ۏ"�֫�%��Op�Q�nv�7�j���v?��z��� :�a��46�86��i�t��G,��%��Ëv� z%���W �	>��t���Z<7�Yw���`)/�r�
+��y��*[�<d%
&"�㉵��>z����s����s?��������7��:�_Ddfe�U�]}�э��(R҈")��d��=��lg�fk���v~��d����F"RER�	�hW��FW_uWeeD��>w�"2���*���UyF�xϟ����lS#�"R��a�4�B�s��w4�l@��OǺc$��wߊ�K��O=	�5�~�inx�.q�/�w�|�"O��4�v�0�8/k/�Dթ��7o"7���X����>�Qw������
g*��_��y�/�C���A��)��[*�J�1���X�X�'����rB؍�b���L� �c�c�0�\P�6��\�p�h��eqiŝ|�mwxi�;|d�Cy(�9|�F�rُG�;4�F��:�� ���pG}�s�ڂ�z㊿w�nn�>w��TH���Z�h�.���=�:r�� ���V�z�ԧ>�9���� �h>	���@�/��������N�>C�=�+�_�bǼ�}�yִ�ͳX���������o[�&���p4���g`Lf�g ��c�Q����$+d�h!퓫�R�<�WZ)������A�/��6����I`J�0���q"�B
	�ep�.)ĩ��&�&�q�_�g�����%��2�����wf�r�JXz��V�+8���D='7W��su�[��U���Y	��'��'����s�*D��P��=oۭkVܖ�-����\��i�{��i���~�}�3���c��^'��*{��<�.P*z3�P݄f����c�]����^	��{뭷9o��O8��?wY�ѡ�VE⦵�5%��޿c׈X��`��xqbP[7Y,$86������y�qC������X6�k7��NLc!U�<����]X����&z��6�|���Xq~�J�&�#n}c3D����%�����G0ds����h�"~��L�O�����q#/�RSA����b��@���y���T۪��q3�1�����As�����&�AGY�x<68�Z*��U=����|A	h�������V�3g/��׮����^BLe|_^��1��I%H=����>읻S���
��;v�7|�~�X�)�=��i�[1^[m�[P��R�sfm����B��.�]'iIl�0�������XXXt_����o��>�я�t/ժ0���E%�'�^�30l󸕱��ko��K��B������Cc����f(������#!�w�����g�_��H�rM�g n���/LRiLnM�u��e�ے���QZ	��-!�d�(m��>��x,NM���'������ga�n��?�m�_�����ޣ�08��p��IIǁ�$'2��r��S�n��T%�u �::>JT?��U��h~���ġi���}����{RAY���y�,{JA=4�'�$dj��u�@D���j_uP+'�>[�9�/X_�J<y�5��X�� k�� �c�C�~�q��8`�Q܁��q��S���}*�cל�lr|�+�G,�?�q�@v
)����F���
w�o\��c\�8��Y06�P��+|D��c�`cgO�e�&��������9>�h��&I���i�~�MM��Dq��8�F�F�b3�.0q����%��#b�v�z�m��kQ��7�'�������é�����X�E���
W	Ɨ�wߋ���^� �@��\P�OH��*�W�Xt���Ohu}��Xap���DVqw����n��n6�8/�����~MT'������mF�\�b<E���$�(���ڀC��o~����?��9v�A1?P�m�����@oP1�y�ノ���ǵ��0�#�u\gl��u;���jDtF0>p�77�nϾY�@Ay5���B6B���`8)N�*���"��P_ȡI��HZ&:?%�Ӭ����ag��¹a��%�FZUaJ�&�I˱�^�J|�����;��hXw�+k����X*�s�[Ŧ�����:�i�u\HO"�wB7Km�e����e�]�[7�H;J�/|�~N{'A~�=�Ի�(2{��8"XO�* 93;C�k�b��)^�@84�a���_~�A�*�gh�q�պ�8��s�NIY
b���}�Ӓ���{q�kHM3B�+��J���&����RiQ<qm����^�A�΋7��I
��׈^�9���={�O�W��M����r�\�ɮ��?�~W3*��ͭ���aŞϴ-=��M�L)"Qh���ކ[�b�(�2�
 Lrp�B�J5@̩1���7���m)��eK���`ȋ�*KE�X�S��P���+5Iv��K��z�Yj���.������Z�͗�rw���ϧG�=��sJ��a߲hlKR��H�9e�@��j�ѱi����q/�&J�~���4&�_�zE+�Jqs��bCC�Ґ��	��o~���S����׿�u���د���e�����ձiޛ�"�X�Xs\j�
����~[����Zj��+Y!�9�R\�]��x*�w(!㤱�S$��>�<
�(£�O��7�.�[�B �Ĥ&[��UK&IT�"׊o����j9y��ඁ�� ����G�SR��5w��«��B5� [�m:$�\T�%x�34�&�\f�����.�+��S^ʥ%5��ڼʭ�{��!��u�4���X�r?��O)`���s�xnq�wP��ٙY�簝��N̻�W�s]a�<+Έ����O�<��}�^y���|��2T�NK!�vH�Z��3˵��������c�85�RXń=gѱA����>��3��}���~�'�f��u9w�v��KN���"�0�%����x�?�я��R06��D�����bD��T9�X����^�d��	}�n2^v�e��a����grr�uZm^[�"@g6ʒ׸������~�:���Z�d���P86���6����.1�R�d�C$)�9��#ߤ�IW����%X ,B"@Y�� ��isAD�Z�~��؅��;u�������W����阶���=��R�8F8���s<�|��1q�ht ��1�h݁��
ƾ�q;�N+��gk��oW�&� �O�(������}�MF�Na������|.0��/�Bmˡ���_^�]��[��9a����$W��HCA�Nx����B6�E�"�'Hу�0�xڤ�j_"�ؚ~q�͗�r�m2�)R�bN�����P*�6J�������^�}��|(�4L!�6v9Q{'��L��7q�ŝN��S\�~s�����8;HAA���ʹ2ER��IҎKT>�*W˰9}̟W�%��@qA�Ek�s�Έ\�]{R�l7n`l��v`l�B�Sɻ�s(zi+�9�!8}��Gi�Y(s����=?ǵ�}`jr��m�K��c�	�N��!r>�"���+�5�t>Фt%�E��y�F�b{�s��]�<ˉ�I���}�vױ��&F&L�&��Йqbʧ]56�ʜFs=����������s�p,����7�.˘/]����B��~VFn���ı!�+�����.�_a�d�ʚ��K�\�LS9%ae�����1�r�$h6#��?11p+��A��+ؘggf�ǉ��@�(�ާ��E���$c���n�O�����%�)|f�k}�N���T�Ƚ� ���ρ^E)%�,��F�����L����h�V�xA�^��B���_ ����y¤����UOlʗ�4[�7�T�n��#��>P���)(g������!�.P(�A�� ���'�S�q B59Agw#B	�2F[�k�#q���^k���k��;uow`c�s�jzǋ/���������կ~�?����S��˼w��W��V֖�����d�=������q�����O~�:����?��������SK�dP�*�<�C������w��Ò6i�1q��6̥ťJ�g#{I��=HHr_][��m�oB}"�ݱ.�>��"���M {p�>%̂"m[&��a�RP���MF/��6EY:)h��;J#�n:T�l���K��:f"�����YD�F�%�2I6r �H�9�eR�ETi�ہɮ�@�����K�h��?��7(��g�޴LB���-��oc��M�K�U'�,+Zߗ���� ��d����Un�-,,�W_y�-� ��G�p�I �U��3p4o������*�RG���8�T8��,� Z�=��
@�]��~�~��66m��(G���z�F��~���N��+�E��ܤ�T�Iw��Ŋ{��aP��
�Zqs�}�Yt�FY���;4�X�,k��y��X�̠J�+�{�G���>ŉp?X��_#}/J7C�U�`�z0��,DUVm*�K+K5��f�cX���ai����3����[&% P�Ĺ�A�o4��c�.����Ě{
��'
�f��!c
��$��|����(Mb�i@�'�9Z���}zv�%�/�l,6�Fۣ��:�{;pn2�O��������'Ƙ�����
@�m.��~�q_�QIs��K�H�;N�(%u����#7�k�x�[����F�X=�ǩ�|й�#Ns`�#���t��S�u���S�%� ø����;v옿�3l7�'�G���G�����s�Q1���щN��������}�ʸ��?�F'F}�q�=��7ݿ���v�w��U���SJ�;ADoy�l8I�W�w<p�k	P'[��u<�O���� N	"ilH�g{������_C�'�.l莭d\�!e"��N'v�٬�3GJJ�������y}>��˞[ﭸ����{��%+����(�=	����p�9��R�U:O�)ayv��U���?>�@�N�:Ӷ����S%�V"]�IĢ�cݻӀ"���R41F��_]"2|����ǲ��:p��N��a���h�K��7�}8����܏0p�y���{s��2tlT�l�����_���/_f*
��
H�X3�C��S#zm̳��V����!1���"�����S�R��ʀ��flX�[�T���06��Jd�U���}�9%R]b�7�b�)t��u=�T�<Ah��`� ���?�N�.��p��.�A�Ε��4�,:W�<�=�k �&�wj���|���?(�Ѐ��<����y�m*2��'p݅�!�0��Q��������JS%
OG^ߡ���hK_���C��$�
�?�[�F&���q�K�����H3��o���e�)� �b����8�+�t���������w��4>1E��%����d��z*��5rȸ�ss{8Ϯ�_qW�$�O����E8b�=(&�:j����gH��sz�r�L�9�l_�g���5���|���������epn����u��#�����������;@_w'�
7$s���Ԇ�oK4�`�lJ��S^�T�m�拓���[�_/��5��[�KH��a��ĘD=Rx@���()S4��T:3R�-�)$*� Ć�}@m�o&�s|��ۉ�`ZI�C�������t��1�G��k�v�{!��'R�{�}���U9O�S���J6��wx=-6��B^�5%�~��We��s���-�� �Jq�6'�N����p����&������)�etpFM*�w�v7���#�p� ��v�*ӕ�.^b��߁JզC��d���gY��uҩ�n�"�R8M	��&K?.Ai�����=%
�b a̰iZ")��H��`�M%�x].�0�Y]:�@� �TTW�_��5��ݑ1�NL7�R�Mbb����_c����d���{��u&6Hʛ��	�� ʞ.��j�Ր��j���{�m�Y:x� ;���O�ΖEEN��9-�K�A�:4*ۮ� .@ѿNV�&�U*GG4+��3��H�a�ұC���CVz���ף��"�g=	�[4.����j��QsB]Y���%���F���h�u�V�UAR5�e�>����v�~\:#B���s��ɶT����Ġ}��o�6�8=��vص�u�!�\�|HӰ���=���:�� \�ۿ�{��Lx���\��?�� ��̷��-�,||�_�ٍ{g�~���~��Iz�ޡYtgϝs/���R.��i?׺� W!�\�V����Y�C2��˝�����c;q`�~����z�o$p�̩�k����>`<�v�	��%�Z��055͂ �vu}A�f����W���s%eU2�:/���6�Xg������J�v���d�]��"�1U$�L��+ >��yJ��t6��J��Dݱ2\��βp�����Iۓ�������T��D�i�ƬA�2j������o���^q���[9,�9 wʥ��|m�^��b�;b�������:1�ѬA&*1���cdfeYDo׽�[_ߐ4���ik���Vq?�4єT���D�d�Ux�\�Ϲ��=qj�Z��E-�i���f�U!߫�u��w�s�:��.��7�ຠtyD��]�x��R���'��?��De@�bb+����?����v��Դ;��
�o�A��T�����r��b�-���	�*���㻆A�5��ޏǰ��X�)K��v178<�E_��&0*�`�L����-�d)Bۼ��	�&, !��ȟə��p^'OI.{���i$�T�F[̱&�!�vוN���p�`L�;)�f���;G)X�(��Fs|��&��̔�~��譻�Z�����x�j�ӳ�����u�@��h�;����?���4Ǻ�j��u��y<b~6�Y��;�����s�?�1@o!�/��p~�q�N�:�ձ�"�s�`�9��`� ��~��ΰn@�ǽ�V��%���sgX��"ה����{���1���}�>p84A��F"dHL�*���H+��s$I��M57U �nċ�+�z��pph�����3�Z�r�Q���'�8mi(l8�FT'b��N$��z3@k������투m"� &>'�*��m�Lv�����x��Dr�N��-�@��2�A�Ů��m�ߣu%l��XÔ��c�'WƩ�c!F�ݰ �O�D�+�PAG
�%۵�4J�KT�5�,��C�.��2ޤw��;�j��sǜ�퐽f9�V�ΝC��:qX�k�l3}�0���J<��c�՗ꃳ��c�=���#z��nu}=��w(��9k�)N��+�� �2+�yM��ܫ�<Ώ���3�Pؓ܍�w�=M?Yk�8�YJ�&��Mۤ2��� ��tJ�Ax��=�ll�k��,�SO�
��2����9 Mċ�>�I,6���!�3C������k%�V�����i�-RD�@�ʜ���).b��f����ޏ�c���WT��2�G��	MM���:l�AaG^�zZUO.j��x�>���N���������_knzc�%�0�0@��V�		}��@Pol̟S'���d��B�(g���D���ɩ�!��5�A�w�����,�N%K�̞1�;��$��Nܗ�{��C���N�/���Ҁ�1A�
A}355#%����ʴk�/Z�����O|������ܗ��e�H[a�cCE��@D[D���R꜓�b�_�ai������W�W���߸w�}�M�vY�==;���_t�g��T
�Pha�G�_�����%ꮀ딥��91�k*�g�*k!����{�7�{_y����}�` c��E�	�Z+�NK�pn�]���� �
g��^p!o�����y�]�r����B �C�{=Y�X^ə����8R1�k��	�&\���a���`��0������� �Ke����`-���jd�#^T��ݑSC�7��3}��;pk�{W]��l�<�K:��lf���^'b�Xr�Yr�O�3};
���\C�(����c�CS#��Ddu'G�����a굉�:_�\��E�߳g��5�eZ鍟��]�`�_�%�����(���+�/T�%����DҰ����ΰ��I�Y�w+���qO�OVU�fƪ�bO�$�C�Et�"_�I��<S�!�0��� �����o=�m���}�Q���� d$=g2O�/�6�
��/,��p�;AYQ	����y���Ȕ�@Ksi��7T��$�8ğ���]5�y#j��q���dH&>���7;YTFNS��S-����BIG	��e�y���w,ڮ��SKz��nA�:H��3���F�	_1-@��>S��d4x}%/&��z��%*�Ђ��Q��It�TX��s���h��΍����8��zXs�2q+kN��a���D�ouM���GfU��ӧ��{1��7������R!�<l��,�Qb�n�^'
������#ݎ��0HLE��΀�Ա&�$¶�4Zz������N��A���y���葇e�`iRk��H��H)�z�4F�O�Im5�z�3Eo�:l���V�c���U�+l�}6ymgz$U,���wz����:��z�c�����-�єH4�*��zA	��xn!b{�0,6���ȹ�3��(|l�} Z���@ ��奆a�	ID`/	�!�E�9�Yܐ��ʜ�pfb8uR"H��K*�7�#q�MQ��d��i����t���z�v�ܳ��s$��2m!S[��2	p�3-nt,8�$"�D���,P�H��R�1�c�a���@�_{�$�E?�o���;僈uh��}��D�����>Q������/q��YO(Hq�9̋�R�(r�(��g��qO��,���oRX�RM��nm �C3nnl��$�T:�r��j���(��/��=?�,	_F��T8�ѐ� w�p���W�K�H�p�M?ø(��pz���V0��b=#k1`)9�	�<�(yb�5�Rn�Д�`�| �ǁ�V`�&e��$t|�K)�K���KFc�L�ӣ�R��S�����(/>==�f�N���1:�H/�0`���i�f��I͕t��a� ����Dj��`�H+H��x��p�IR�D4�<�gއ{	�Zb��hˢ�ߥ�S�?8�S!W�D1�DU��董��}�G[Ϫ��M7���C�ȱɬw*�9%m#�٠���a�pH�M�@=�gOai}aN����Q��q�gd�5�[��}�{*��i^Fz-:�@+���A~|�go�w�>6E�*%j��}ܿ�@e�1���a��p�p�Gd��a��x�c�|�c���Cc�3TJ�3�T�]�ScP�^__uF���\UdQU�T�}�_x+
�P��k�������>�⬀+����~���@�*!���)�+��ݩ84H���)S�H!�Aud�"5�7hT\1��͉A���w����ja�j���Z4�{Y,���G��\D������r�v=ߠ0��R�@o��8�#9�M�0�-�=��-q�6o��y���p��6K����m��&	��PzA�R��s6��ﾦݫ�W�1�����3x�6��dP�UhV����+59$Mw��{�~��pIHՐ�5v�E#
���=� D��[���Fz#D�2I!=�B���D!������gn��M90Ή�r*琵����ǹI�A�j��`�a��Y9g gQ�����^�ߔ_HVe���sRQ�ڱF4V�5:�H�oi.V�dU[ 4P�Lx-@iPJ��у��C3��P���r&ŵH�u�%*�eb�J�gZAUT�fA�G��P$U�/4�&����+�`��$B9�Ǣ���G��<�9P���VH�P�on���}�v�]�͟�#6�MY8hc�
�?�p��X���e��m��s5UR1��:E���]�ҨTH-��@X�="���&s��eo��i��4�z�}ꓟt>t���3($�����/ B��H���K%��?���Xd3����glw���9�Md�\9n[��*��l�8��F�D-�aJ��@m� ��`��(��,�t�F	���:y����qF�B���M��ҕHQ�R����ə�d�b��
y��6�,{N����p�˸��~G�"��<��;�b����UĊ�o:�-751��x}H��F@ih��O�Nbu84Hբ�����yO�O�e�z8p�_~�e���Ƿ��wz=���L�p�Ю� ����R����۟�q6�2�R��Mu�U�$.��]���'NMӀ��[�a�J�Zځ�Ͷ�x�s[O�!��
���7eVb]*�X1�4W��E6�꜇Ceª��i�@�܈���<A
�L �1y���>������O��O\t7��,^�����fhA��J�-���"h�i�Â�9ܘX��[][u#m!���J��֭Z�O�Ԉ`����������׌�w	ٗƬTc����V�&F�.u����xa���&h���"&Ur�h�BY�.5�D�.���`��0�2�sF�R���VK�)6��K�j�����~B�M�ӌ���w06�������>Dj�si:TW���B���D*�a;//Ǣ8���TL}��b�k��D���E�w�>n<'Nw���$+���ښ��9��c\���+��z�ɏ��7���Hl��įS�d�L�/�})/6����m���i�D�A���ǀ �1b~�楺�'��jkУ����6���k*
w��TT&Q~�H�s)�����j
���tD벫M2�H�ٮT��@��C�>�T*��p��zH6�y%�F(���q����^[�o'���0�[�3F���<B
��?�c���7�.�3<������w�w��KUfK�"&�
�=�ĉ\'6gw����,�K�_۫�#Ƀ���S%M�Ҁ�=�~���g|&�A��e��[t���{9��,�t��JCK�\��Ya�∝:)~�w�r����7����T0�>!�a�@|�������YF|����~h3�8H�
/l �ᛕ4V��	��bÀgoKs~��
���+6�9���B�����}>��O��=Ffe.fp�	 ^����-�F���2>3��t%Dh�gFT����o��*��-c��N
/�a^)��}�Xn_ZY�#J��"&��#5�G�2�k�9����@�4����e�R����Y�̀"�����Dn�X~����E<���	c��]~�)��yI�}"[@g`�1/l�?u�]�/ܮʊ�@M�D�/D/�6W=��EB9�|[n�r�6@.d�2A�8��ɉI�aT�f}�Q��~����M����n�;�o7H��u���b���"/�G�M �����1l�@��/���;uڥ\�qfv�VU��P�'�,�R�DPg)�6�¸�c��C�`���A���
BnǙ�L��I����Q:iD��jć��\ݰT(:�\��6��L�Hl;s���G\.��B�j�7�s"hi�uJ[tG�=�b������r_������l��ь�Ȉ�?qv
~�G>�a���t`oGr�T�2W�M��S�sÎA�f����{e���gG�D�k[2�&�,����qϝ��'��!�Vm�hݜ1��k�`
�Z�\8K���PC|FI�S��6��,*7�(sJ{3~e�Y��M�ƞâB�Ä�b(�P���ٰ�@P��0v33�~�Y���j�H�a��[nfz���;K�<�����<��K�t79坚�{�� �����"<%��ը����FqA#"M�z�P-���!r�J�R�=�E�.B�$�#F���MJ�9	B�dc$|�U���^Ԙ�+����<��V#6�vd��a
ق��yq����C�0�?y�5�S�}{�q>!�.�mF�pԥ�������k�9I�&991l�;m~'eN�M����#t~��,��s�׮]�s|^����4}��H��I":�T���ύΐ���TPO+��a�����\(�1�P`��\�"���ĵ�D�-	$�
͈�ɭФ"R���v{Ln���t��h<1�KMi
�:[g�#1f&T)��RW�t��I+�(�f�*G(�\d�[��e�9Ip�̮W�3�o��l��n^}Z�&A�䚱�hu��[����fF!�`W>��ۇ>�����?���~��Q��"���3����N����?����:J�nFi-!t�(��@Y��V\��s����d�y�	Y2���.���a���Ix��|S�ߚ� :y����{�SF�b�(�y��u�V<W945�u0o`�+�4���QT�ђ��9S�&@s�#��oO*�jk�`��i5�;�c�6K}�a��n�,��J�6tY�d:'-���c�X֢�277���nmŏ5"b�<%KP.ŽI��{Gk��V�e�i�#D�����_%I;���/AT�E��\����\u��~���� �ۉ�����SUKM*gKr�����P ���lo}����t�Dc�yP�ޘ�����x'�ي@�ۇ���Ž����p���H�&0I2`"r �:=��vυm-�6(zW�P��3�΍evz��iD�H>�?9���U6?�u\��J��a<�#�~���Y}��|�s��E7?��k(�Tn���f3b$&Qi+�>����[3��lP�ٛ���H0ΰ	��YdI�t�,�F�}���������F��q����.��Ij�(U�?�WRW	ݕR��E�&	�I�TI@o���lr�k��a<��Vvº|�s�����C��1<��\ʖ�9�jϡ�L���
bNA��j���Ӊ����K���K��I�VZ���l����_��?��Ò2��>r�k�~뷽S?���4�e&��l�bf�n�hZ� W�m�hf��}�>��e#U�W*	�}!b�����mw���m�a�Ee�5��H�`���۷������FL��;)�Q���9C����J�.��^m����K��ՐK�V�	~������O?�>�p�u��;��;d�c�������}QU%�����~���Y����˗��ry�y�ƑxKO[��ɩQ73;�xF"_��Y�iM-����f�E|�h;�Cme�t��w�R�9u���4�W+82eE�*&��N�&rqjVAX�Z�������*�P�r3#s+NJ3M���y���7�褎&���~+��؄�����H��KR� ~�pe�"�D(J����0���QX����v�@�@I���j@� Y��WX*���E����=��'� �GZ��͵W��Q6���̵����(��8j΢��q�8�'+4��d��o�΢�]��������A�J����������Aޗ2kbǆp�*�N�\xd7��h]mH�u��(]��lh���(�L�������\l��7}{�n�+G���RM����Re>s���l�jL�@I����.Q�
��WeaĦVCn�;�^�����H� ���ŕ��wO��S����t�@���v(���jk��0��9���a瘓��;���G�|�����X���� 路V���H�k9�����'L.���7�5Xslz�ذA�o��y���[�D��i�u��ʳ_���Ϙ45�2�j�@Gc�&ʊc�c��|<ӧ��<v�1W��J�l�Ჾ1��Ͳ���e��_3-/�j#:,�u76>J�gv�G~�8<ҋE���X�[rc߼�A4�"�
9���su4>i��zsА+��a�T�h�}wc�:���@��˾��K���tJ�9�g8vzߏ�߯ƜN��@����t��TKS<4������u��s�e�1TµU;Ɉ�V����� Վ���p0�=˨���S��u@�O?�:��#���_��%�4$�#u��7R�%��?�<�R\�g �E*�An�:&����2�Ð��Vٽ�݃�1�)���]�͗�Zr���=8k赅oG*׳���="���C5�ϓ�$���,�K\K(�����i8$�U<m�{�]���
"?\����Se�����n���:��<KE�
i#����sg/0��=Z�(�
��ȼ���B�����wb>�5��9>-mc��i��*A��_�m�����5V5{���LK���� ��2�R��䒚2@�y�����'��M=X�1!5�a�m�}��}�uY�Ğ��!�*b�50�Z�m\�8����A�� 5x;oOM��!�b���/�syi9� "�^ZZ�c����6�4qS������E7���g�W���E�P��P㝡&R�	`��ν����.)~>ͦ!k��^`���)+��$rj
k{K|k�X������4�����Q��4�2�4�e!�!]��-w0߯T��v�5YGD�p�����?��?� ?��#䥴Z�am�2!r>*���H@ML#�0p ���o�&�DT~Xk��N��_��_���ŋA�zY��q����:[w�Tv߾������X/���wVg��ҷ���܅�����m�WK����`2|mD�nr�,E=(?&Hb��8��e\��@��iI��3¦9�ks��ع�k�"Ҧ��k�"���K�y.]}��w�E���%��m�V�]�P�R��ϗ���|�I$��Q?g���e����B*m��-  ��p`��*5=�����#�|�] ���czz2�uJ�G�J*"Ԗ6��c8�ukǽ�/*�bBC�4SQ�~%��j�E/�JS���+�OB(,�3�YN�$�4&�o$����,	Z\b��0��+T��$z��G?��7��� J�H�Y!!��L�^O�bGn��p~���^h�`ヅpS�n'N�G�k2�-���^�~�\pS��F�=�6�%���n�E�.�M�#�H	gEXW\TyP��aх���������wI�׆�$���c��F2L*$I��\{�`��E�ߑ~^0<V�c��8]QD�ӣ���ñEe���C� /���
�2�.6��[S�%�{�1�������EPRR ȘpQQ���u�ޤ�_��G��8R��s�Yn��U ��ܬϒ�5��-{7�/1g�b�^V\��!q���4?��c�T?������L��5��	��y��İ�T�c�5>�gʍv���]vK�+nH��<mi(��.H�s�[�ńX�0�U����T3��Ú��aAK�6�h* �,�Xs���aվ#�^oץ_�j�0��V�����68��Q6D��1�����/�KD"E UDL�����e�$T}"�"��J�H��B�ek���:�S�[I?�3�������uh��H��p��g�<!c��L��H��R�Q��Y�ʛ�����q�tjb#��>�V=�OY�!݄I@��(ښ!f��))[D[)]K1� �Kj�u3��R�s[&z�c'���r����}�e+��SWQ�h�އ�uW�^��cm�z��Z|�B9%E���G]q$m�J��f�(�ȥT7���=w7=��z֨ע�ˀ����V��JA)m1
���!�F���r)=�\C yuT|Aaye�Zp��$8	����6G���kw� �[��,��߁Ѐ|n���l����Μi����9�*Ϛ�B���#���W����T�vh~^9 �VKE�ઊq������a@��*�TM~��iqX�V��c�7ގ�󎎚�dR%F��*_�.�aL�A��0�JM�=�Rd�l���R�fm?�W���d�1b��2c��j�8Y8\�֡�kM�s��G�L>�מ��$�\���ƈP)�
H���y��ZDi�SWaA��eX�|��tJ��B������ޢ3��i��5#�cn���
���9~��V�AE�@���m�kgV��s�X�����<O��RB��xk��8���jK{&�CYm��������@L7��7�}����J�5�������R�me�f0c�0Dk�O���cd ����X�*�pSʦ�M]h(���ʯ?�����*�fF���\t�%���uX�o��f�88�:J�*�9
5ʵS�Շ	Տ�%�aѕ��i���Q�)h'e�Nȴ�?D�8�?�8B����ZpR��F�:���'.��*2M�S}Xݩ�?jؗ��1��K������L&�(�?�V�� 1��1�W��[喷;n嵻y�;��c;A�t��N���2�8H�X "*�U�"?N8�����9	G	����%򀮏?N�&�LA(�4\�gm��F�#��bJ�#L{a�w@ew�}�Vѳ,ԏ�M����3�b?2%%[�C̙i~�VhO�|n����@
��4�pN�q�qc�2c�u.J���P-k®���9�FӲ1nK2h_�����7]L�h}�ꩢrB�A�Z)OO���T�n�nvМ�L���m�����������d�մ���=���*چ M��xc�&kR�w�R�Z}^��ի�Y�g���)�%�P�3����d�y�Wk+��V�e����"h��uEa�hqS�"8�N[��[A���qOZ�aг��Z���Ŋ�~/�5qX�f���im�	J�MwP�[N�n��m���J���k��5>�IXo�ʰ�i2Fy)$d�
���1!S�kG�H,=X�mI�\�v�-/��hv��J%2�R:iv��HB)�;�:[pb���=g�_s0£E��gi�VF3��{�1�w�}&��AE6+[��#�V:9�4ؤ�+6�i 6܃�Q5P0��d�M�"n�(_W�w�9-�gzɎ��9����O��XG9]B��FY7��E��2iQ�PQ�U!��j:�ϒhx��$�O|������c:�7fH`�ۿ�[HѲup������8�?mi������@%�m5.�S(��Em}��aUV1�t�b�)��P7��v�kFZ�<��<IN�}�tgϽ���%{����)A7z�4`��!�H�5\^�:
Q�t�\��R4�'E�h�NT,�lj�D�� �e�k�T�*q����
�y:��S����� 2����O(f�d�)�y���nm}ս�������ݷ��&+r-�T(��E�x[�K��������\��O�!Rػ�����i����)���l5c�ر�C�L9~}k�#s� �Zо����X�Y�e��qϑ���h*�����&i�Pd�sn�q���yx?Q�(�S;tlJ�q�4���3�$�Ǳ�&p]�|�I���jK<D@�$����Pr��y*ȇ�1�>81�Q�,|�fO8(k�pq�ۜH�ȝG����Ӧ�����d���Z�97Q���2�qP6��I:�1l��*m �J�g\��r�����F��0�7`���
{������n��|�!�+���	*;�!�v�僆ؤAE:g��%(�X���[L��ퟣ�W������z�G�C0G�����(��T�����o��Dd�|�Y�X`}� 9�ʮšQ��ҩ� B��~���_#h����6�H�H�!�����DD�[�m�/�Ҽ"�[�v���8���C�y*�:�?�Un�j'0�)�P-���17:n����Jg�c'�v��i�gC�FdPwi[p㒚�MX�Pu�Nh��=�^��eKNk�,J�8 ���]}?�'����}@d�gF��������^y�U*���?���t���(�!�m�6Ie�h[���>i}���5��{����z.�w0��6�����}���͜yK�3��m�\6@����)���� ��1����VpW��&����`l25S��-�3�o)�z�q��UƉ��8<�f��+�w��{�0��9G���̡i��U S}:"bl&��0�����'����qϿw���f�J(Dn�>���"I�+C��[\V;�j36��Љ���k8:�RqbjO9��A�Z�T>��$�	W��G�D�@�P���<��:�U#d�;1�C�Q�%������d���v%�5��$����#޴�8��ı�fAu�O<p�������+��L�[�J㷠A,�{sԔ2o��	���NJ���Ĥ�����۲����ѻ��e�<��%�؋�����K)B�}��O����=Ci��y{Qe�*2gV�A��|����5�5�����*I�|����' 7K�W����~�i�A��P�1˪�$�JC�2Rm��M\�~q������99�C�t�	Ъ�մ*��M����^���V��}A�Z-�����G8b��p�I�����6�Murac��� Xd�:c@��4����/��/�/��J3(�<��?�,"(i�?򑏸_��_wgΜ���l <V9��i�lh@Q�sNQ;�s����Ʃ���en[ە���G;9�(b�v0@lKƥ;�	i�����=էe|E�w�SE��w#�Je�f��L�hN��A��T�c�d��+���97_Y_�����y��\�
�V�P5��Ј]�E�8,�f�
|s�⨠t��E�Ҥ�M��tJ���]\X�糇���K�X���!�9"�ЅJ&��"ʘ���F�j�⍽9����������9�+�TA�v;�$DBea��r���K�K�K��7�����7�eXUO/^�G���� .�C��Q�uǦ�}6���qX:s��9�����qcA���#"a��əK�]�.���T`ޡE6�$"�f�u�N�-�bD{�Q�j���aS�����D���LǼ��Lu�<y��lvv�׃�'&'��Q['�,�*J��c Dt;s`�qL�����A��p���N�>�Ν=�z�~w�z�]��FG�n��^v6��G��x�؜ҟ+v�����F��2�%�yt�aІ�ޤ�{=�4���=%iT�s��]ڪꋳ���T�<�F�9S���x篃�խ:��k�Z��"��RH�s�}�;����� ��0?;]759����˶)H�B��ߐ=8w�k���E�ج�_�ܯ�ٙY�P*좽�rhv��0�;�������ٰ%a�T���&�
��k�Y�ZP��Ǯ���&vs�)�膬qc1�_H�D9�?=��G5Y���Z��)0����Tlϼm�8K#�r�ܷ�z�}un�~1nQ,�ρ��^~wTJT��)w��!��T8�ot��c�KDٱ�jsA!������0U^5�TA��o��BF�$��9���r�
�ұN�Zq�˛%��ȸ!Z蛩N�uC(�qqf��$����˗�:������+Z�p�iV�d��m�P��h�Zzi����6B��7�R0�������?��`e\'��M5e9�{��z5��
����11j��$�@�/�����D����$��)/�#�q�9�66������&�};���ϔ+~ ycR�3�uj����k���?na{0���x4�O�87�,�Rӹ����ƺ������O��yԭ,�pW����Ĵk�wy�K]�qZ״C�c��G-��������X��
l�e��+��
J��m}p�&�8hje�2t�I[��-1.��N�Տ����`�[t@�����f%A;�.K�P�% b{�y�O�u���o�g��{��Y"Q��w�~��s����;v�;z���Y0�&��x�!�r��/XWqk�80�҆4��R��4�vrlo��^X��x'�+�pAGq}s�%��;q�K�˅�������������O��u��{X~�i~��|�`dh�A{I���Oh~7�d;�w"�����;����}�	�UL�N�8�~�W�������Q'��_��Ϻ�{�`Th��Z�bS���͞+G$�>�Q9D��K���j'ʼ��&g@"
)@�*/sV��fK��,��Ė+e5���p�P|XqB��+g̹�s,�J�{l�B�;�_�N��
�oߐ�D���cKK�ܙsn��#�#���+�Wh܎9J]�/p�� P��c�S3� m�n�U�&�s���ZiI���i��p����m8VV���h)(�����cw�Z4pj�Ai�%Zp�,�cH�A��-��]H��b�#b���(D�._����V������sB3ׇz�]�O�}��*3��Bd��av�܅{t�)��,�>�I��DL�#�ܐ���h|tҭ�{s�ڲ�1��F�c�Y�u��,48�z�C�R�L�qK�T�-��[m�r�j��Q�ǘM)}1����+�¥v����Z+w��5�\�=$a�����[\Z��'n��n���4���I�����,8?O{g�����o��� ������~���ܦw�_?����?�C��㏉��u��|8�3Sb�
�@"�}τfq�]��vIU�Y���ȖDNO<k��'���ا�EU�T��u*���Bڕ}�|౉k7g����qϑ�ծ�$�l�8,���cǎ�0Ԧ�d�y����JP�f��b�a��Q݁��ڪ�r�J��:W+k�v`����XRR�@�Xc���'ƑM����(r���y_�خ\��<����Kչ����LVW�u
G�E�Xc���M��6�k�����f��m|��B���E��N���E�@��_��p��AX�#��ɟ������c4J(���0�di��wx�6ix�9-\�t��#@D�k�הp�^z��������ݤ�� _�Âpx��M�"8�p���5<B㟪�
z5չ$!�!/L+��`�z�-:��� Qü��*%a'HVN2�s/]��5�|)�r�N��>����c9�#{D��d�f�c��K/�ǟx�����%w�;��� M{��ӘFhY|��}? 3�����m�א8A��=��a���?~\�CI*m-
%��ʬ*���yJ��c�;�s���x/��SS:��&��{��E��7��]�����J�:,@x/�?�~��tT��?�g��'?��hem�C	8�J�\6��[����W_u���7�=���<�Xg/
��˘�Y�:�s��a<7��<�' �p�H'I�����WrI#�~Y�͋�{�~�?k�	՜#���gˏ�Zh\���&xuW��?+&<T�M3:�ǐ~ ���nu������3��3}�� �Y=����|�M�O��O/D��<��d�`,�Ώ��lB�Gpl�.&bm��K9���TA�B�!�5%
��Ԡы���5<ߐRנ�xC���J��L�\{�@� �]���.^���:̔�p&�� A�4NL�)�[�
�ƫ��m!��<�)���`�u��i�2"U(Kʷ%��7��[�ˋ~|�h���<���Y?f��{���wz���< �x��:�.2�F�ϵN�#Դ���b)ɞi+<[�E7np���%�j�䛮��	��vgf�TYZ��%E8�BW��l��a���Rt�~䑇��?{Ž������O�{:햗ܥ��?6����?�PBtj|�
}i�5�,����-�Ο�7�G�"���ڂ�
��U����tYY�έ��!�t��u�����)^�`@d�L"%�9���N��QU��3�p����(��7R]뭻o~�������/��U�i��c*To��\�s��~�����'I���q�E�T�����7����^{�6����}E}��Pt �T�N�4oP	�ܒb�B��~�©�;Q��0�M,,ǆy�M7>6�	��v�}7���.&D�S~� ��׏���n��X�C/�v�쫯��{�dMLZ)�+mI��2���g���o�����>��:D���G��:�_�ī¦�s�����uB�푌m��⧉��V����̘6@A@��h�#^4h���"���e�h�X�۫,St;-�1���t�4F��6�>�M�Ν�ov�w�r!�=z�>�]Q�$m6�Y����7lH���s���f�6�K . Lw�D�0�>�����s٭��u��i7��H�G�S��w#�g�8��B>ל�J�.�8�w���aDy�˪{��[��0e���$�?� f��{�1��/|�<#�7�x?/G��R���f'1���{���ܫ?}�ےkމ9��]�;R�n/�k�\o���31CԱa� �B��Qm���LB�^�dȚ)+����*�J��(���Uz��_('�sL��Wo�+
p�R:4pf�h�Lu�;��ha���s�>Kg�PD۫�B���o����?}ǽ��)w;������p�����+��W_u�++�n� ���I,88��5�n�I������|�i;��	W��3�=�3�V����"q�}rkv��[<i�a|�B��J� @�6oL>�eY�*�0�p��ܰaW���pB9������wy�.����l�ׄ�J(ũ���g�Y�!��ayX\Z�� `�K~����wOq�>��O�� ��s�,�\`t1���t�G�>z]DՄ7^s��2�ED�yl�����$�#HR"�b@�+�Q.�"�Xl�^��[٬EZ. 0M�>�'��_Y����3�98Z��8�es�$*���&#y�4׮-���UJ] o�=��
��6������wgc�y��B�~��裏�/~�7��+}�dn=��/s����Iw����ۢ�K���xK��(�ECKhX������cl���$}�d�I+�1"����J�5V]�9�g'g������~n�T3�c���� �����G?�~�W>O�ך�W~ۣ�2��!a;���"�x�T�f����f�-�ҀO>�	rE����Ǽ�3K���WT��C���d�)j�(W�.m�4Z�Յ����Y��U/0.ư)����q���9��=>��+�!�l��Nš���yh����wS�DQ@v�|�:?�|+��w���~���,� �GcX����`��T�!%��K/1io��� )aVi0��5��S��8|G��̩jܪ 3q[�{�ډaiJ9qz������;|b�ҸjŰ~��r�3���:2��iM��A�������V�d �&G�7F0�?jH���X��*�y25�B�Q�e.T%	g�Emӌi���G\�`������#�8��T'.�;"*�覍���	�r�60�O<�y8��7�3���0v�"�����"s+��ܬ0��c~��(-`3^!g"m�Jusw�Z�� #7�k�e�������/~�uͶ�����{���w�Ue���?��y ���@xD)'�}H)��_a:	�&R%0��|��+i�\�*0f0v�N�tX[�-evp�U�RNÎ&�m�c%�H�����0�/8����xljj�=���o������:@�㇏����� �?w޽��[t�1G�ۂ!(xꩧ�:l��D<|8;��
�D�ґ~�z(�>}��|�N���l�#����c8���X�C�>���
nv_��2&����l��p�h�p�����o8��=����~��;w��uzj�;��}�t�|)�&�gt5���C&�O��T}ٜ�u�N�{��1�sA�'\����1W�M(�0��J�H)W&�OUj�ܾ�)s8.	k�Nο���w��Q�t��9r?{�Y��5?�-ɭ#m� i'�-U�i�`�
j:-#������f�4>G�o�=op=-��E�� �&��.���z�nF�5�Y��i�fmw�}\
�`�UM��	�4���s�S��*��8�͈����.,R֒[GI4�Cj��D���-z�lu$�N)Y���n4i�S'�	��q��%�C����,��j���d?�}��pD�$�*�ϡd��N�zB�eS��W��gg��v�Eb,�.^\���w��s�3�����*�S1��\��"�T�O��7J�+ǧ1�΅R��,���E�oRǿ��*Z�`qlp���՚�|�����l���E�0�4e�0�V��e���Ж���k�mH?���T��{��烘��	��o8
�G/ !��_�|x���D�G�U�{8��c?�Ϻ���q��3~���SS{8߀��Y���S��A|�+_�
�I�v���z���X�N��y��;�DC�`(�@Dl��]�����hV]5f�Z��q���� bK���Q��pL{��~�Ϲ��~Ý=s�=��~3�&by)��θຣ~l:s���i���p��N/�l�L�����g&��V���P�fE>aYsfj#(�W<E���"w�e>0��]���!���>J4�Q�q��Ϲu?_��D=履M�rG�J�e��L�%q;��wc+|��s|� 5��Z�6��2n��5���me��I��㞧�Z6b�����F,��X�R�6/�D��ٿ���p��Rq�����QI�Ǐ���YV� �7+9�����b�&}u� ��q��VXT�>*�v��YD�؄@Ĥ[Y^���m�YC�bzf֟����T���&>��w�%A06��n0f�#��ӭ�m"ee���R��ʵ��0:�ث��x��$�gJ�����s�7��z��ri�bA��{�_�c����jN�=3,U�FZK!Fh_s�5#��� ���u�̷�q�>�,�6Gho@Ph ��i���sp}u]���Q���w�3:��AM0?֎5���Bp��3�?N�,�
�� ��k_�[k@����Ҳ8�m)& ���X�������>^���/�(�L�\����]�vo�Z��L=���@wt� ݄���2xSۄ�
����<Ga �ˡ��y����� �l��?�3��c:Bq>:1���*�	l��A�q�T��ih��*�Y$Q �AO�>szJ��"0�:�q�ח�4�DSF�B����a�t�/\��)΅V��|��!r�T4���w�3\\,9~/D0hJ�ŶM����p�Y�I'����gA�Ѿ�!&�z�)�#�۾��N�S�g��/�tsp����o��|7�{���RLV-d,q#����
�3R1���(C{�P��;:�!�� '��Y�ZIy�p�a�x�$H���!d�_�l������MG�z.9M����	ӣd��W�#D���x�C�&i��U�N��}~���uF:*�T��+�n#����h}���cQϑq	Pf�.R�(1�����a�{Ej�����C�y�]:40�@Ӑ2���{����9nޗ/��{�i��IW�)���793�<�N���7��;��'���._~���5�� >�:.���ȁH�5�(��^;�����O,
V�9e�a�(AM���M	H�����O~6G<&cP�p���đtC#=�7��l� զh��FH$����BD{�G<��Yp��U�T#d<�3m�x���|��i#_z�y��,�A�޽3�Sy��EW���'��r>��	��29���u/�� ���͂���v��t�����C���T/c[c/�Y��Deyb)K��V܅���yء�vfz�]�ׇ9t�3]�6��J��%t3��-���*�f_¡�&B��G�����f���cجގ_z��Z*� j�I��p��̋ܽ�=o�o���766j:.�˙W�Ɉ�!����^H�"�8$���l$eڕ�h�_S��k
1�XL�t��Q�o�>@�,�V�k�\�� 6qu��t��hؼ�O"�_�~ս����c�?掟8�._����3n$ب��M���n�����Դ[��
��I�D)Ƌq7�mSgќ�1ÚWC�H�)��,�j�l7vj���K����oM)E�2r���(<�DS�����wN���CNH������5�>BCs9�6@ �Ȁg�1��
8{p�Pe)�&9�f�q��?8�_��Dk��@(�N��1[�[��V�E.6��-��~]O�%�}MUf;Y?2�$]\jW۴IXMD�`�ߓ����Z[Z�y����jZaE��Ś�7��rڃA��ε�5�ޫ;u+s F�,��`�1jg%'t�(�96�{�!�F?^�����z�i�3gN�M�?c��^�_:��n_�#��'%A�U�Dj׀��i9��ki`VO|��NJ�܊�ˑ�#[�2Cn�-l~H[)"q2�6�y��N�:M"�fO�gmu�E����Ip,��6a��{{p��r�z�-^��#m����n��n��\�1;y_#�j��Ww���j�:"�S-;ᔁ#q^jM��qO�¸Y���+�����2W��n��9x^�!x#��ҿ�v��a�"yۛȽ���Ю���J��drl���(��=��.�%�Nx5[O��,Uuҥ���K�k���k�d��͡ÇY���̆cݮ�l����#ڝ�j�5V���\.���Je�&��A*���F/� *��uX�mqU�cF*���%�;�^�B�)t�-KBgN>GϽs�{��W(�1���?��xf�;0o��&yG�� uZKi2�N-
�FA<RUԔh�5=�a�̽2ۀ�w��2�}1F��)�ڇ
�wfb�ӑ��;̣VVjUb��ؘ�6R��=ׂ*�.S���Ҏ���qO�< ]��ۅgP`mQ�+����ݮ$U>�zVQ��*C�u���JAӁ��
�@�o7���mX�Ҕ�}N�V�=�N��.�ap^�Fǉ6 �
n�? W�&L)�ӟ�v�<I���7�X?����ӋK˼�(�X^]�9?��V	֘[�y��ҕ�Iq��[m�!HUQ'�Z>�2��i���ه�ڝ��y)ixL���ݥ����N�Q�����%�Ɂ��ޙYꨰ-JRyA��w���ع�����:��ӭoV���Dv�4C�Ds����.ˣ6�؛ڼ����}(�m:6��R�op:5P�m��懣�B�馲����#�އ㞦�lq�RJE-r�����L�^�:ȀȇR\^f9���zHņ)1��`�a����%c�o�P��%Y�������Ml"�յ��aQZ� XEui��͗/�����w�>L���gϻ�ǏS�M5�d�MJ������r�	�~}�N������ Q6���{pBP�*�%��{v�h-�N��.��[�������T�ne��WL L�g ~^_� Q��wh@x��(�Q�p��S,.���|�=��O�{��s�w�fD���5ONBչ� m�8����F��yPn�x��~U�g�(u�����뮿�nFX��E�6�z�`ﬤJ5T�LCp/S��W�iߛ��1i����c,��T�漍Oc�=i:5��͔A�>߂#�<bt��ӾCv�TU��P@'��J5���ǻtt`3a.��$X���>�~��#�W��=~����g�;�7��r�k�x��ڵ$m"����T�z�I�����	b��#��fW/���08>a>@�Br�/#�����m;�lH�B}�m��>C�u��~rm�_���V7�=q�M�M�Ay����@g����t|�a�ԙ3���-���v���BK���Um�U�u�GL�F��ﰢ�N����ȶ��':*D��-C@e]<��֦�>b|µ������l��1�k*����=���5�F 6It��4���1���il���Ō�ak��|���,�Ne)ܨ���i��6*�؀�#	F�V��`���#/��w��NO32�*%�|����Rf���@k�}�Yv������9�1�>��-UT)Eʰ���.IUq����f�w?��Ȅ�vXB.�N±�H��]%��d�]A�ԩ	N���T��`7ц���*��&�7�L�^�t��9^���:������;�ע�e���6phZ�w�ܙаU1�Z)��G��q���W�m rپ�僒~�Id��q�O�ᲆ#u��wNjLSh�Π"/V��O���U��w�k�g��|�#I��9���3�ۭ�5Cϳ�~����(�����<ѳ�F�n	7)����O����?qgΟ����3 �wUG����)u�ctf�Μ��ٓ������|dc�
Ħ�����h���R�1ShUU��Rǁ���Y(x �b �8o�Y�����ө}�ч�Ύ�`,l��ǂM!!�T4��7�$�#FŚAI�x��m|Mx>��T�J`�Ec�LD��?��T�����N�z->'ZK��a��!�m����o��?mN���p��H)|1�U����=Ejp gk��XG(��&V�α�M�k�;��h��hqld��x:�$U3�p.��$�*���̑�b��o��n` �����V�7,=��5���n�w|İ5�������ܓO>����A�,�	N�HDg�����NR��)@ٽ�:%r�Hc�Ot�ؠo��ON?��[ Xj���*�/�B�c�H�@I���Kuf�y�؇aB��K7�g��;���8!@n���w�<�(�:8840p��Bc: �c|�y ±���a_��ל�a���ӱ�Y��<|�'���X�$lP�㷴D�\�q tF����E�	���N�&�+���$URpc�:EF��T�n�V`x�A�����WH��t���ʱ��Elrb�;���@�|�5#ܨ��k>��Y�_^��$Y�ak6I���pl�BzS�/@Q��J~�.�X�H&�ÀT
66��)��gY՘� i�n<��2^��qӦA�:�mA�^�w7 "��`��z��;��ljU%�<����#��E�/�t�R�X�i��[thn��;�A(�@�JkO#�C�K\��DaLl����a�qhj��� 7��`Rꀅ<29��k��&x�#b�o?H3!����8��A'�H�q��f�)>/��&�/�FSJ�ɧ;��li�KK����y��ōE�RE 7x�6����a�\�J�X����T� ώTܚ�dD�5HEML�V�eaLJÖK%��Oۉ�9)��;�JT&cS��j)�ҚTRu����7n�7����D�3�Z����.���/�kWo�|�=p�!716I]��o���H�� �s�����)F�~�;���pS"$Ĝ�xsL��7�N�9^s��w��~�ܢ�v�;���l��!����Z�g=ɰIC�|��_~�s��T�q`�Î��5{��q"g΁G�+#�����#��ߠF��J����i�v�I�iy��R�杘T~��g�K���^����ቤР'''n�S8?A��Ho�4p�Ёi#�S:x���)��8�?�\��9�Y���T\�'��c�D]��]͛^g.Rv�H�*A~;�>�w�(m�/��<, /X�[e/�x}T'��
�g�85� ۡ57;�[T����д�/XIw�0Z��u+���nb̉�=X�@�)0ua��`R�5���x��#'�9`"S�A����M��Å��8�y�a���0�&~_S�	�n5����d�q��ڻ�?����C���K�N�YQ��Ļ�� }�>쮖�z=�IKJ$($�����񶧽�g��q*���j3�=�tlNwձi"߈x#"��������+�s����W],Zׄ�,��Ҳ���E�*JtKQ%I��s��o|7<4`�v�!��)���kl�l�*��f����n�S0��ٺ��V=�$Ǣ,B�+�eI�&�{w!��
)�o��4Ǐ�4��}Z|�|����02�S +�Ks��9rD
f�� ���	0A��v�@�v���Lk�f�:V�o����aY���|.���:Ӧ�&�~J�Z}Y�8�:P�v��(u˘�oY��.{���ܱ�w��,5c��X�8��� �;p�>f�l�]�͍k�fbl�80c�s���yi�L�OH ���.m墣
�e� �?ÝH"If[�:r��k>h ʅ���Zw
K�g���!y���$k�sG�*��q?��M���~睇,X;"��s��yxh�_��;�9������ƒK��`��eMO���u�dn8��^/���d.t儬�w����qX�,=�E���̽�Fg�ɛ�Z�̭ܥ��Q[�p�S^M��ָ����Sƾ�b5��c˓�����#�����wXnB+N(��#�I�����S��Q#G��&�y0l��֛0��F�f��a���n.]�'O��w
B��\ȴ>�o_����*E"��PJ$
V�%�--�XX(��Y?}Vxr�|��N��n��#i����^#��d��I�BU�HJ\R�e�j[p�����H�9yn4!�k�����1!����:u�y��G��ܢ�p��Tl��.
hEKC�u����3�<#��>�J����/,Hb.�k��H�Y�>�$X!�I��$ܸ�jd����Kq���j\z�(u�5=/�Ѯ���jc!m�0kQz����deq:���>�%;W/�m�+�߰�𝦿@2�5�Gʣ�5�er�~`��u�Pc�ݿ��ڱc��zgg�ٿ�Y~$��c���B�A��X�Jl�e!ro�8r��U$r��e81\ų\v� �M��	~�V�y*�2��Oz���N�C�I0�dI�w�"2��+����L_ `x�דZ�[���n��f�ĵB����#�	U��8����"�,rmn�؇��Ţ͜�Ʀ��߅g�#?�Jυ��(V+8X�?�.yc��,�1Pv��c�i�'��8�d�iPEp����<5ժ`�
�������AG����I��ڪɕn�cѢ����QëరX�l&����]��eo���[ Q���(BMh�"�r�j��ea��KlN%391+�BСA��Q[%_�]r&_8�d]�hq5�ȼ������Gۡ,�|G�纬|P���ẋKes��E�N�2<pڜ8q�jl7�g����z%>�������@g�Ep��G��Λ�f��VXX�fK��oT�ҶȾ�XX�Qs��&��a��x�5I�(�d�Nq/]\��s_6��$ǋ=gKf5����9���>k 5knj��x浌YZRM_��]�U(�@z��	��;�+W�H�I��Dr���U�`~�|��v��1'���k��\�rI����%.��РXm;;�MOw�}|*�/��b��0c��s���4�` �����X򙗱�@x1J4�?�ib}�ܸ�{F+o��<�'V�ٙR�J�O�P�#�h�����340l�ׄ�����.
Ler�G_ �P�PjhMŅSM�j��99��+�8j��K��R�}��ͥ{�Z�X��3���Jͻ�,��JE���4�C;�Ċk������M�)%(�$��g�\_�96۰6�-�~��AI+�NUI�an�5����������9�I���l�������Ѫ?��`M�6
f0Q�yCĒE�j����,LI�o���,[�(���~��XaT�i��	�$e:��r�*�Ai��Ju�E��8&����6X��.�C���A �	�\N����)�#s��� �abbZ"7J�eɠ|��I1�B��z府�㓓--΋ ��9�s���|��S�����f(�l�vsjT7۶=C�}���Q��	�Dͤ`܉Xpk--��PI��[G���dGʍ�՚,[��Mֵ�A�����X���[82(%��cǎI1O,6Xh���H﵄oHc���{�>;6c�cffj�,/�����()�svӍs�V��w`�>+��s3nc.-{��%֙奥$r���	�q�Wqw��9qc%���ޱ��-̋<��;~�9�Xh:d��	��eil�l��,�tIu�gF~��Y�<���1��tH	���.#{�g�6��#։P�ٚ��q�F�)�A܆��Z�V7S���v�f͖��&cnݪ�u=�^�����xޗ�aﭹg��]W�9f{奶m�ҭ�S&��iB��n��rK���+���tWA�R�5h+�ib!a�l�18#,l�y-�� ��Έ6Cx<&]���,z��,�e��H�C{��P�]��&��W �F
V��C, �� �e4���I{/!�>��"�����Ǻ��I�R� �d����Ԍ���>��0��K\`�qy�׭��*rSt��(V( �8|�9}��hR���̰I�=�#��f�rm��YO[�ٖ����\2!�z��fSa#Ěǘ���-/K�X�J����D8�ۂ�Li�ꙣm�=i���6���}c���|I"���-���@�7�0O=�� �Y'Q�(=����:��97g,(�kyy���,����ū���c�G5��r^oO�ȅbq��T+Bݵg�\wʆ{�(=Z�E,�$�������E!b�-����1�J,5��|�)�0<���ٽK6P8������r�뮓���Ιz��
�b%��;k
X�;j��+�i�7�K��I[�����x���Z9T�R���,�U�䧃C�0��ؔ$9$�K8�E�`*YX<.'B��gf�[7��
�oe�YOK���>Al��xB0��ѣG��.����V�-�Ը�i�'�)��E�U-��_�u��4�Q�56����J�k#�jZ[�gj�ZXZ07�n�������b����@�uS���-���^7��l���4'<��w0��;�h8���N6=� ֪ya�����K� ���F��������\9�;;R����KL�T$�w� Ʌ�OJd�rxhĜ8�3������!>�k�}�E35���
��|��Q+�m�'?�IR������P�C�d�^��lu˺�	�2hu�,��8�GUb�L�h������MR7q|���_��?+���/Yc�֚�.lu�5X�6ښ��=ڤIF��.@Š�3�w�v�]�K4��9uꔬ��{N ����+V*��k�"�(�	�p�ߋe3=5g��QZ���ό�MZ���pY�A�ݽ{D��B�g��zs�F��DK�#�P��F�L�J䚺r�*_��)vt��׮�3g�H��{���d��.�g}�[=h���7\C�]���h4��u����;bub�Q��x�B�kV����x,D�>ݿ�|��ΐ�\��������ł�{�}s��yg�IZ���Y�/2Xkf����o���\3f�:f��ح4A�|r=�r�17s���#泟}�\�t���D�5��ն�82oU�2�ɐ&��Cx�M��7(,�u�V������pq�j5GgY�D��s�vR]�d)i��}���Ep=���R�{Ԃ ば��
����ĒC�]�*|��9bȌ	���wޑ$]������9,cŤu��%�"��nr�|�I^�tn*�fD[;��jQ7�`���U�OmH��B�������+��I!0s¢$�ׅT�J�@�U ��8��G,(q.Bȣ�>NrF����via�V@���Y��K cG�#�[�񺱈�%��m��_���_l��C��:��$6]�����ёp=��/��U|�~O���y��/|����?�Ϧ�e�5L>�˗/��s�������v�@�9 ���~3k����d"?}�~qQ^z��v���DI`M 7XVǬu��<����`�%�|��Ysc��ԟ� '�S,5ȝ=̐�v�<�����wV�V)����̜$�DviT��Р̥��*9dx�a}�
k����:2й��E���M�ɉ)9o������f7���	 �{?����.����9��Yq�	�Ƃ>�T�k�L�k	���i^�FZ�c"����"��%GT�{�*)�5"��ж�L�
�0�L8�r����>G%%e�`ڹ�� �Z@Fx|��v������Y�]ͯ���X��~��?q� Vp��YЯ,L�ۼ�&�'̤�y�/�}V X���aAt��礖ǁ}w�Ż/IL86:i�oN	7�[�!�R����O�32�� Ӣ �U�F5Q�.��9cJK�t.{]IIi�$�+�.�uJ�aj ^�x�LNM�5a,�ӂ#4OOMY�2@Cb�w����gW�3 ���4/QV����Z�k-��LM�lxٔm:xgq{א|�=��s .�@�ig�K�'! �9M*g��Z�Bxq.6�w�7O>��y���ec�{TH$��3far� E�SO��������F�|����2��X�{����r)�!�)�������{�h�T���)g�~,`a��=�u���¡�!�2�	��FGo���ʇ�CB6�+�{p�~�o�>���l��=VF
�� w��>ʬ�eb����L�:��h,��cy�n���.WMwg�<8d��>34�C�x��M��pD$��K����l!&|�-�s�FvH�ܙ���D��4s�l�V������� ��K8��Ҍ���d���vJn/�;�~Pq��%QIrz�*���I8w��Rf�4�\֔*���IsmVS� ���V�TZ�i���Gǥ��Yy�#��kW��7~���3}�S\�z��*[Ω�4�34K�w��s��VYZZ��p_n��6EѲP|�����s� �?3��V�ٷw���P�y�X��w�^�w�^ӿ��[Y��LK�~��.c����;�&��2K�9�ِ��
�Ŝ,R)�Yp7���ZEH~4jw��=e��(�.|�$�7E����@���PD7��Ʀ��>뎝;��dE�9�N�=o����!�����G��F�e���C�㕾O�^��c�׿�٨B5q밙�B�1�!�4_�rc�p-� ����� ᕍS\VR�����F��T�^6j�w��C p�Vm�5^;ظ�66*�r�C��={N�}��a��,�0����a�c!��u�Q4#n\:��*K�uq�-�{IȇT,%G��kׯ9�U�Kt
p�㛓0�={�5�rL�]q����7;�8-�&�9b���ćr_ ю�6��}V��ji����`�Dcm:p`� (� ���Y��Z7�&�X'�u��L��u���m_a�m_��Ns�*kCC#���I���w�Z��z�
�����e����m=�V�t�		�V�P|Sw ^Q��d�]�f�:s�|��O����d�-�(y��jj�х)����"~�m
��ζ��s��b�>&/�q��Z�ʤڹc�%���5ԛ��J܁D�;�L�L��ZDA���96.�H� #���%Y���	o'�yd�Yju�]�j���'�XPs>���A$��jh����s�/މ9�s�= ��������Ry����&M�z���r
�V�+ۍ}�q��֛v�d�&��s�ϓ>7~�ܚ�k��?A�>�G݅�q2� �h����]508 37_�u�o/���������a*��/j6�6Q�l��j��N!Zr��߀@
�Ϧ��M��	Kn��bn��n���s�tA,�(9(�%@�f%H�8�+ѕ����)��
0�xCJ�������81�v�3]�CV>�Yac��TQ�wu�$�/�}�l����}���3־���ې� @'�	9F������^��>i^��/̷~���WS��5w>"�������T��k꜠��X�<������L��k�n;/������rI� �Q\		+����@���K��m[�|/�pè'͖��3�k��o�Uh�g��*��Uh�
L�}ق
��ޟ��粹`��w�`�����A�P@��u��V�;h޳B�ƍ�y Ȩ�,��A�sYec�P@�aJV��k	@�^����9�U�^��A�?�}�L�,�Uk� C�I���G�\>�;w�RR�\T]�w�\��6���qkR2	覵��"�G�^;���Z���wl�j��\�x��H�u�ph�����-����q�9&�Ěwk!ؠd3P�ʂP���+�������(l�槒Z�[��0���]�Nɚ~뭷�2Y�pl��ʲ�Y����r�p�\�߲X<XK�ʂ�mU����7J�I�z�b��\�5]���v��&���`��Ʈ_u�(7Ku2�7��� ��w"p��vݏ�i�}ժ?ӟ+��?�P�2�SN����a�����Q�������g���=pP�9Qf�)�����R�Џ����	?J��������h��1��Y�^�v7�C�4 �f�'?O�\�9���Y5vp�������Z�[j��dP��Z�)�8��(ڒ���V��s5�+h�_���BH���k���#9�}��'Z�:$�,H�]��y��'�")!ɂ������5���	���%!��D[lb�}����}�I��O����Xi4y"@-��4�*��A����4�"�H��Q��9�U�N�{^��C`��^�}��-���[K~�t��3�Қ�wRA]�c����!�;¾�-8���F�M	�kw&p5�*Xr7�	Ӳ�\uD�|`�f]�u �2�����~�ǅ火W���VXKX��g��9��1c� SX�<��a�X�x.��Zn
M�� Bj�6�Ǻ���@����UZP��A	���)	���Q� /����͍�m!�����}a��a�_ȵ���f��*t�Y+����3o�c�8t��Y�����|�}�8�*�(����o���նY�Hm�k���}�DA��
�`bj��*��:�W��{�\Dd����Vs9ɶ��d�0�^��2��K�*�>
"<N��R�ZeJ�N�o�gZO˚p���r06S0�����p�(�F��6zG�+%�̤� ��)����dJ�DO���X`(��2�ΊPs�ϊӴ;�Ԓl����f�d)�J3�-,��;�����ǿ���HB�iݮ���6B�����i3�}?�M�V�/x���Z�q�y��m=#��Y��i�mؒ컫�kX���¹�b�,S�݈��T�1�GM�?��!�}�͒�[�Y�g`I�����y<
���RKlc��d���r$�,s��y�~F�9k<=��F污/��Cְ#߻h@�����#�MXCW�^w ���%�5��Eq]a�|8��*�sS];y�Ͻb��5d�Z���z庬k�c��&k��_�s�h�tq>φ�E�)ugr�f׺N����1q��߱(#?nX��0��¶\"7Ό��l,�?{�E����j�9jb�'�x�����l?:���o^���o�Yؔ��u�Z]QzN�Kbs��Œ������>�9�y�e��ζ-�'EͪEk$�~�-D�Y��V\��85�f	�V-}�Z6��xi ��v��G����
��
�
��Y�Y���g�u �6}��hx"�`c�aQ�?J��33SUE���E�\�ٽ�4'�J��,��A\V��/`ghh����բ�KK��:B���?ό��&5�|=��'ڑ�	����c�����y��s���~6�쫝���i� �)v
?��u_D���4�QC�5�H]�*$R�R��H޸D����L��yW��U�a5�OK��*n��{��ϴ-=���k�5NJG�^`���:ܼ9*��2�䗝E3?��x5v� .qi���Zp4cn$��bO�ڼ�'�+���M�-����|]:�A .\ʜ'ܙs���D}8ޚwd.i]7-��6u����e��tFչ�"�䘸j:���:�E�L�H_�,��^O��(�b��Ϫ�>ܿB�q���1�k�ak����-
9�Lu	�j.�p�g��Z�qf�R����/�V~���VO	�����bx����i����j��p����T4�Q*wS��TN�S��-I��C0`�޷o�9~|F\R�{�fT�����Ѽ���ɲ�c��,��� �C��]=)W�����ꢵ#@��e�LN�=ro��i>���ݒ�S�5		Ռ���D0�o�:�7�ph����5.k&����>k7���R�~bjcO��BM���XO� ���
.���|����jB,7
F���T`E|�r�|�����j7�Q�Z��|�5>��P�*�q a�N  ��IDATQ(P8��Md�4�E`��9�������d-!Pn�b����Z#l;�/�H��|+ʟ�M���Â�|�<D� cmb.�#�(�hދq���|���0�Z)��Z�(F9/7˒p.�=+�Ϝ'�����*�  Fz	"� l����#�9��zW܊{ϧVVM��^g3�����G�*����=ϲ�6Twr�Y�;\M��ж�Sc�+��Nù����h�uf^K�J}�nr��i��>��	�6��a�V�Ņ`a�!�,P����8���0w�}ʜ8q̂�k���rC/��n#I��D�j�� g�)&��'&g2�J�l/<VN�_0u���3[�"���)���3� x�aA�B$��#�C,���
A�b��l��졛X�w��M�����Y˘�Ż�M� H�9_6E���y� �5˘�����'I�N��F䞁{g�uR (t�m%�g5�&�sIO�"SY�'��V3o����t�9n��=��-k_�p|�)-㣒?W	 ��P�&a�h�X`]%�Z� �����b�ޜ��9P�n*��޽�Z[X�0д�	���B���()�
H�W��i%�]�꿲E�����5)��[@�'���b
����O�ih�,\*M�d���>,-;���ZU���YS�f=���h��� ��y�y	�����±1Q�Q����� �tk"
ӑ�(�[�:90���tal���K���J4ӳ����X���7/֙;�Z���V{��<�!n���)!��l�ZR ��7o�Ι������p?
 G@��h��{z��y�,I��۞�\�]_Xt��%���]��Z4�?�~  !�DSW�����|64�kJf�o`�o�"��.���ZT
��{�;�de��f�K^s���Xp �qR¹�e����Фwaۈe-k�X����� u�v���h�|��~��41Q��)�U������!����s�<��t%������a}!��rm����bUuڹSbԝ�V`��� �Nǜ�%�=WA ���Xk�
� 1�-P�\,柺�Vk���&~!I='��U)�Q7���t�K���Ւ�6���t�.�L.�6�������Zծ۬&�񵀖�7;��$( ~�Rɽ������~���Ӆ�QM��淕~�P(�s-�rd��?�~+�y�oB8 H�M�'�@G��{���n��+x����K�sǰ9j�=0�mrr�,.,z.MM"^�*x�"d��b���P �[������X�ZO���K300$H_
�Y`jj"I�g�pB�����b���s���7�l��Ih�\�[��b�'�U@j������+�H'6(""�~�m��}v���&.�$��$its2���F T��V7�:[�7z���[����%�Q�Ɠ�׭�Ք1m��	��*_�UG����2����P|����;�#@Hg�Kr�(���Pd ��+ 	�R,�!�r�W�r���Z0�;愻C��Cwޙ��4\_y7(*(-|n$�ͼT�Fт�ɲ�-v�Y��Ǯ��H�ry�tǒ#DA����y,p��"�`�5���N�[�Q��۵����j_oK�E$�ՈF2Fwt�H����B"�c�8�VwoE���'Z���N��M�o��*���/]+˼�q���M��L�v������5|�,�~'�� 9�L�� �FTӢ �q38t�Y�1�}׈��z,��g�[�x��.I���fA�k-
8����O.�H�a!��?�L��� ���wX^t��c��fm���D������џ��j�����YO�������8�M�7[�;g
ܰߢ�Ó�eる�w�>ŦA����$`�_#���	�r�>���zƻ��wo��[�i���y����56��b���d��n~AH���p�f���R2u˸�K@pe$���|�ő����# ��\�H�HwO�?�T�?�������x���8Kм�<�Cw�4򟘀���Uw��{o�X����K/[õg�1��bəЫ���D�5�!���5�;W�[1�X�#Z�wUƦd��s�
93��\�cVF�G��r
ۖ��TѨ=^��"����K�Z�:����v�JC'e�Y��e\2^�B�H�������.���i���B�+�)�J�Lv�9 �����_�a����L9�,�`�LOψ �Ѹ��P��i .htHΑ䨀;�٥������s3��V}�!7%��Τ�	�����˾���U�	�f���%	7����5��T@����ф�^;y�u�y�{�6|����<�Y�������s����6dDjՒ�	K��\0�ujj��}�]��=�H�޹��E�l��k�/�R#�n��v��|S�^}V��q
lN�/�X����:X�Y�Xg�Cb�X ,������R�!tw#�aZ��8��渪!�qDlg����Ϻ?(g�.On������Z�}+Ι�$��/��8�4or�dZ��I��y;�$��6����0!s�|SǪ��I��&��g��܍<S;&����l��Ӏf�w�����)���>^&����oU1�O{f�,�C�����q��˵��p��T뀫'�����F�Y��&�W��֚4M�~#m��d|�S��;�#k��?��v.J8u��f;�-kn$�&�(�qf�{-(�e��VJ_{5�l�3D&U�S�h�QxR~ �ONN��gd�n��O\��Q�Dw�>�G� o�Io������'�$���] �I=qO��xL=6��LL�%nf�i�R�����4�N��R�6EVdX6䧅��{��ܬ�l�2���9��u�<D}nƁq�1,n�+��Ы���+����u,����>��v�[�~�r�LOk�;��e)�
p���߭�%��pT����V ��h�&�3���^sO�|%^�(�	�Z ���Ws�(X��8�,7Z4Q�<k�.K��Ǵ�e�vѣ5�#���蓲����%V!ж�
^L+�O�l�x���k=Gx�Z=]��Y�����ω8���"������\�T�.$��T�븫K	@�r�����9�}L�uD����;��>p�Keqy��]M �O�R��di��f�Y����[ڬ�VJ�v�V{]�-�J��32V}�i�P}d/Qk �+W�ف�IЇ&,d>T�"Xun9��}�e�����I�9�SՅ�5Ѷxğ��o+�{;�4���A~O+����WL�Rq��]���t����it�Fe�4��rx C=��N3k&j@��U�h����m#�>J�K[�����K (Q2���$
$]�i��C�4��=K���xL+���l-���e�*B4<6,��u=w�8I���}�����65��<tH�k����ؚCFI�XNIL��$k��W��(<??']'���39=9aΝ;k-h��
���E鲌wHh0V$0�����J]׸�= /�
^�z]\l{��àDP]�xAjP�wL��Ҽ�p����RhY�����Y��.�q]��eѴ�z9I7�=k���3j�s$as[ږW�V�������tA�ߺH�:��v�Wk�˒�J0�����aZ^AALч�j�P��'�N~��X)W$J���c>��Z�A�۲(JDf�uus�y�v+�����-�+\����"ﶉ�PAoNk=��
 ��ټ���B_Kx\�7��ݬ��謣m�KnP�O��C�]+��a�ƹ ���A�����~��d�j�Z����]�����l�*�bCfa��=�jղld�0��'X�FGo�w�}W>+r%	 �{G��'R���e����Y���iwO�����4L��.,��B����a�;����?��y��%7�P�fYl6����ޡ��E*@3��Z29��x㍦k�^	I��$�c	�nu@7!*L�e./V��%������a�Z�L�~��SZ�Z�$�.���Y���ڱ�9i�,8��!���U���[����M��8�9������J��49 �!L�	�Jb�Q�Z�ºA4%�R�j��V>W�y��r���X#��#�\2�!�T^�\nT�=C%%m��3M��/��=�o���-.juџB��	���џp��r����GO��au���?-���.��(�j@~�::LX�	P�PD%{8�g3#=�¹ �@��m,�w�$���؄D�u�c��3e�㾃C�����CVs�.H~Wp��	�ְp
�&`phH��g�H������]O������Z�B%<�T�[�����EFB��Y�ZY 9c��7�WXS �������O��^o����j��~Ҵ���.	�ز/`VL���E[��/k#iwޭT}M�/��̺n襏����=\����z�&�lJ�Y��GG�@���.�F� ��<$�bR4��Q4�3�q9�W�7��D^jW �yNB����՟Y}���$��-�
���<CK���;qO.��-Z��;ă�$�" �IR����s2�����Թi �\�4��,พ�	相j}uk�U*�L�rDP
� ��jb���V-ہ�~�K��$�� ��B�!V6�%`TemJ�<c�+J�������;;��	��K/JE�kׯ�\��vM��b�9������o^}�es��%9�豣�MId��9�QT�	��r.lހ�0)���'�O<a>,�7�^fh���}�I_E.ߒD{���C���@�0�Es�
&���͛V�6�&��\�t�_��fy;��*���^ý"��\�"U��&�E^�����ވ�.��U���-��Pץ賊jJt%��*�&���ȗN��|[��r���Vi�jx)p�ZL,:vuu�<5yBJ�xj�He�zP,���,�,<���Z�E���m��>)֏��z�L�l>����/���y�"�#mu_���O�2O>�����(��	��R��B-�����?�Sʕ`�PK����%���|�o�~�iq-����?����k9^^}�5�W�W�j���f�^�s��!�S��B�XXX�E�(�,�;)u��O��{��n�X}�$k��S��ڹ{�.(������tw9K/�s����?/yu�u{�A�j��/v���������/����tKֵq�~s�Yij��
��R�Z�C`�+l�T
=����䢴�D�X����U艹�"}L��!C�Chw��\ʱrlb;���]^J%D�%|��@z�ۖ��i�>42n����V�&ߣ�춺^2�;ha1���V$���v��J@�v�i��jknBse8�����������ś� � I��v�:��w\�93ku����-����M�=��p5 E��Q�Q��-��>�$e���af{s��_����L]8g��¦n��!�EpE�r`�`�l��[�|��t��q��o|]�s�N����
y㍷!W�VN@
��;��{W�^�zO����ԩ���+�F'.Z ���o���)��h=�Z͹��֬d&9֗��~�ԄY��2���v�}�� �Ii��Q�ieL_����H�	J�@��&�� O˥���dmh�V�����~�8@��j��r3��]c�h�h'_Z�gg�@�LAWڕ��B�?��p��u\�7�w�7P�����rs$oO0�4��j[j��NrϨơn-��kn/ٳ1��m�,5� @�����Z[+b�FZֻ��d�8f�?�'��u��R�#���J� 'c��۴z֭j���H[����^?��lbk�߭@�~���b�2\JY-y��Y��m�S����9"�
�rذ~�ۮ]#�-k7����$v�0���W�s��_��y景��G�J����Y��6��9	�&��C?by�Q35=%��?w�}O������?��c��[o��� ���ϙ�E2aq���2�}���[
�vqa��  ¸�K�<`N?)���w��Y�-X:���X� Z����l�̢a�[�h�dQ�R���6j@�SO=%u��l�����}s��*C�����9t�X������1�`�- ����]"�B/l�w	�an^�����K[��]d��)W�Mr��~+b�w�H,vie4<���K> #@q7�]���۹�+cG�՜��F��F�e�&�Y�5m5�):I�
jZ����3��W���S9�� �,�\��,�=6a��|wl hղ&W��f���uW;6�^0I���K�~O�K�3��-��~��9$ 	� �k�h�ͨm�ֶU�h9�}}���C&�W
И(�,|K-��o�5ö�믥�S�`�(ou~�d��� '��eY����߂K��/�~��+�(n6պ��]4a�<��C�Z`�Ǐ���j@�ZJ�e!|~�_5_������w&���G�gR7�%T�ς\LG�3o��ԃ����\��$׮^�m������qSr�����*r�;vtT�ET����$�]�0M�/�������{DN ʾ���>,������=,`�/��\�uW� T��Y�[)�5/ ?�������� ���y��/��u�D�|�7�����	��
���~�i~���g�}V*���}8�t�D�״�e'��I&��D��!��>���KX�boI�fo�9e���UΎ��E��8�L#�������.f��{�� 	��c�Í����t�Զ>�U7��*�&4��t�r��+}��
	7Q5_��3�.w�ȇ��u�I�mY��3�[Trm�p��8r}n��ϴ���2�D����*��B	�oe�Z���a���Z�ڙ1�g�[�J^����K/}�z>%��^���i�5Y�nx�zYc��d���H�����.�@ϮG���Yᤒ�V�o��%+��b�ݲ@ҳ덅j���8�l��3xN��﫞�Z�Y��FG�q�ɸ Bط
9���6��l�
�Cw�u��)��͛�2�b��� �|�d^r-\Z��{�g����Y@s؏�j��<��95�FFvKvajC�)�ie)�'�KA�o�Bꖼ$d�r骙�^0ݝ��Zr\!���|���E^s�L���k�������פ`%V(�ĭb��a}Y��. ���G��r>3;gJ⢫���9� hA^Gfn�Ӽ�ht@��=��w�#9|x���~!C�NWŭF��/}�K����0ǎ�~s�թ�-��~Ǖ���}����H"��u�p��DP��z��bY2uWH����ݼ�x���\!'!�2��b͂��L�I F.�wq<�����%��˾�H ���;(q�)�\�1��_��R��p��d�?H�8Ҳ8�r���-5ʕ�^I���D[+���uE�����%(������k�e�ES��U^W��4���g@hzf�t���
5��Kz�������/�W�\�G�zgݰC��j��Oj��0�g�.Xa�mҋi�n������vXlZ��r[ԃ�}
 ���M3 ��l�.��x �.9�壶Ic��'6.P��k������&�C��6]H�>љmb����
�D��� 2�}�S�����S��iS�1|�+�M��_��  4�L�@9[N��F�L����bب�3zs�[Hz�e�c���q�'G(ttY9�%������3��VE�ڣ�s^Y�T��u�قݰ;,����ݑ�Ěu�w�E5�ڲ��]|���zS$d������'��O��O�J����<5)A�}��O�?��?0'O����R4��_���8�ꫯ&�b%K��t��8p���*�4��(��ٹ�4���V�΢s	
Iγג�X��aAL��b�����{����?��? �L��J�br1 �p�u�^K�<�'&� rznnƜ={��޻��ł��j���۾��DaQSګV�,E�I�@k�BZ��:��(�	�k4�������DCb�"/+�_�:`#i^S�3&lww���9,Z��ܬ3o���mªo��M}��,�P���Qu�̲8����yZڢ����&v�����F^8J�6���I�j�.�Z�F�G��`��6�d�%1�&���/-'�%�ͭl�-��( �3zƉ5%J���:���klY@�壶�N�R�o,!�2�b�Ep�3��H�D��?y�������O˄hc��:BS��;o�-��mz���~O�J��o��o�ݻwY���][7ZI]-�b#y���K��z<�UZYw�Нj�L�T��}OY��"g�7~C�CDn��ƛ�?��E�V�����.]���GyD8�拗/�ٙY�8n��N8�z#t���A��yg��]w�e��=�7�NX[l-�G�D�py�����$y�RɅ9�����[އc 'B�����-�9n��k�&�$���Q��E
��{�XjbU-��T+^1�E�e�rnvo �"��%2���UB3r�&��nN��W	Y��e�ȒryY�&bb�BՂ�%�Y��k9Sfϒ&X}��B�\4�o�Ŏcdj����F,Y.}�Z������tri5M�� ���['l���04ɵ�ϵް��bgrA��B�� @;��2 �������Z��,E^��)d,�R�&a�7/��J>W'����Yh��Y�����?��f�t)��E��b�~�$�v\��U��AB���u�mu��v-�}ښ�8�,7DB��k�W9Fu��|�В����&kr�ĭ���&�h�ߋr��	��}cEH�i�(GX~��9��h^�����.D)xµ��5JT]�l�(:Nr$c����� (����ƗGhvE:�/��y�Q!�%�;�#1�}RƠ��Z?���ُ����� ��-4H˼.@��볟�lR����` X�
$�R+cϼqF�=�J� � �űK
��R�����=���7ϵY��98���^{M��?�����=��6G�M��������<���R��ҥ��T�k�ny,6X}�V�m��%�M>'���.�O\w���~y.R`�ۭ^�����^��,�/�Ż����b�+��:*�J�&�bI������Ғ ���Y���D�T*��A�%�ʒٷ����4==e�����b�̋�O	�ޕg���27��H��B��P�ցT�/�3i��L��Ǐ��4���Ȥp)����;����0�_���g��7�;�s���n��2��p	�	��Ň�GQ �������B���'Kˋ�tu�ryI�#x/u���w�Ur>�'O��>�U<܏EJ�!��|xf��zFLj���xct4Y�ӽ�ޖ�R���ZCJ���.p=�`G7�SQ���%���;g>�K]��'�>�'��O2���ԗjYX�E��G��C7SS��w�R�`�\I.ڰH��nT/�ʧ9o}���#�W�"��ՊX3���wF6�̹
Ijr��v�+/
 ��0ܚ �*�kpw|�[�J� ͊��C# �S�=f��8T�eȹ�Y�����:PD��w�Pr�x��XE�yXI����ͷ�2���3�#�u�
�8��'��rpRp*�3&n�W��Lu۸D�b�<ע�Īm.�}@�V+bpظ�U��o���>���+��ZC�qwa�����\�xI����|H�Ed�ۙ3g亪��^u��Is��{�X�9�;��H^/��i2<�f����|'��ӛ���V�هz�:�jW����̤)-/�=gV�;�
����o�@R�频ݻ���g�\�n��Ϛ��^0e����3a��i��jmYfXOo�X��Ek��h[��J:ٻ���02?RN�>-��Da�v�ԙ��ȡ8��c�wI���8�-�yl̛���.]0�<�y��d���;zv������M�XB%q��$� 栽��Ԕ�,B�Ü:=7%N�$B,�k�Ӯ�tN9a���o�?��?q�̎BӱAy�|����N����gFo�p��Z�f�K�m(���W|(��G��֮е�DO)��Zￕ�Yx�-�	�����Y�E�q�J'$��e��4ܴ�����w�d��~`����{�PH>]U��{	�Q��m�iZ�~^v�tJf��,v-��Y�/U��y��l@�f�[Yk�����H=c��b�E�h�ܐ\)���p�!�	�4qn�8!K�sgͮ%���g~e��;�ݟ�y�=��(������Fǳ�ٳO^�2<'�2%������S��0C��d3�7������9+�v
����A���I9��gj�g,x�y�Q-.&�I���!���%�o�֤���� m����������r<5�ʎ2��q.��D	Ӿ  bu��?�C�O=f�s��iW��o����Sr���F.+I�gǡD{�lz,P��-efl���FR��RZ4W._�@t���]5�
ނ^~ _#fd�^��X���ől�X�v��{G��+��jS�#�f(�T��d�����<0.@@-�+W�ֵ-5:y�R��������f��=����5d��?�}�yYL,J��9��F��{��Iי9���恇�������^1��a�&ك�#�ϙ8�b�u!J81T�������N�k�CX�?�D��I3)>�Ϙ?��?��[m�2N]kT���������
���jK�9~#-��R�M��� ��uϧ!�<�JCZU#�"Y�a�zݭ<�(��sm��r�h���w���q�Wd`��X���6QgN$VL�?wY.;7f'n=���J�Lk--<*l������ئ�p3n���%��`��AU�%R놈��6�{`���9��C��[���._�$�/<�is��E���l�E����R#�/��A� ����� ��as�±��[�F�=6(����U����M�!�i*�zS`�Z?�$S/4n"�!�iy�(�#���;b��B�c��y)P븒%���4q?>gc�A���m����I���<���`�D֓q@�!��An+\U�G��2<䄱Ǫ5?�ʊ^yD�@���~:D^E	x�7B��@
���:��Z4-�H�� H@�O����}>��r ,P�"l��j�<�u����X\P�?{��y+K����u33;f�U;^��ٌ��ٽg��Es��9��dqnٔ�˦oz��?p�ԫ.���1��NQ�0ؔ<߈��3�3���+���G(�����V�-5ʝ����BUTGs��Z��� f���Q��a!A�RWt������+�ۨ��P��v����K6�("�����t	�	Ȃ��%n�dr9�m���T�	c+��u�F]�.�f)���~�$�9�`ba�6�t��UɁ@�9�I�?b��߼ς�;�?�����쏞��j�s�d���i�㴑cӂ��V�~3�_�����+��)�vɖ�->aJo�<�,�޳0Y��W�~+�sjJy�F�D��o���u������tYA��P����h����ǟ<v��9v�
W�[�VӭV��4w�s���	+-��0���,WH�\�3��9<Ǭ�%�I=o�9Km	�7l�;�_�y��3�i�!m�#��k�]��VNtط�90h�>u�y��wŪ;=3).�ŹE��#��G����3�ܥ�&��'��YD���p�<���"B�=�����"G�0���k��?�/�w��kW��QR����Pr��%!�֤����_]Q\����Ki1�X���LtS���}T���F������O*.ށ碏_~�e�����$���w��'� 4kA�Z�t�)g�q&��7 ��J��@��G��l���K���;(����'k�q���[uٓ�^��4�r��_�\K埀ͲN�2F���}�x8�&���f?P˞*y4��c�e"�����9t�����l��R�k~a���O�s+�V)��E��9������)k #��x�.ɡ�@�Q�ʒMy��eG��F>���-mK@MZ i��B��k����j&׮]�A�p:���_���cY�L,�/�$F����v�Λ���77F�xԜ7�33���ۢ���V����KUId����C�Z��#��8f������;�s����?D�a��^hB�*x��eCb��?U�)�H�>�7�؞���jk��җ�d�߸n>��C�W�,�1=�Ն�n�_0h�V�B����T@� ��8��Th���,�Y������תm��)�ڢ�ժ��� O�"+9�V3�YPs��;̑Ç��g?��ДXSps���#��;�_��/%
!'�՚�gB|Ը��ҭ�J `�;��hk�I%���m�I�����lҺ>��#���~�ﴊMl�y�]s��e޳�fjz��6���fd�u�·�����}�VG~߱c���#��X������.�Q��+|N�0�a�ƨ �����c��k~E�l���Sj�7�P-!�6A3%TyiA�f�TB�q`9�p��LB�;�F����G������ ��q����~��l\=77<��h�� �1F�G�MA�ȭ���_�%4=���ZQ�<�0���S*�� 5r�`� �/  ��Ν#�(�I��r����.�N�c������f~��I��2U�� -�A.6B ��w��~���otP�:��v����m�i��g�+/�B8�1�;�fyiє $�����vN8���==,��kE�W�^(N�����C��Ȼ�<4�P��5��Q��ܚm	 �E��P�f�3!)���탉��!#�M슜�d�H)@?X?4�5�>�&&�W_��]��d��@.Y�{�
{Rn����:�2d�]��	�`�r���n'XL�$�����g�?h�<�xᢘ�t�}�L@����~��9�I%�A2Ӧ���@`r0{>��3b������P���7K�o&f�r��?4�v�ёD7�6��t"����}�&w1a}�0�a�zJ�G�wneMY�+i#Mݞ�7��;Ⴄ@���\���w�k�Z�,�/Z!�`�z����2���l���?>+�����S�n��o�ϡю'�����ílk�"�ǩ���,�´��C2.(.\���%��nWGo�љiu����n53��d����~z:�����C�c��S:��)tM�����Gb��D�Eeh��0��u�#�� � �_���}W�ܖ����$��j���B��$̸f7F"od�.EW��SM65�!��ܑ�ݳ�&��(t���P��;�p+9�W_סXbP@s�
�u�b������Pe-E9��1����@B���>ĽQ�!��3��kR����uB��B1�����]�w	?ڄ��se���+���5%<>j�D��gL:Q�^���d�T�@ͧHI܋�����9ϿX\�}nvj���~�p��l��J
ɽR�G2���*E�Ū��FB���}�]V�Z*���/��+5��$:Ym�{�Z�"���m	��rC��ݘhXh0M2H�$p� !�7������$L�V� ����^�`�$��M�"�q��v�-����|�#��GX���L���u�֡��a��LW�31Oz[���պu���~��^{�z%��
-����y~���0�I[�6@�F��<ɩ�I*���f��B��y5Z��9<�]/�9�Ƈ�J���ݬ>,�(����s]��K�mI�t�$���C�9�9|���[m���5w�k�����t�r70�S�(R�����pi�čt��y����KX��3hńv2ov�1=�}f|r�\�
�����[�7;,^�Dh5��Ah�k�V�K[2�
��hE�i�~�5Fx5r@����-Ǩ���e�g}�!S4qfnт��lXq������JJ�ݰ�Ee/ᖉ��4wC�Z������ \ 	�R-�*C(�qx6\(vjU�W�����V�@H�&�sn�0�_�711n���M�(	ݜR������+	��.��;��]o���Q"�(���C�壏?w;8�m��c��(�����	�Կ�y��G�{($�r<��YZ
�vӲKǇ~XP7�l�I8��VI8z��-EbU�k%`����/|��w�w��9k��.`L�_�.�J��B�{z��[f4,���8�y��������j�&���v��Y�Q^��3�|[���WMO�����%}�x)"��R����&����|�ʞ��F���{w�9�Ywg�Y��jK��_bn��3Ʈ�Dqކ�-���R/ͅ���Q;���g�r�MR���E��S�����ʻl��k1���
Zt)�k��3o�7�|G�^=]�r_�#3?���e�T�v30.|f��nS�Pu�.�N0:5ݹ��,&ͤ����s�H��$�b�jaJ�k$�r%Ĭj'\���۳��h5׉�[�!d��{�FZ% TV%�mUP�ᦙ0ݘ�I�8v��.c�+n&n�v�6�\�`\�pP�;��ұGH/-�j�\���Ñ�*q��Ws�e}�ހ6�J�d�ϝ;�\ ��?z��Kl^}�U��j����68�vݔ,ʛ��.S�W3��f�n<���8w����%R�ޏ}�s�����q��,wV�wk%��n��|?�����6�eqs�����ԓO��>x�||�����w�6Ǐ6@*�>�P�9�T1Kܪ>�v��9����b�Fv������\���+�((JIi��_��
��#���d}�fjU��5�����r��r36v����ȼܿ��%y�J���o^=�W�ފW��(��:����XnD���NV`����o"H4�:��C�g�"����>����������Ԅ� �?����,�&�7r�0@�QM�m�.�E(_̍_�����?o�䬀���O��~�i���jËbq=c�޳Xt.Nn;�0�<s����9r�**	q�!t�='��Kj��d#a��[��d3�}-�a�"��,�~�.2��vdrcN,�ł��{r�%���q_^�7��7�'������P�Ǉ��Q���U�=�ݭ�Ԅ>A�� ���ʤ�3��ᦦ�V7����nġ9�E�0r_A6��N��P���s���{�>}�Te}��'̀A��^��0��}�z>"��^���C]I���fe-�Y?s&ê79�UR�'�/LP|wo����>[f�%Z�X�bٛ�]�	���A�H���c����r�-��`�R31�!QƘFm��|�s:^#ؠy?4M��g(��q=��0�cRGx!�4�����@X� ���m�>��Ss&^��O4��v�;����؄�-u=��g�Z�6��cb��w�}���﷛A���� 9|�3o��������3"��ln��-��Zpu�bgn37��̭�7��	�r%��8>���7���{lԨ���$� .�&��nZ�5k���|��3��6�Ξ�c�?f�ؼ��[�ʕ��d��/�4k���	�,�������]�C�5BP�ʫ����.
�U�n�axxPrlE�-���&M.��ٳ[ ���G��k�n�sj�`�ў��3"��U E#����|x��۹)*�U�"�|i	��$��g}uJpR\��9�z+WhxxH��Y����T&(�A�#:w�d%��:y�W买��~B.ѰV��:;o������%O�&u%�D�o.�߻�g����ɼ��Oq)M�`ƅ����E�!���%�7�2��rX����|�����N<�9Ƶ�e�ƪ��|���e�-Q��g/.�]R#�w4�/����ʼ���8;v��{����f�2��G�w��[���R���BTMH�f[ڶ��T��E-�Y�Y
�;��bC	u͙|�g���	>
�9�N��v�J>�Q���"�2�z�a�П6�V+�I��X&��\#�v���i3a7�����YDM�l�<�T�ͻ������YSA\ȁI6XWu�qE� �Ơ�c�d�u��r9	�^������p�@�>��w�r��Z��)9
Β�Ӻ#����f:$r��W@��[444V�*��={w�Gy�<��cņ��y�}�Q�[�,й�=єy~���=�x%��~��ߗM-�Mh~Ns��/�>���<� ��p�H��	�J�e@MN���3$�*lt��������������fbr�,��͹�g��̬t���-���%J0r��[m��;�5���y~�Ɯ��YO���Z+���W,ۆsװ�/�h}�Q2�̡Çe�b�x�j������z�p��^B��̄CCf[��o���Nɦ��ܼp�t�S�r��xZ]�)�]����/qin �X��åa- ࿐���U�P���]
jP��gA�q*��Ve�]󲤐��F����{�kI2�
GΞ���'2/�������J\R܍IJ�HΚ��$�"tE�[hU������_��T7���%gc������G�㐕IE+��Lʏ,��y啗%�`WW���Jx>���G��ݹd�s�9~�;�7�^|�|�̎T,�����X�jk��{W }���#�+��8,n%;��D�s�g5��V��o����ފ���ID�K����:|��1�l�F[�3�#��4�'��i�	�ʘ�E
�a��^7!��ϥť������� �;�LP7�� �hA��2Ij�[��B���e#�0uł�e1E���>>�DXUk��wg����(���1���!�w��|섄�u��Ӳa�$��="��e%���`�{�q�Z���:�#�8f/�������啩�>���M���wq�ۗ�Jfڂj�޼n.^:���#3;7o��^��/����A ?~�j�{$ʋ�A�5}��w����/�d��K�I�\Cj%�y��H�.�זtLB�V"t�F�f���[��4oh�T������7%����yb=����tS���wfzjڽ��W�]3�$$<�>��Ĥhi�D�~����f��B�~����w}&�mWӢ�ƯU-[��i�Ig�||����f��Z�˼����`���$	��\{��k�y
@�T��X)|�9�4 �Ͽ��o�yt�*\�*3*��e��	(��`H��+�ۄr�^|�g��s�A�[�,J��d�5��X����S��kiqGu#��Ѭ�*��p�([�O-C;��xw� $@ۿ�ĻH(��Q�Raq��O��ʐ0�^�I�K�y����O�$V+�
��w#b����%���{)W ��.^�r��jB����P�� �����S@���h�]RE�s�Yp���Kb�j�R�c�D9�j�����E�W���|�W��e��Yy�{1�c��ppF���6r�
��Ȧ��N���!֚| oGR�m��ȂH����B�"04�[� ��O�����>'SK@��x�l�s&4�F� �#���A��₶o5��/��ɂ�w��I���K�����+h\�H\P�rE������d�����`@+2!�F`!`y�0#�F�7����/�"h��c+9X�D�	�t��13+�~��:�Dì�Y�Ր�M	i��!�����L������ȅNH%
 -ד+�V�ʺ���FwO���5SV⫇JCUW�KB*ۿo�9r���-n�iY����wR��3����4����(�N{qUt�o��u5�����4�<6��֫�Lb�9*��:��|)W��6��F Bh�+[��=��E�'["�4=��νl�I��� h�݇[���W��*h�7^�l��������V�Z,X�cB0e|�m=��Ľ�O��1KV��e�&�����bb4��9��������K�k���^�5���Dl! �Ͽ�������(��`��9�i�q�/X.���=2��.��Hd,(�,��EH� �>�����z'��m��B�>���4u!��Dӧ�b��~t '����$.w�2���M|�*�D9��r4(ؐ�uu�_J��m>G҈�1�#�$:�^�r3��(X���Dv�
��h��w�<��D%W1g/�7����U�Y(��b�Vp��?ܛ�����K`�rP-˾F��A؏~�HbG�c��--2�O%2["�jV�zK���;��3��0�E��׈r<�w:"����f�A0��(�&M����QJH�?���������S귉X��F;[�1p$��O.�ؠ&�)��,r ��dQ��Q&K��];e�h(��v�I�0��#װp2��Y8d�<}�^�D$�#�dd�N��3mB��b)�^q$<�տ!������\ v��P/�>B� .aN�_o
Y�"u�~��XΞ�8r+�W��ZH�4,[ ?��6[͜J��{�g��o�����w�۹S̨\<��XlZ%�C����$'ɫxw�>9M�����<2��7����>{E��]᲋�w�U��KJZ�ą��y��ih�� JJTVOvd�RBc���8`�j���Xq��w �U�n��a
�c2��2Ԫ�)��"8����aǇ�s��W_��5,��K�)Y���x�+���ߥe�w+���+�-�	�$���c���9U��>�l��H� 6��f���|-��ً?�
�ň�魯X.7��z7Fo�B�߇	�y����!�����A	�em~���Q$���~�3V^ޟX@�f�=g�BY٤k�{j�.�ڢ]�s$�,v6YO����e����[E�ޕc��,W�I�+Ƃ���)�$c;�ໝ�#���UT��L����k���~S��~BƒM_����:�	詉��H�N��]���9�¿o���K"� :nh�I%+� ��/&��ܗ[�~w�ś��}5?��\>���1��Ef���"�k�"K �Xo闅��2�P~��ڈ�(v�K*o!�?������C�sfq96g?����-�}W�˥� c!_7=ݻ�<:(���,��6�-5i�_B���N�J��qG^3R6;�)6T����i�}��%%���${�rv4S#ד�va�=���Ӝ�d�}ffjVj�C�:���/frl�,�/�A��`�S
�U-p�s��������2��_d9'a�� ��* �9!�}��ߕ�W]4�4`ɲh_��j�֬���ШyB3%���=�yId��J���M�hN.\��Uן��]V�U�3��<��	 �Gb��<���X��{0���7�g��F8�ը�����w���ܗ�F���?�33`�52�B�!s�� w�GO�ǽO�dQ���>k�տ���0�Հ7b���%|؂�N�p��+R����ե����+�6՜�||!/�����R�����y3����J��Ӏ�]K��v��\+��[��t��'�Dk?�˾\���e\=2�Y�d�.��5YV%4[�ʾ�_���ú߽��9���ۦ�ʹ�� \���)�=6�;>Ga@q`�T�ӝw
��b��g���� ǆp@!c���@b������@Q�bu ԰�X���ͱ����~�{68N�:a��J8Ys�329��e�r,��Q����e��}���c���#�:]�,�9�8D�b���U@�Vs~����;�#�r�����������2�K�K��`�ǫ�9N�����aM(�d��T��* OϿꪢ�� W�8�-}�pTZ`�D�Ă�=qU��� 
�Z��R�fJ�~$�Hd-<����Z���Vq߹s���/���ys�����s]�,�J	�Pp������~�F�i[�$�)�5�&�S��20j��-�����y�11���.��8ݽ]�������'�Y�^�@���)S�&L4B��>,�6��n�.?FN4����}���v"H	���Q/.��c�aq��g?�we� ���K��U�3�I�>d[�� %����3��?�z),��i5����Y��!��{�
2���~b\n�5|镲�����s�0N���������=Z�3�;�IΌg��D4�3�)��!QK�E3?� cA?B��y�fp� �Ĥ���
��ĚU�.l�X zh�~jۃ<(!�� 2sm��) ��K'����i�?Y_���"���0����4��*���N@�r����k�V�͚Pn�@�ʭ�, ��jsw��Zx>���s
1B��oA��������7EhDn�h��(����Փ����^���*@����';�bP31>a�XM����w�#V���O����� ?q��͹"�_�ʗa��:W�(�bqb�cef�F�~I�G4kT-����J� /���N�A26PI���@�X�r�Ň��j[��h9��J!�hEo��x.�Wy�J�2.џ�����y���B��Q� �]��9�|��ե
d,k���,�4L����;�$��'�P+i�9�rph�󜜂ȃ!����͊�ː��O!
�L��W\��R��sD�\�`�/�e�{Y
�ο�<#�So�s����1dܔ�������ܶ�E�L8%5��jc�@a�U�/a':ڋv�.�ȇ��+U�,r�"��Τ�$��IG�f]E���
�,"�����q��07Ʈ�مq��x����jioW�L�b��O'�Y�o��pC����+�����}�"h���o)�A|�� ��ёL/)3sZ�ik�yh�V\z,
����s�k�]xD6-�贞�^Y<�[o�-����͟,��:�}�sͥ�R��J�I�1Ɠ w�34�����/:xJ����AG�^���6[�lk�j�Tse�y�����:w筛Y�P��G���;���>{�񻾋0lanP��<�1�|��P�9K�a"J ���v����.��6':t �έG�9+��9y� ��[�M.�
!�����6
��=�a�RM����7�[�6���ǏW8Oo�c)�j��S:��~�l��K)��M�������a��<b+�G%�������Gh�A4iܽ�����?o�\�#E��ۍ�-~n�	o�I����O"���)�9^7�k8�I=� 3K�fs�U:�룿�QO�!�u��7�;���=��^MXS�Զ����ŅŔ^Nߩ���"���T���P��L+�Ew:�.:��PV��G~���D�����ǏӾBf�G�"�'��������"�[�a�T5;E*�C�c�#��O۸��H	%oD��=�ߑ�KQ�{�H�kC&_�J����Srΐ+8B|����z�t"\��c�\nJ/t�N�
���ʙ3g�}='c�����swx��8�EG���SD��H�tk��
��M�i�!D�4���37;>����y�8�K�Y]�tE}猊����1�w��2<��l�A��K7V�o ��T�>H�P�6����hN�ԅhP�&g'*˜�yI�$6⢖,��zUW��+���}��s
�B҇�޸xV�y]�O��=35-�������p�dO^u�rq���`4��($7�������S���	�k�0	c�ʣhl�k2.��B��l E�Kj�j+�L��k��a�R2z���hK1Tv:(uE͚��?x%ꩧ�e�g�+9SYV!�R�R���
��!0qW���o!^g���a����wh�>���J�� ����������>�g�m�ya3%
�w�D]�F%�+���>*ARA�4c�I�*�l������3��<�)Ej�2J��PI�t� t6��!S4`sRx��nQ��m����Q&����5j����vPñ���Ώ"�Mk���8�Z��/������2N/i����qm����z���(2�9�1��*~_�Tǰ���ߨRm���(�m�K%�L�^�|�%0~*�l�{
�{GQQce�C&pƃ�{��$�8��؇��q�K{��SEE`����:x蠘{q�0|�;�������� ���\Y�Fך���`����1�) k�^��6QY�V1�x�^1���^���!������g��|HNՑ#w�����%�D򉢬��W��kW���q°�Z����X捔 cá�\33sB�}�����'����A���$�����ѣ�QG��[�~��N�%P�td�#3���u\YfP9��)���d��� ��X�yƤ���"X��W�
�2��yܖH���"���lN��&1���9ҡ����&rB�n�������~X�������|`�J{ɐ`�r~�B|���U���;�"�xH���V���� yꋛ�]�4�W���*9K�cNr%��)�>$n��Ρ�F:�*���д�1Fg��GO���a<<���������pN�N�Z����Q���T-g{���բ�AXeN�/�=�R9ߢ-����F��|���3�	�lrl��*=O�`�3�g0���&�
>
B��Im�SG��^���� 3v�!q߸t�?&�ߕ7�n��Q����4��%(����ѫ�u���eU+�Jg�
mP#e~�(�[��Img����?b��o���ΑRF�"�L�Bf���w,��(�0Z���m���H�����@��"\��{t��T�_7(�-�'�f)��f��y,������(O�k�h"�w�u�ܑ9�#ak�_�=��Z����^|)\�z%�E9�~���W�"��ܘ޴�j���=:�i?�����$'7�/��j'�nXX\_�ۯ����GDqX�39h�y�B8e��D��g��0d$p�|\N(��}���e,��<����;UT��ۃ�"�@���ݛ2�����gO$Z����h �tI�Y�X4��g],Fg�VPZ���
ب��4@늎��Ǖ���5�hr0m�yժ�x^k�0r"6�1�>M��� ܯ��PY(���3���s�0�}���"I[vg�|���'�����*�%j�������4�_��Z�K������e�r�ٟ�Y-*�6`d|�P��B�wJ�?���Q���*�U��l3�8⾭ª���s�<{*�MI����;��ڑ�&5'��ٙS��t��2��`�f�9���΃��g�}Fcx��G����>��~��.#��1��w�1<����L�j�嘚2&��(H�l�Y��.b�C�&A����k�K�)b���B�=���j=�ó!�Ee���!D���#8.��1���*C9R-u���S���eT8��}��J��Ԧ�4���)頷:�q�ҫ�<��ę9��{˾^]P�w� ��ݨ5�qd��%�f$ґn���Γ���T�p����6e2f��@z3�'���
��=�e���2��ICܱ }��N]¦�OVV���С2��*P��da�",+�Ǽ���6���X�4�"��8�MP�8ҫ��@k uZD=Pߜ�����{J�2PRy4�"�T��p���F4��Av��8.�Hm{��m����k)s���%2��Y��0�<*��0l8/�A�b(��OV[�!��}�ݯ4�!�1�U��L�&��я֤8ܦ���"Di<�S�d�"�N�p�|X]^�k���4(�ߞ��n��Q-�
�f� Hj�m���V��8|�Ĩ�ܫ��oH�8w�{�X��ZLLIX��E#�C�>|0�>��3.P� mU!�ٹٰ�`dZ�S}��Yj�� �'>��*^Ξ#�U�3F\D�<@��U�ʂ�`񲸉0 8�,�EH9"s�"�^�_J�ɿRb�
�Ͻ-�#����� $6�3r�J�c;�9�3��/6��}卣����3c "����KtY�F��+1;3��D�EE�l��{_4�+�<������m�s�^Wć�%��������޵s��/�	�EC��1�k�t����L��!|�����{�i�`���Q�����*��j�[rP�e�~�H�?8����/RT ���-Z��Ҡ&��"�"%C��N�v���V���+��w4&���Ʊ��9����%e@J��ao �dzx�#�7���9%5v�o#�T���m�%�f��^+�ƽ����>�|�"3lL��1��-^�Fg=�oQلZ]���ƍ�m�)���GD��V�ן�(j)Z_S���crj�򊴖k�0gͫ츴>r�h�#��ަq�<^6�����b�����{�W���q9:cn��'=���<<p@�JWz�)�8��鶊 �6$Ԙ�~��@c�F�:�v�c������H=�P�W�b(jޡ��Z�����9�[o�o{��5'/�/�����0zu�+Ff'��,�R���As�|�����֦,8�J�A�\܆㶤�r��+C���������k߻*�7D�P��"����ע�m7SY_=*����6��;�b]�Z������915B7Γy�o�O<��0{}G�6B�֔g�󩥔��N:f��RB�����A�+��+��r?l��D,D���G�G�H���B�w�r�0\����?j�����Gu�o�	�f6�ư��Z/� 
�)���s|	�MJ}�W�x��k�z�AAD��°�Tݫ!$�z��%�jy>�m�CX�f;�,���hhq-��7lc��h\dؑ�TK$jq��N(�v�'��cl#B��4e��2���7��m�'����Y)������3/H\[��J��:�C�
%�6l��o>V��,�����ˋa2��p��Գ���|��a���z��������˕Ѩ�'���ߢ�V2Dy�fܹ7�5�H���L~��ٍF����n�/ބ��~�00�pQ���0��o���k���M��C�n�^/S]�z��0~Ir�4�V�uS�L\_.���<̓�������d�DI~��~�c���?/��DLR������<O��	.2º��z���;t���wiG�#��A,�	�D����õ��Х�|1�<�H�_u9|T[-.���d����x���h��@խZ6}�u�����W4���5+B��f��m��) �TfA�;XI}��BjnP8�U��t�,�:�4��L=2x�<D�{F������pyF| H���ii5�ğVcJ�Ŵ;@�
�Q�Br�#,?�A~��Ǫ�V��_�Zx�ǔ�d<ޣJ�~u����3i�z��b��!��1�q���y?�I��P9X"3����*p*��йw�����o��+/�� l(����N����{�0��Ӊ���"b�*f�ο��d�	�~�ۭ�!�G�;���T����'�U�'�c�y)�ᛖ���Q�p��h"A�z�1%lM�3E�\�IP�!1�������{E�S�S"�-�FQd/��F���{T׈[)?ގ���B9l���j\p�p���˸�{W��H�R�wҗ*?����گ�H��_��]U2ϔ�p� d_��$���?��z���h������0��Hs�N��ix�3��w���t˸1������g�d��1�G�@�9���ܐC���c��|s���{�1�7W~�7�q�?��:���������IV�r�FQe"6/Ɂd�%�S�khY�Y���'�_���rR��;dd�w��y��%�X�"ڣ��T9N|#� ��(i�n�ݸ|��"� ����+��"Q����-a&r�VSLR��S�Y�,$3A�JE��kS������Ȋ��w�U�%��6�3:nC�Ʉ���\;�����];��Xl� ��F��3;6%�w5Z� �5���PX�6�ka����]�����A<��o6����	�7u�) ���v�H�0듨@�-�xSq�D�ѢŒ���g�g±��u>�A��w~�w�Y��$zC� ���-�y!�����R<������_�e���~��*�\0l�E�/��� (s~��q���}��l����޽K��}�Rz�?���F��	���0X�xD�Pz����©3�����Ǣ�f�g��aB8��yuu��4٨B����="�����o�7��8�	��0�$nfcw5�"�������J�!���V`0ƼO�M���Q�S�n�����Q8�Z"��_a������u��\P������0&��P(��'2Hy<��T��Q�� ������<�{�v�����E�+5�t��׻����s�S��cƑ���?�Z��{���19�_�,�:C<�3�=�4����2�T���$��n�+���מ��Ң�7�	3NVU�I�?��?(z�8�������(����YQ>��"��QD��k�6}�K_�a15�V��̊���gϮ8��*G׋Fh�,�V���)z�"����޽�?NU�/����W*�j6�g��Np������-^~�K��9��OQ��\`D=���x7j���_	/����5S���k�jX���b��y���~w�[�sEe^0�!����M'&�`尜��!PBrVNY(\g���c6 *t�ƒe������*�ǩ�R�YU���+�AT�9��>��x�(l�s�h���#�J�3\����O����1/��=��(t�IC�CB��{�=��0>"4 �Pn�ӳ��h�5�� ���(k�M��2LDa �X��H�M�,�N��sN�1��*"��ҩ��j�C��(Tʸym�X��t�rQ6+�c�����B����Z�e�%J8'�r&R�Bŏ�ɐ���`T�|/�B��HD����;(ү���;�;��5�;�+1���Ƞc��f 9��=5���q��n�3zl����_���L�y��/�n��ѱ�e�Q�_k4�4�Z���׮"ԩtٍ�ɓO~RCd��"��acm
�%x���p��=9|�Nɘ|���}�E��Z�� O���h�ƽ�o9C�ם���N&�ͼz!^�q�^O⊱F�׮^���)9���
T|V���ːv*3���gcMQ1�0�9���3��9�~�J����S�t`��}H��Pf =��6�Ĩ%�a�Q����UFC�Z�������ˑ	��=�z8}愰�9�����Q�?���jV��t����7PnC�!�t��4@�i�g9]y�=�3��fH�`|8E� N>�p=4�.��4N#���(�t�&saN0܈t`�q��d V����v�sn�Ȧ��r��f않��⩥�2��a��%8���z��ޯ��pP�v3lN�'<"$0��z�FLF�3@+��ޭRKM���5ό�y�:F���u��Δ:ór��Q J��t���r�Ѡ��׾�2N</<!���s5���[��G_�'F�g�ldW�T稀/����r�ƣ�<Obn��L��;�J[p��Wʹ�7F�s0:�u�������蹓�=������NpU���U٦��6��b��r���~��8#%��vY��qx��Ɣ���z�r�:�d2���ѣ�§>�)�a�=�U"�~=d! y�aD�iჃ�9ܨ� ���U{Q2�?�h8r�p�%�,#*�%��H4���>k��Y�!��6�r�bP$��ğ� Ȗ$�A�͝�[��kz�����TƑ���cK�um���گp�>9p�V1[��6�������+P��*�'���t@b�GD�P"|)Z�k���j�	�̈́�����q���A?�U�4�ԊWY9n�?(��o)�`e�j�V:�^Pݽ�s��\Z��!��&�b�=^��M+�L�����ca^`,8ʂP#6��S�.[n�ќ������-�{U���̵���'����p����G ܦ坯��WiJ��x��BH�=6�w)G�ad�8qRx([֗��!��qN8 cаdzqL��9s�������骮۵0(����zy���ٟI��]�4Ȧ'�?Qn�������;�������e A5�Y�Ѻ�"[a+�SZ[����I`(;ӲG	�{T��A0L�ӟ���ϳϟߓ_矺A�v�Dzm�z[�y�'.ow�o���=Ǩ�2���%_G[}o���$�#�ҝNʭ���}�=Z���!;���;��1��������$�b�7���L�����F���g������k>�!%G\��VW�Ɇ�f�jF}�
�֔U����U�|�׭�K�cFH)��
a��D�WD�рvC�JU��VE�Q��4���(k�s^��m���]�m�~�p> W��<2��c�ieQ�>e�n�x��{U'�z& ��ɵ�KX�d��n�仩.��jAr��}+��V)8��5�v�����0T�`�h�M膲�
Q��J�x>��ݣ7n}�ƗVoDt��S^��
ۻyXxt�{�>�i����`p-�a-�����q0D;睊�{x!1P�CZŸI;q��1p0�0�^j�z����:�D{J�&�u���7�����¸�k-l���Ф�⭽�h3�t�(օn�����#_\��8`W6:8&���a�CO"�[����fF�8�?'?�ҠN�5j��\h�{Ν�|�oś�j̣�	���)������6g�@�^���hDX��Ȟ�\�^�������x�c�A�˶:F��Q���^;�(˶��K��s*��ǝ���i@�n�w���Iny��Gs�y�$�>T�y�6w�����;��y�J�
7�F���!B��Ko-���V��8%�{���`7Ed��K�	&aN�"��5�>%��h�Oq>kr�\����� ӳ߁���V0|�9��lG�;�i��sь�8N�9$��U@A�W6���7%]U��aj|Ay
ÅV�Y��0l�xȣ����JIibY��uބ���0=ۗ�tD�W\�G����Wػ!6�:X�s��rO�5i��zO)��d�S���)+���9�T[e�$�nW~��<���R�0En�y�;��X+e�:|���~/l�-��,�n�Avo���U�9I�J����ʄ)�="p7�S�Ɗ��� ��mr�",��80B9'�f9v�̒*��h���>����&�3'�.̉����UW�kr��05�1�!�a]|������ ��؂�Z��̌"Y�����~�R��k�y��g�}+�8�s�َ��7��PǷ@gJȗ�4+��1<�Q�v�b/��8��L�����P3��bv���b�S��|\��[q�Y]>���N,]���v���ILP8I�W�=�n*ְW�}�X�؀T��HF� m�ꫯ臦�jO �,�$}�?t�g�w+�td�l�;J�xvSrן�Ǽ7U!BY2�$��u���j%$�\�w��s��������Ͻkמp�Σq\���3auiEXdG��v����p���p���p���µ��q��|�jjj̹B�d��MU�o;X��5yߍ���%_|��&��O�Q6(�A�p</��3�۽���kׅ����A˫+aq���Ơ���ë�~U_Y���������� �ח�m������G7�������qa������9W(|8\<,6�IY�;㣥}gf�xIoU�����r�*�����0�c�L=�P�܃En,�憩+2�J�P��T�&�y�7�N6ɠg�-t�(S����O�&,<JY}=��P+�gϜ������X���!E��u��)#���!�� �,�	�ZTa!��GzA!4;�c�J�׽�0߇_%���������[�����������}0"�q�n�K˟�����h@e�M����$ʂ�Uc����aN�IUi�l�{������v����FD�)y
(O޲��<����!?�����*�t���(=���AY�h�SP@,J
�&��Y�Q�& �����=��2�]T�
[SE��jHl8*� �$=��4�d<Tmf���z���g���7&�N���Z]8 @��u�����vw�59���U)�a�Cw�*��ξ|��Ka~i1�ꨯmE�)y��������C�������a~��zəF�������bw|�m=n9P؍� �.0�:
�o�EL:���������|,]GokѴ��Z�'�@In"J���� �z �¿�v�ڕ�oϾ���gC�����p���(䖢%��r��n$��A����U�%Fd{ g�g�G�,��*�a�-\��80����f9�"�5z�u��dn1ؔ��X}<��������SC�x�kﾽR��98��Y�l"�_O��Ż�JF�=���I=��J��e�Cw4`����h	�(n���8�{��tqjrZ�M�����k�������K����������
�D��n�̱��xv���'$��u۠D��z�󄗉 �g�]��f�)F2���9���Y�#��=H+�/6U����q�b����e���x��p���W.��o�5��ux6�9�e̖Zf�t[#��0��\����S9�ὶ2ީa3��*B9�޸�e��'PS��|���֌������FFwi<LD�� �<���ף��_�>�vÞ�<9i�y k� cE��a���CÝH?����1 ��_d���d��������kŠbFo�����b�vO�1+K+����s��ɰs��P���ߜkp�3��!���x���7�~�reT�azF�
�g�
atخ=�Lf�J��}�LM)���m�����Z]���a��"<\RAT(y��B��܅By�>O��������Ŏ00����2����ƅ�΂y��qc�8tP��P�>�ڪE`lcX��A1Pkf�����Ѻ���E�EN��.54�	��d0{�Z�(J��gl:��%�e]�h�W2��o�|S��yą�~'�c=M�TS���V;�����{�1�Oa�tc�C���$"�X���f��D�7��CncnX��8���=�������j���3�{���7νO#�r��+���81.��+)/͞���Z➾�ԷmA81ߔͳ��!-G��3�n�1w�`��f`��tb�Qn�4���|4�b����<�ψ{aM�}�1�cZy<x@sB����a�1�a���c�0��@�����F���q�8<F�4�E��3aoT?H3��i��XO3{U�=�s�此"��cPut�R����x�*6*7Ɓl��ߛ��z�"�Y�.�4ð����f�\(m��VE\�'��#���iۜ��(7n�ü�c��u���F
�����%9��NƵk���"&�% ��(�h7��`��W����z� �/�Χ3�/.�+�q
8I?������I���{����71ӳ��p������(Z��A��+���G��=�/,]_��]+�Qo5¡CG�=τ����k�siU1J�� i�/,�.J���e����㖥�8l��exx~�q'FJ��m	>91����0V���.*A��w�d�4��[�
,z]�r%��g���!�h!s�,� �����T�X��m��C�n(\x�ҕp�r��m�y�)T-�~Ue�x������I��%@ʂû�vR��x��/,�(S�F1����?/l��1֌��!V���l��^N��g���9n�c"W��^X0p�/�����RV?��O�J"�kO�0��q�ҽ9��z���6"=���w�P��*�Ξ���.\oF�E�)���7t���|�y�����j7�阋�P��ꋑ¡r�h��R���?�97�??}挌(�F4�.&hk��̽��y��n�MA���A�!��?q��O<��S�c����ך+�'�[�5�=�B���(g�Z�-{�"� ��0�6�C���>���b
gn��>��#q��:����(d�����z_��x���+h>k|�g����1����b�|�ǝ��7�8C&���a��z�Lw08<��`����s��&�������%Ŧ�s����nZ�~��h�Ep�ԓ,�JF7��>�(��=������5'?�"�E����\2�[}�w;�<���IF��c�v�,��g��p�=��1��~@�8S�[3J�q�M��;w��W_و5;ߞ}j:LU�8��\^Z07;��
�{�7<�g��4���1��U# �{���G��f�޽�����N�:^~�h��D�C��q�?��h��|����W��~C���t#�\鹕�?Fη�4���JDj��H �Z,J��� ���R4��J���(,��S�����vB�3�%-��e�S)�Y�	��J�n`d� ,�L�6�T����:|yޠ���M���Sag�?�S�--@�*GeH���,Ɗ��M4�lB���A��]�h����Y�7�qQؚ���Y�����Y����g4�&�QQ�U�K�MC�g�j '�˅Ր<ϼ"?גq �f`�6S��s�}c̭�Zi#�,-���y�p�&E;1���y~Jy��c�����4�3gτ3��T�ãK���b���sq��x� �W�l�'�>&�cܣ؃����c���d�gu��u3X0?�����'%�8!�Jc���7e��4M�����ʍi�����hм��Q���~9�+�<@m���q�<�Q��|Fx&zӠ%�S��_�L����ҡ�G��{���|�G�ݵc�n�1��z#���ݪ�y��� �fE�G�gg��N���Q2����{�Z������]�?�����LD����2��9Yog.ǥ�8��-�W}�xꉢ�JYՊMM��ׂ{�~PP�`��߽r'[mE����<��xR��bh�#�� �0��ʋ"�ֲ4��秄�Y]]
W�\���&�a���S'O(�s�(%����B� ��/6�Vx��B�X0Fd���')A��Gkdy0%��#��0��}�r�&7f|a�����-Y����;�E���*Z��'�J�7��BX��Ab��(�}�RS����+am0��С��{�x��dZ�f��\���W�`�ݐw:��J't7z�������+,ί|��
�#����5����H�w�bʖ<.�d|�!���|��P��{�Ƚ���}�]p��h���B�p�Z�)��x���W��`�Qa4y</Ɔq�\Hz�yD�{ZQ @�͈�ia�ٸp���#r���H���Y}(g�ȝD5����y��v���A��@�K!�jCaJ�)?x^� �G���O��A܌	!�t��Ƚĭ��M���C�@�c=�ZQE��������{4��r:�t��၇�R@Q�:'�2�u��kc�O����S���7�EEa�~K��B��G��:��QΚ'��s��cr4lm����=�dTH��f1�%ñ��pl�q�y�іb���q�����ת����Gkc=���=�r��CC�D�f��bhe��b���:� v�q�{LQ�zM�X���̐�Xè��*�^i��ר�1*7�{�ek���9
#f������q����DB�P���E����X)g^z��� @쿂=v�RN8�P�`�\�p^M���D`�=Ŵ���ë~�EL
�^�Pd���_����/G'�l8r��Ri�QN*��nzX�K��Dc�4�i��+ˋ��sS�+Y����F��V1L��^�`v�-3jr/������fr-�U��EECs� �o9z�g��D �._�,aJ��"(�^|��m�x_��,�����,��ɸP�x��4Iቫ�q0�^DfP�*K�V�,E@r��6W�lv~�{"��s�=/��Lz o��@�?E*g�#�����.ct���0n�0RXԦo�g!��U�̈́1 ���Q�w 24<� ,QDO�����{���,�T�-^�����VVd�~x��£�����l�Կiǎ����#¯����<�����-�7C�=6�G��cN�Za>6��mæ�Xx?J��B�~�|���7��<v]�V�|��aJӍ[s-Ā�:���;�j��w}���z�3���ov�����Іh��!���+_��*E���{���;��:�1"��eӍ�!�0[��4\��GE»� �Y���i���g�;:n��][9%�a3��sl�G:<�dG�s
7jE��MFgjR�4O�ɐ�:D�����[_���J5�-�I�w��h�t^�Y�w b1�(Q��BQw�6����� �0'�����W��o�n��ϋ��rY3/A4I&�Swr�}�E��d:oˢW�n0w�ԍ��%�9�*{ǌ���g��4��;���Z��|����
tAi�~b�'K�7R�K�.�a���+�:��D&Y��%�q@;����7��p����5�S��]�0���
�^��� ��qK���_�lF����@�8+��!��`����ot^À����)��A� � TANOl�~	�0k/qMr�1q "ccQ	�9����7����E���:k�Ю'&�`�ޣ4�kT�Nu�øb,�3���o��80>g�@�7ClU��3!�Y���ˊB 8��kr��������rPyD9'�p����8��o��h%������=>����T�ː#���������_�A����wP��ݸpa��z�/�߽�܍�q-��Zc�%�3j5R��P����Q�����Ը���'�`c�?C�u��yS4~^7�j���c{��a�T��84�7(4lb���>�� {�4*�	22��}c�����D�����sܷo��%�!���H%�0�Ln�.�UQlez8���}3�c�v�G��q�?�`�n����.j;����ӄ|�w�(�����W��q��A�b�*z�n������g��}HM-�xa��V�����a��s���d�Q���C�7ҵ��#m���	�z�;tB�o�/?>��FyoF�T�Hi��e�HrN򱴪�V���:r"�QRCe0��b*�8?n\��9�5r���0�U��3�9��0�����A���O1$�3�1���b�~G�����&;7��q�ui�zt:ߨd�ɛ$S{�1m)=�p=�s`=�0�ji�����ߡ�i� �6���=UQ��{�����@=��&,��</�Aꦥ\a/\8A��#)-a����(�^-�ݽ$|h��h8P��^�#C^�kx��`$H1�&#���W��+av�\8v�����v�is�'Z���΅�9n����=`3�\W���_���VM.���oT`r����y��p��+�o��?�Ϳ�B��F�(�s��ń �>1*p(9ܫ������̋��w���uDQ"6$F%��{\�﹭J��T��^%U��M=YNJ��� ���������k���zճ��T�e��\0���͎q�/O-��Z*��j�m��pC<ϟ��������=�*�Z�x|+�r�7H��r��1Xl��a�z��԰��	y�F�(H��@��Y�?ρgO$�(#�*7dhn��ycf�������������D/Q@9I���!�����јZͽ�ty�k�/]�m�w�Cg��e�#7<�2B�1�M��]]��8#f�X1b>��	�������RvP���%�Ҩ5*��0�w��R�ߍJR'��?��j_�8C%�>�я�s;QE+
١�;c�T/2����@�iY��|��������+B��茿�c3:����˸�NC��<Z.y��gq��)�T�-��2�}�}E�֓CO��2E�H�#��s����P�M��3&�0{�{"RnFK-�h7[���r5eC�����mDۋh��ʚEYʞ�����щ�������aie9��Z}�&L�v�񼓨Tj�t�S�xm;Y�M��sƴ'�ԤP�k�e�^S?��y�b�V#oB��y�÷tzU��q�^�=��I�F�x�gp ��{��n����Q�\���e�c�� !7z]`P���-��r���|s��h�}T)��c�7H$��"�� f�q �E��`��}��_UJ`R��[gq�I}<����o�A�!J�_�m2@i��-t^�������������w��fܺ�X��D��LMMH�r}�o��e�|%��Z�W��_V���4�����y+s8z�U�7z��N9�|{��`=�`\aWqݪ�X��ǎQ�m]s뉍�Rs�uk�WW�|U�R��h(r�N�$a8�׼�=H,���j�uB���8'I��U��E	e�wFy�j�ŗ�/�s~֍+(<X�ι�ܯ^�굫���p�+q���8�(	�s����`�(C��s�FJ��ǥ���.)�p#�����=� ;�&�o��oj�3�8�R�eעz��<}0tR�E�tꉧqT�J=1�%��S½}�k[){R 3;f¿�?#|�_|*?v\�VJ��f�J�{m�o�&��sw��0��o����(�ˉ"}��n�{d!C�@:��6���j4��:KSyH����īTY�7X�WT�;H �^�c,4̠���Z��πf�j���9nό�`��!���}�K��M���`@l�f�Ko`�j��X�.�g�f�P�Z�553�j*�U�|����5|�?�(P!M?F�u��
��F������Ø�S�>�6,]"(<�];wǅ��J@��)H��A�54�V��5:��5��+Z|p���X˼������/xx�P\�����_��2LL���m��L�'�Z�܄��H��Ln,��c��L7��mw�ݰyu����ks�sa��}z�T 
@'ʈ�
F��]i�N7( �#m����~H�a)T+ h�6�Gj2l��O�<1T%�C�5H84V���i��|�r�/�j�̠��>no�x����s���|��˜+����#{�Z�����u"6⩉�O=���Lp7���MX�Û�Z��x^K���V1�V�(�a$Ƌ+Co��
��n复*RCԆ�IIay�K: ���yy��T�^�Gu1jPJ|a�F�չ���Ｎ=�cю���P:��-�?�H8x�N1~���	˫���U���I>�6Uxy�֟�0ZUV�O���;�!�&��Kk�QED}ai������zz��i"�V]��Tà����Y���j��WѤ�J{��uU��*��R_�P�4�� �}ɛ3gO�V��x��� ujF끱����^u�od��Ӫ��= �(��y���z�c��Ũq�|�=�U���gÇ?�a�ؐ�<�}�C����K����Z�9�p�4�'�}m ���u�ⷛ�8~��>Z
���LP�*iuy��Vd�@$9�R&DY�ୁ��H�]J{�^9]q���*+�����@���B8�Ͱ���I�S
��v���0Ui�Hs��!���fʑ���w���=N�87�U#,����Eҕ�lǍv�RX�F��[�f��������Շ�]������;b�2)�{��W↤c����>��-Q�h؂
fw��������V����5���Q�oe��)��#t��+P(N�/�_2f��X�HB�6ldB��*%���P0��{*��*Rc��cl6�T��Kn������y˽���B�9	{71c����ױ:zOW�J`��9��/덨�ŋTF���g�	�D�|�n��0�������4Ji=^�U�\����&9ʁ�V���{������v܀�+���X�-R��7@�(W>��PZb��1� ���Z�pb(Fx��w��k�����bY\Zܜ޳[�9{���u H����2%���l"��A���k�Q��x�x}A�~���f�$?����y(*�f4d�i �P]X_����_�����@|��W^/���UҨ�s�u�w��y��9���!�Q��?����O�E�V�eq���I!XJ>�F��.��B�A�^L_��cmad�&%�3F���'6��|^F#d>^�_��_��s�9�=�s}�ē?�d�W��_��#k���g������7U�g������b3�ל��|(
������'�7��w���N+ H��.]�V�������1����d� �0��1v��b�@ɰ�N�>#]�,��)+,��X�	����%���ۻ���8n9���x���w?fR�H�juLL�Q@׭�d�h���f��Xa�a��A(�7�D��ffw�t��(Mx�	���бq�5݀��쳸�u�M�WՉ�d�M3��JV����y<R3:�k�r鹧�n=�|�k���A�^��`���O��*�����)���稱����\��c�kB���*�W���AX����h<�457ބI)�Q�]��z�<h�a>����w�TZ|J�C̕����,LUF,ŵNzi2*�/�K2h�A���aE�������6����[�M�lQ*���"|^<�C����씗�[՟�m�V�����|���s��c�l��XIX3�;J��o��]���ʊ�ep9�+r'����!�.����8r���;#l��U������V���+��G-����F�¯�گi܆?�%�	�46�	���Ɵ���W��V��F#.s9���%>�	��)d-4
_��W������!�r�����~��ͭ��I�}'�c��QY�󼢳��#qPF�~H9���9=��
̏,E�	�S@�Fkk[�}�SEd�^��q�2ڍ2������|��/��ƙS#�^�"XS�m����3��as�z ���0�>�я�_��_S<����Kw�؅�K�T4ܯ^�"��Z�[���WC�,*}���|�i%�xtl���J��,"��ލ��9��%��F��ݍzS��F�լ� >�Z��bo �ᅥ��;�<gש	*9����;����Ik��|�d� �[��F=R��-h[���/�8�x-,8ZPp,&
��� X�|G\5��G���'^{M����@ޤ�0�a6�oƄ qtz�0��0��9
T50�O���`M�2&�����\���Y،�ƌ�v�L��� ��9����'���*O��$@bY�*��y?���x�;���U �[WlUn6�Bz/7��jU�ѵ��F	���qsR	�0db��%���s�j�;�E��^���;�o�"��z��P�8 ��\�|4^V�g����O|\�I���a� t�f�[G����u���Y��9^�w�'���Ԭ�|O��R����<�D�ȳI�����?�� ���y������=cW�2D��L�ǝ�p�����R�Ґ��s���3�|/|3�V�{4�a�&��ܒZ>��"�Ic�\a�c��[1�}�U4 `��s�C<<Dl��z����#�1<OZ�` �"�v3���9F
ʚ��O>�d8?M|m}ٽ\J�o���?*6Z�#�)G��;*�G�
�[���iF�2�R�����
;S�=�x���Ut�(	�	>���̉�Xk�z����:�T�T4Z�{��g�g2r��S�;~} -�o�6�ȏ̓=k�|�6El�y�qoE^���/Y�c�X1�_��Oˠq���<|X���|���@}@{㜈�c�=.c���Z_����� �T�;�����4�Nˆ��<_KΞ�Vl����!URF|���"N1��A�JN�V�{�a�_[_	�����{³Ͽ._~!�oC�ϰ�h�����x2<��w��3��{�LQۭ����-��n!�`���.��~��?���/��r���Sʟ���~F�&����P�!5"9+s�:ו��À�تk�����X���햛�B����a�A��>//���#a��C��k���I����r�p�#��#n'��h�`T1��Ҹ��s��ow����a���O��U�o�3q�8�	߄�=��h�j�vQm�ͷ�8�� ra�=�����6��=�<o^�����h���s\X?����k�Ŋ����<�n��Ri6&dxPI֋� �Fa�֭z;4i��o�ԙ�\Q�ν{�P;
	^��!akDy��Ű8��*B�N7�'҉�@�����=zZ�s��*��#���O6R��*-Od{�F���6wT�;�ˍ��7I�6L��Om��o�B�.�)�a�h�]̨yS@U�v{:=vw�x�Rx=*��;fu���E��`�Pp/'�t��Ud��������}1o`H�)����dl��T�f9fN4��:����3|��PD���,-�肘ԫ��:9t�@�����������Ξ;w���T	iڮ� ��
rR���G�M�iᙁ���!u��3��QCԋ��00�2w�w�Q4���G�"S��`]�������xVl���,z\A0t���[��o	�5O0�s;g���k������#����}���R;�V]M��_)���]R݃r�ӓ;aǎ�<Q��%�����>�V6;��!q��!�#�.�^�,���}���a@s�}��0۫����wHG)
RXq}�k1���a`��å�y��5~��pþ�~Bȍ��W4�)���3	�O��Ű���sߢ�Q.�&�jX�~!��~����w^m
F��Sa���<���ZG늽O4H�,��P�c�|c�o�^��+��r��֔/��ؤT�M�J��c�u�	h����g6)�<7ɑ��9Χ����觪��(�@p[�2OI���U��C쌉1R��Q�DN�V6��i\Έ�(|<,y�a3N��s�e֧�,+��v��U)�C�M7jn&�o|������7���ʅ�u�H����X�`tδ�-�ls�w���{	hn،�����l�������u��\H嫝D*�$e��!р�3ަETܳQ��c�r�t�'}�(ޭ�����7���h����avvR@��V�hg�A+T�x���(����r��^�+� �b"?S�T��B��-�?�&���3���TXK�I����8�z/~��OF�^H�˂���yH�FB��ZJ�6d����sG���|�c����D2FK�+W��]s��̩a!z���)E_O�0���4>�햵�hS�0�ss;*CEt��iy�^���Z��~a͒�}�V³��D��x�x�"7��"Z��y#�K�
�Í*�}� "
�A�k�z��I���Kq}��]zΩ��""F�PSJ�tXH�slM�����x�Z26�W��#��C��u�$�,:��̬��u�πG�C��U2h����ޭy#�j���b�wc�jHq����~rn� �0�� k�?��1���O�T�"k<i�l���q0p0}���S�kb�䑇d��)X�J�=�!�y��1*��W1b��z�F��)	|F�>*�>�l`�̻7'f|\��7_�s�� N/���0�7[a�Bd���w����cg#9S5�T�t����c�ˌ#@+����᳙}�As�U����<O���TX�(�G�I�Lf�t���M��۱s�8���	ɫ|͌ �BW	l�[��9g�zGU �`ag7�\���_�` (M���AP�����w���X6y.E_116-6(�`��0j�O�͌�Q�ƣ=���j�!dƚy6y�gv"�&�a��AS偐�t�[���!�bq8��Cw��?	�fR�F^�rU�?�bF��+*�k��� ~O4�Ge� ��0/c���ѫE�
�@ͅ��ݴJ�i�wk2�߽֖�Z�H�Q�4���Y\o���*
�����Y�:Y��X���X����j���u�F����L+�B�Pt���/	�v4�(�%�?�x^y��?[�w��hH]Z�V�ek�Q�{�+*������� H�q���w�١
L"�f.]��X݈��!�)3�į���ݫ�A��7���M%�[����RXJ�j"�8��	�����H"Qf��i�Z�dlD[�����'
���_�=�\��׾������JUb�!s��U`A�V���jAc�E�"��NI<2��Y��8]����j��N��h���(����� ���s?p�����7M�cd�ͤʭ1� ��կ���� K�d�w6�
� ����#�<G�j��^����4Y^ui}��*L!�7��x4"�s�P���A�K����)-R���������a�l$bAoi��6羛00��!�h,���(��R8E<�&�nq����l|��K�a��i����W��;��q[��rC���\�76mV(z����s�%v�b$��s,x6&�����:�i˭�Ъ�:����$��x�:�v2͝�A�EB 1V���k	��`?T9���
�v)OW�A�.�A��	����4���1�v�??Π��؇B��2^��GP�����G�����S7�Χ�p���@ļ<;��9�͸T�1�Z�o������%���S����ך]�~-
�u�<�g�d�@�2��'.���`��EON�Cw
S/���{���yY�(����SB����P�6�Q3f&�JY��,��	?sq=�L΄v���6���v-L�L����k!L�gC'�wmc���7Z������F��� �R.�`[!h<9H}�,o�Ua��/�z�;���)ǝҊ�i��U�uM��Z�eM�e��L���������h����3�,]��:َ^�TKsq��ǣ�rUX9��8xPB�T�%U���ǎ�)=������e`F�~�T�������/	
�+c�S�6<J�a]��+餿��oS�F"�A���BA���c����c0h>��S�g��?_z�eq	��7�����j{B�#�������nsS2�:��D��mi�x��܉�
3>����g��c,I�l�+�;�B�謫�����S�r3e�ƃ�I�σ1�9慨����p�ԉ�r�:�u�h�#�g�����ܞ��۝�H��0>3��9f)bŞ���Ta�r���eP�Ew�|����0�1����O��d��s�@���j�?癉\ob@��RqF�4ܞ�j]!���g��7���p�je*x������X���[߭8n�Q�{�N��q��h'�録>i�1<��|�Cj�X80h�6����Q)d��� Z��u��(�k�_��U/]I��<�������>��.������n9i��7G2��1��b��8�$��뙗n�,�[�[.D|����q�ZQxھ���߷��G��L���کo�칱��V;�\���B�f)5�D /.g
��{��p��{�U�������?~_��_�l��G\k2���`���ڷ��W����ط7Y{���w�
�g�{F�ٍ�Q�/ ���b**�h�~4H�V��R4� ;��ЮGû_����w���ep��Pڈ���Lx�P)+����J	LD㻳!���j
ɸ�}����*̽0H�%/{zzV{
�X`q��T3!-mjPQZ��-��j�T��MCt��;a�����
xljqo��ڍ��0�Bh�q0|������8V������qC�K��(1;�#:2]y�ȁ�'N*26�?�e��'e|�������o;X��f�d���ԤE��,�Z�$}3@Gϼ]�r9q��1g͝��<�}�c�?���Ar�۫�F����J�c��`i*�E#�s"_݃��4P����Q�&Gi��h�aüz��D�]����_����<��?8���"�Tb�9�1��a,Ťi''�A��h�s�A�!ҴDJ<�1�c6���"�G�:���
�\>�Lpc�sx���C�:c�:���i-!�4�{�R��b���?��X����g���plD��=���7��\wmu�:��߮�}36�J,�㬲�iHUZ��X(���zK�h9�xMt&z)⴮���1n�q�#5L$����<-��@4�x�	;lBf�Y�n��0?�#�s���u�n����Q��ٻ{OسwOX�v� ���O�UBt����F�7�aQ���y{UQ�J�%�����;<�����{,��R=>�@a=?���=7`sF��$�|5�O��i��ÍǕ���gG��Maذ��ո�=��_��������|3���^��kUjt�|��3�bp�9@��~�6V?�3?�1	/��?���'ٳ�$<X�ʁ;�0~�Zv� �^Z^�UU�C�g��5�ʊ��7��/�76��s��.�`O���������*����l�>�^�QRDS,<X1�����0
�Yk��#���̬x1�H����J����T��b�M��T}F*U���N��hܡh����9:�p���9��h�|�ہ���~ �ij�-���ј�����{\%ZI���\��Tա�̳�� \V�?�AES���:u����e4j�W��`��M���&�+�Yx�b��(�p���O|2|泟�3���C�V��!zK8Q���a5��GDڙq����Ԕ�� ��ZN-8<h�$��%��>��������1/�O�T��J�����3o�>x�r���X��fu��30d�������ȩB�ِC�N[./��A|+Q���,�S���>�S�
_��/��^yU���c�^A�0�ɩ�bs1��ԓae�vP$òE�^�><X�o?��*�9J��;c�i}������T2p`$}�e� �ic�o1��y�VC{���1�h���u��e���T p��5�ܨ�+h\�{�i'�
B����5',�y%�[y�|֙E"G8-=�������B��TS��� �F-���G�@���L������*�F�n��<lzﱤ�o��s�xy��#`jŐ�!O����	��
勳hZ�ʓ�#��4)<��]�~#Ng\�v;|�+�����q��xzp�A5FXT�����1>��
 ����a�=�3lF/aƊTz���s�bL%��MR¯�&F�^�v�f�G�D��'iL���P��u����Y�k���S��UW猵�aE���81b.�A����n����3J�!��p}�zF5��t�)2![_��h`�Q�6�P�c�� ����9���]W�ְ�o�w5o�@�<`���;==����q�Oڀ4sѳʜ��~���T{Bc�h�ru>�F�K�KT��'Upr�+H�Z�YÛe����u�>V[�M�ʴF����*J,[��^(�F:�0C��g����nK�c(c���|��͡�41z���ܳ���b�56�a���j��zY?����5(>�l�9�
Q�M�5�x��P����s�[[�ø �c��% + U��9����X_�Y�����E͈ܴR�ܸ4Mn0^��wa�&�����O�������^Q��ǎ��zH�]��l&�0� ���P?+�m
���U����1=� ،�)R� �ȉV�S
n\�!_Sy�Ϟ���Q��Wк,�ϔ	'�
����U�:a��4�)8(��Cp��)$�t2�n?�F�m�~�	u��	#�n�J�4	�X==��s��2�1z��+Ǡ�F��g���u�?�@$gA�ܙ��c_�g�JI��~��=���D�8��1C��r��U��{l(��ظ��|�H�8Q�m����@�6FZe��2p�}�}9�4.O�;�1ॗ��W���r9��7�Q#$7L}�">�9�77F#�Ȃ��zv/]���0��1[Dl�
6�&��9���A���񾑰dO�=�~����k�Q�N��9�9(J�����l(Q~ⴘT%�s:^�L�f��I:�A!�bOac�ЗgC�e�T�:��޺�����K�Z�hK4�k���N�Њ��>���B�IO6㽷�^����?��1W��,F&\�/T����2*���)����.�	w�x�����:11{J��ٰw���s�����D����D��Q�޵SϞ�¿p�Mu5&:��{QMDI��ն�x}m5��y��n������yf�����;*�S42�#�A(k����F�["!(R�4��q~���^B
{�\:r������Wح�N��R�HL������i[���g��T�#�T��#�Y'Ǣ! �G����$�r��j_������GtE�l�	3���j~�hllll�C�
���iÿ������C^�O���Y�t�:O�HY3�G6�6������J#�}�=R?���;Ϝ��l�R3�U����� ��0b��,EEe;�wC��i9h�V���{_s��Y����{�^�2>Z�*���5�er��>�r����a�n9$8'���v�#dL�}k8�"5�U˔f�m��0ü���J�U`�B�p~(����L��9-r^���b����mf�5��"�Ε�F�"FSS����\j�B:s�JA��@�Õ�q�}� O��}�K_�y��vÅ2MʲY���.˫�>�� Z/�2��x<�oVt��[��\�J(�v����#�j^�<
�)l[lN3����#�{޵�So�~n��/��T�1b��z+�s��=j$����	|���k\�����8N�q����*o���r\�Ki=zD�����y���=Ǐ�G}$��ß��(@����#j�'��8�]���s���h���o���Qp.��=��,&+
�B�G���ʲ��ӫ���X.�l��Յp���}.8��`��DC��4*�BY�
��=�|_�s7aK�}5�㚌0^����-�n����'�Q�{����6:(�f����G%�{��@o���?��~=��JT�����Z�NS�U��~!�_]��[)���U�4'��<�@Kb����h̨2�J����#A�AA~�~���Ь��|���̳��00���k"_ˮ��]��1��~�7~=\�zMD�^Mɿ0{)'p#�Y�ѡ�ac����;m������bԠPQ����41Dԓ�拻v�=J�E2zS�������0��G��	��"
���DS�|�a��0�!�*���5�ּ �5���;��8��Xp�@�#)�J�$Jd.�F��h�,5k}��dO0^k]�'�x�.]���zAy�<g~��sJ�}�[�Қw��%����������2��D8��SSS�#IχsR�������|>q<�R=+�<[���*ݺo��R�(ꀥ�
:�i���e圆�~�r���cW�,�Ec��!�[������2��}ӻA���y��N�yG��(A���g�l�~��4�h�\����(� ��r�X�:\3�S��8����ǽ��XB���ڛ��c�ϣ$Eb���k�$�ǅS�.A���]�ʰ<EDʛ��7Q�����^��/OG˲�*�_'�1��~.nnh�K�������A�x&�t��'Ս�q����H��������WZe�c��.^"�f>�����#ѰeNϞ=������`�z�Z8w��p��I���p!C�cH{슊i'|&;w�<ҽ�S�N���:"��5<D�Y����]��N�>�{e�xi!\_XQ��+<�l$�TC� �����m�_�S�}}e5��`4�bd�;9(%H�87%��
˞:m3����z�bZ�u�H��sT�x:����Ҍ��f�t�t�����������D{*�y����ܴν����,+¢SXk7�׭���XY\2z��q��k_���qx��g��ˡ�E��בGS�ߚ��޽�������b,��땔"�g��z�5�K����2�&ֆW����)�Ѵ�3��C�%'��R���M㊘WԜv9�C��H�3.�9��aV�d�GgwY���2ݍ_�:���@�����*���<�c<�)E"&C.3cW��,����e��T��ɟ����p0�3W̤`0�qBh'�?���I�š�pt��/��/����+�eﾽ���(j�w�=����`L8�W�9k'�@^�ݶ��;�v���	a��n���mG�Ս�^G��M�rd��ժ	�G��fQ5,�H"%x���k�1�$�t�e�Ni*[�eC�!mh���'�;�:�<'�˕�h��*�nmƧ��b��MF#�y���Vǌ*[�<�k�_�_�k6*,h/9��L��~�
)ִ��c�0�K)��%kU��a1�9�/~�>\�}�G���4�6)��C#�����k�{��p�LR'�������$
 ��q{Xڄ*���ڹc�x�V�V���<q��huY1(��nD/�	�3m���H�1H�y�}�ɏj�SJy�)�y^0��>gP���*}����c��98k3*���
�?�?�|�����Y���<*��	��zR�~�W�I�=���sGْ�X�_TY,���d[�<�2zɏ�ȣa��T�K�wꍖ�6pZH{�s��z4Z�mU��9s!<��+an��x�E.xf�.��t�jCE�wG�;�1���2Vk��7,RQ��J��µ�)𮩊�.�x�X�*��FgEe�q>�{~
k�1�**�� *��L7"8x���V����7Ë/�`XR~��R��>k�^z���㼌WL��t�O�~�k���ԕNo�S'O�����V}����˭a\�k�F���[FjX�GS@8}�����o�����Z���rE�C���/�E�u����~�M)ok�wܨ�"�#�6�[�{/.���r���W^IF��vz%��Fc>K�Յ��������<��3ZC���e| ��� ��E��g��R�8�!43�-ƌ�	��c�gID������yi���1��� �<`~��Թ|!������^�G��uQ�O}�)�$�}2F��/��2~�C�����{h�&�G0`�ѭ���R������L� �F�x�v�:�E�'���k/O=�Ǝ�E
;�1ɫ�`�-�cR�;��эχy�F�m����Ϭk�_ֶâ6���m]�ݣ���<��br�St�+6)`ΣpL���'���m��u�vD�_����0�X/?�sWST�{��>�'\�x>�j��'K�Y/�{F��R�v~%M��&���)k۰��Mp��%-\6�7NۜӴ�Ç~�x�����e����kj�v,6���13�M^R.*x���pa3񷑍�$�?��+j ���ã`�#'��x⃏+?� ��?�7�KJ�]X,%`�����0���!!�z�"������Ƃ@Fq Mn��������10a�n$%���1��ζe�J۽��.�h��d����Xa��ak���_���ף�XϿ�!�v�HG/,|S�z��)��`�7���Li�1%�j�`�m-Q�c�\j]	��s_8v�������g$5*���Pt$l$9�*���@�feҍ�3̭3`+����M����{�1���2�1AW�&��)��aF��:�;e��.{4�������Op�4ʾ�����X�x�>�9�ǖ�B�ǟ�5*�(��5�+�JT����skZS���*>�+e-�F�|eM)<Nگ�|�G�����;nZO����Zꥡq�� M�� wc�f��=�Q�<�dk���a�NW�ð����Ξ���<���y���]Ϗ;�����S�uS�����p�.Y����?)����<(�z!H3�9{6|��_S�#���W�?���ի���p�ʇ�2�+A�s5��:�vu')-�Mc0׬�ovvZ�{�	gg����.�=�S�έ�_��7wh�2���0/�O�p�H9���vK�{��o��?��^~E���E9xZKK�:G���R:�Yc3�WL�8ynp9�T��,ך6�ng���)�z��0��:�%kJj�*��|���x浞�Wj�so���&��=�p6>��蔶�r>'�1>�Yʐ������-F�����@9{�cC�� -@ҿ��H7��@٨�k{BF͊,Ӎ�E�p�<�p�*�ڮkq�	��b�l41������_��υ�������]"Mu4Ot�f_M�R��A�
2�9�h���#���/��^;�]T}\m$@mZ�z���*�M4�6��!L��FL�V���x���X�(�1�|�Mi*�D�+�Q�7�0M��j�J޻^��,�������Z�~_T��h�-�{�=w����� ׳\,����E�h` YznZ�fK���4y�Ō�BQ `xAt8 W&�A*����s�,�2xP��)���A��Tѕ��u�W��W2�(�V>?aQy��}�꼰;oFco�#u(4z��e*��_5.c\�*Ò�>��R%���t��(����I��sכ�V�����XC���r�w�՚a �����M�,˪��}�sV�<�P�MCC3
5�	^�2ْ�-Y���o�'���?��pXDx�~%Y��d[Fb�n�y�93�r���߳�:w��Y�-���H:��瞳��k?k�g=r.$�ٙy�P9d�]+U(N�ӡ�K�����F*��wG�M��Z��p|�>ʺ�4�H���A#.����Ȝ�W)�9A�d�mzr�|ooț+�B=�p�@bD��5h�����ָϜ��ƐkR�!~ �?�f��v!����h�����\���zt��O�M%�W_}]ߋ��@
'"�υ���HQ�~*�l��c&z��Z���l}�>�������B���Z�R�V�-��U�D�6�7�gy��ڋ��JzKڔWWW4>W#؁Wv�ԙp��M9}|�7����q3�R�-�#t��ڌk���55���s�Ԃ��-�SOsΛ���4�����]�-�C�[З��%��Wm���4��kVn�ޅ�������ڷƩk1�zMh
A/������S���L��Ր����Vq7-0�:m)ҕG-����_�jդ�Z���)�811��I�Y���9��v�h؞��;�f�P}"�f*�	-�=o�����S�g!uX�E$����J�?� �w�u���r�b���p87�I��?Y� ����A&B���s��OF��џ���:^��?yG�ĩ�pt{��W��$�x�K {Z�SRq5�O�C���xK�U*�v���XP��``����w_�J˓���k>�㎜�Ȅ�wmS���B���3o_��e��H����2Rd�\����a�O#x)�;�]����r��Kb�^嗕���Ϊ�{o߾�����q�~��bļ=��D�&�O�MV�S�ra6U�#��F�2�8<G�3�k"�)Q�+�4ɮ��`).S�l��N��7�Z7�,=�%�eD/�v�Rt)�g!u�p_K@A��Ϙ���ı	~�;�5l�h���J��hGtsq9��Ÿ����h<�,����;Vj��+O�1D��nE��*�\���d|�|' t`)aZ4S�j ��Pss�oV��@M�[`�4���J�+C��y�mHů�[��N�1sE�m��������H5Q5[��f�M�Zޝ��.aT����tJ�=\������ԧϓ��u�?��?Q��	��O�ѤGg�:�����������k�j����=��"�����(�c�M�M`'�rH� z>�O�kU�µ�[��y�����e5.�N���l�EkT� φ�C*�7���߸�"@V5	�.U` K�Ru�g�W��+W.k��Ul�'Q\�|�T-m��I�b�}�4�Gr�hJ��!bx!jD
��UENȣ��䐜��~��9�F��l����5��u�Jb� �|/T�wkk�<wY6M�!2���Ρ���XO����}�̙����s�$W��L�S(��]�wxm�"H!R���ո']P���U�^ϨokM9hռ5D����u��	3�a�����6L��Xdl�^�"!�I��n@�Vj~#:�� ��(��ٜ�����3�)�U�JD�<|<][6��٨�Z���S��DO#"xT��Y�|�d�����(	�xa�c�/u��!��}��Wë���{�T�h��8�pt�.7�y�(ρȤ����!,޸q-z,kZLֳ�^rL�%��Ѳxx���x��(�SX�X�0Bh�E��@R?�j��K�#���0��*�:Ec�1�����6}�h0� a�H�z
-��y�g��*��fU �:���q���������	��`z�-���I"yN��ak��R� 	��!(�"p�+�pU�H�z����Dc�E����^�P��8.�Z1@%�j54����'��8"]��r�;J�tXHH��[5�����g�̤� 7c�Xo�o�k�
)w[���o�d��u��&�����b���b�-��W�i_Z:��Bg�<�8/SW�7��R���A%�=K��Tu)������樰{��c>�<?oS@���cM�����T� ��-q�.��A*�t2a�/�N��� �'��紳��� b�6�qC) �`���W^����R��- 23c�8Gl��J�8:�J�H�����Dzͨ��Z;���5�M�nl�NU�^���U�8M�ī��{x�拓��`�pOT���$OG�'~k��������!.�/���K��$N���z��
ػ�|���<�����������/ \�n��v����`�������5�P#cC$�~`��)���|�Os���t=�ΝU?��7M���]�� �/,�I�'�58��7ԋ
s�@U|f����B�Ȝɞ�[;?��?�!)l'��s�͢�a�~���z�ɘ�#�~��9��B�����;
��c0��3S��u���`$�!1ٯ����|+<����]�!�vD��բ>o}N���0��¦��	-_�|EyZ�b�����ĭ oq�Nǉ���UQn�o�Ϳ)Þy��;9�ϫ�Xh�)`������"�9`�;�.\�^}��p��~��e(]���gh)����v=�Z��пI�Q�̫���BU<p�G��k�T(o�H	ߍ�bR��³�~?|���/��g*�Vb�?���zP���Q���.P�5U`��8?�����/Y��dn��������3+�^K�"�%�r�M�R�^	�rLmC18X	�G�r�s#�F�H��ҵ��r^��͵J� ΁�8Kq.޼qC�X�@��<\��H���ķhH�N �c�~�ʯ�R��S��t�����,Pb��x�a������>+�^D9��t|F���C�~˞��94���25R���sˣz����;E<�����#��E �G�<��ĜWsJ�-s8�,6�7�7�I���(�;b�~��~O���|���&��i��~	��������UG1o^�*��^-\a{S��w������_J7
���g�iuO�9_��x#�&�ܯ�Z��"���|�l�kb�roت��u}�7���xm�F�XN��:����g����FyU*��������c<H���
�cֹk�dOR�O�����τ/�����>��u���w�wu��C��Hd���I�}\�u�瘋�
R����Ժ�&��\��(��>�����3\`���J��L�EԲO�\P����>�^����ET*F4.RZ�Rm��̨?=涶�h����o�"7�3
�V���sgdH���DjF�/5�o]�i���&\�`{�̍7���Gr�q��|��<}�� �
����"��""<�G�l���Sz�T���e���×ԯ�IaџIM������xw��ߡJ�&z��?=5��s�{s)|t���]�>�RՑ/�:�	k2�O��?_�җ�Q���A�VYݔ�|���5�0/��UW�O�x�B;�������u!��g��F�+�=���z�$�hϺ�z�T�³PrO!�~�Ӯ�$N��?����q���h����Րs~�-��=��s��;s�TG��\�h�r�5O��w���)�D�݁�wz�����>[��RR����G�r/�4pY��L������囯��P�|�p�N����;�R���jͩp��I)���:%�sj�);C#��s��4V{�:*K�/>_�ѐ@M��e}��wa�!��B�r'#P'rJ9�����K��A�&gg�y" ƙ��d�*u���x9K/�<lk�Rn��a����A!I�q�3[C>����Q��ۨq밬����w��d������?���X��@i��3g�N�~K��(�%�L�l=>�Κ��_��R+�^�w�P4��p�hbS}=����c<'�>@��VE�a6�fft�||ܾ��MJ�~]N)�M��<�]�}[8���E��]t�f�g������>i�'��^�;���U��(���=�[E(�2�P@����mw������@iޮR�F�m��Q�&y|��	͈�H�p�JN^���P����s jh��ÙI3=�9��V>����x-c�=�4[DyR7�MF1�� �p��|㲤���i?K���t����F�����?\|��x==�}�v�gE��T����p0�pߎ�B�	�F��N%�n�<���èL$���P�8�
�O3:��Ʀ�#�ʶt<���4yx����E1)c
��Bܸ5�yϻ�����h�ܬ����I�,x鋥�L
���S*$B�Oݫ1$DX�|7��wl Q�˗��҉�ͽb�0y?4��Q���/�I�£-<��.��X<v���-�����DX�^���._~Cj��� U��vokU �y`<�V��̷(�������S=öSzf�� �{�r���!�m��.�٣S&Ɩpl~8�+?��w~6n^�bE{/���d�!k.e��H4�>;�v}� �\3��:Q��&��:� <WSV��X�D���"/��^��������d���I��xT�J�V�Ӡ~Ǯ;�ݣ*JK�@7x"�E2��~ܐ;UU��&Q{ �x-����_3>sEi�n_k���K�#��A�&���`&e�����KiS
#)�<�����0uἦ�RO��A���s��!��؍k�B�zP��Sl�8 DP��JH ���6�����KD�@�� <Dx�k!G9�k񼤲�5l��Κ�s��o^�)U��ZM��*��'���v��Ŷ���_����;�u��� Ro3�D��b^����|A����o~S+�ҚM��#����;������s�sŁ�������� �H.�Ԃ����@��?���ѥ�-�(�疃tT�S����q�,y����*��4� �S�� P��<��I.���e��:�GSe{�5%5��D�a��aI))����dKLl ��Z2��Z#:ٓ�Ï>r^=ў������sL��g��[PEp�wP��~�� IƟ������t��p/�7kߔ|�3�𶽥��τ_]_���;���-瞚����"@Q��&�437���>��	m�;Ϟ9N�<+���oF��hZ��\�`�6����^��O��5���T�������'������!Jh�`��u�?��&!������RXl��?��05�qQ�|狈臧^�ȃ@��2��2��9'q@���"�X��o���SG׺�F�4�a�R-�AzT��ƬL������(���/�rgϟ5�*�a2�'\���31��3�>����3��%��(���cx/U[D��`�/��Z��������y�7�l�� ��9B)���K���;x���E=oUfu��}NT����f@�N C%�ȉ�f�`��3�7-Ҷ�45��&�MnUO{;{r ���=s�D�d��&~V5��i1�v?�i�iU$4 ��4oB���<���ޠ%����j�`i���N�Li�I�O���C���f}'�P��r-�QNZ�8,����â�yĆg�(szC幍� ,�ؠ����)�6��3�;�y@P��b\5�8 v�sأ�po����/������h&N�~���6� ɏ��6��x}u=>�����;g�Q�6g���US�����?\�9�q�nM�©&�:YX�gN����Ö\����.�A�6��,) �~��㢟�����v��t�˽US3�Ar��\Y^ZV��1��h{�i�$��_���������o��;���Qq� Ό�Y5�ְ�#"�:CNF�@�M���p�|H��B) ��n�}+�%���~C� а�vN)��(G������"c-V�Ѷ#�"u�)Ew�7G��{w��H��4�S1�7/��j���7O66b H�M�囗�P���^�k6.�0���XߚFM�hR�q�OM�TMM��F��W#�ؔ�<Ǡo�V4���(��Bm����Жib0�U�-����E��?�-d��yɴ�o�^���b�a<��+�rP�^?F���^���ܘz�Q	�vI-	�ݼy�ʮ��q�;%�7���*�l���ZU��ZmQ�h*ÍZ��`�F\쌈���lx(z(gN���,e��'B�p����@����D��{Ā�V�Z�i����*!m>��w��v�xl��ߌF�_��e (zN��E���s��~��<:����|��#�ڌ�\9|S&�B$�#[��[K܂VR�'�/D����W�΅͍-)���7���|4~L9:���Iw��0;UG��F����iye��)�YOy���_IiI�s�k�\[5!����u�80Ɯ/�hUU����(��y�����T�e�&�VoS�Q�*���a�g��d�k>W��2n�sP)�?KC�3-#h)�z�NM�F���"ƫ�,��"��x{�۹�$�$��ڳjK�9s��U��u�;N��(���:)����?�h�*G5�-�9Q3�e�v�EJ�񻱵�-oc͆-����>�����;^<aQ�n9N�wr�糱�usS�kSe['�� &~]yz���e��瞈N�?���<���oß�ٟ��m�Vذ�4"�D@���b��T�Z7�@��u O`���1~�{���񴵹���{ ,D�}~wZ�2�̹3��L��E��`�?a�d���J�l_zcj���~���Rآ7�d��HС'��ѥ��#�m@���d��<�.�_�=5f�poɥ��S�^�K�U^]�8���6��-;���ST, ~�p�ܤ{(=��?����ɣ�=h�G(�ZD���i��f�<��G7$��n:�"ǲ���R����S��i8 2�Wn��>&�#��j��빇0r�C�Ɯ�	%^�	a���YPl�xC�u4L!x��*�K�������#�z�ݒ��C��Zoc�{sO?�sO)�"᪸	4��`�%�����OM����IB?iN8����~��Hup���`NP*˽���a` �>�F���u{9�m���+���i)�7�c�yt����p�b�Y�^{�Z,�S�A����T�N����DC��$����^�[�/2�N"؟hTZv��МokS�s���JTfyy]�7oR*���p8T��)��(�
��RزHQ +�ֲ*�4�((�B�|�H!~ �w6Q���$ 
oon���W��M�`<��+��zMQ�\�s+~�Ʀ<vƉJ��)�!��@��u�-��$��f`�9F���O��Áɝ����7?����6��F�Y���������{��.�I���H�L&;���}0oY��el�>�I���uRjw0h���JއG2{R�(-�M��%�����=95l�7n\ Pd=~7߇�{v�����L���@�J�[�v��0r_�rg�!�kt.c%�b�I8DH܎��É�����Z�8�͉�\?��D����#r88��G���D���@{Ʀ��s��w�����?&��Wʯ��<�lzF�VBL���S��;�D֟�B��o�������	�iűvp�vv��k���棑�՛.���^{5:*�w�����������#��r��tDj��k޲�̉��/��e�X_��e�!��i6M�q-H�Y�^�`!�;{N�o֍X(��9J�=��H>�L��p�71*3�����'�E���1$����ϸ���}�r�3��G���R^��0a}A��f 2��YH.�?E�o�\hNX��M�f�V Ǉ>����­�m(^��z1�H 쐞Ԡ���/�@x�0��`�k�\ղ:���]7^�j�;V��J� ����A����7 �{.�Ϲ^�;����)Dԏ�Ԝ�1��;�̥
�0S*)M�P�|x���x�TNa�X��  8�j=0F���V��}����G�U�^q�.^| 5�R��J]�=�w�# ��g:���j��EZ���=U�ݼ�f���a���"�V�Z
�EG��dD3ۻ�I)̳Û�$^�l�z�Q4>ǐn�/�����������H*��h+!s��Sѻ�bq%�=hfvRc����� ��~G����8��/�k.1��4X��\r���Ȉ92DH&dc�W�Zƿ1����|1i�E�)1o\���6D�h�<�"q��r{�$R ����k�bR'�<�"��I��������~�_��1ଈ8���	��ެ�f-P�ZD ��Xv��0DH���Ӝ��3���׿�qQ�^�k�qD��J�'���Ӛz>&q@�<k��׾�u��YO�������]˳�m��J)��cɸ����ߴ.�(�p�h����i��iS6b��MUZX�XD��{����n�]�4sdu3��-~�O�	|�аMɐe���J������{0�B�xzzN�Ѫu�sF����p�݈�Vv17��3'��أ���4x�x9��o�W^Y�%�M��lJUk��r�<ccw?�$Owp����	W�?BJ�:��j�`^����g�����(/����߮]��)���Q�����Q�`�J�F��<�±�x.ć}�D�y�R~�2�����
כK1|��髬N��qQ�/E��g4��ߗG�rP��գbyΰb��+(+`xk{&���M�Ǫ�X ��:=�,{��2Q�S'O+��lL���'�������|H�����U����ɩf��n�ã̈́*�*I��&n��.=,���B��-��UH�2ß���c��6�OG��FvD���}��2LpK��pn�<�F������᳀?ԌG�3�0>.�Ș�2'���*PN*�~�6>62J�-*y\z,E4��z0<���`M����1�!���,�����q�u��h�&�v�ڡ3�����T�3"u����x�h��~���{�>e[d���[PA��Kq� ����wy�fh����Ǎ��k����=O<����M�;m1vI�wã�R��d�r�T�T�aj�jǏ�����d�1��#�׈o�2eqcU�����t=,̝1�O|��d#�X��[[�|�vı�����O�?-ϛN5)fג`s�5xv�s����D��`]1(K����a�f��"�j���8��q��ڲp�~��(E�6Fl�;�9���>ZQ�\%"A���	�4�d�}s��^Qg=ݪ��i�["����Ôk_ �R	��,����=����� ���(��X�9�`��������+�"R�ZM)��T�2��"_��i)z���k�{�����'>�1�����I7�-�?��j���l���T��\Ze��`�pi��gp�������y��;�B����T�-�,�����O�?CYͱѤi9/̳+W��G.�T ��N->�7�"Eǚ���É�|�B\[8_����rk+��c�d�+�g���e9m4�Gu`QZ�24��h��IE�sE���Ka�4aI�+}�V�Ү)��eT=Ĺ��w[(������8�z�`{�3�x�}�� ��>
���/�H��k�`�܃��'�N�<n��������0A/�v�@���B����ga���'�I2y��bp��#4��I~�r.�����������ʸ�����p�~����ލ+�r���LZZ,F��(�԰q�w�yu�s�H�y�R��c�"iK���D�&'�ϐ�-yΐREH��TjQ�Ng/�Ǉ�����6��xd���4�_�Ơ�(� ý.��h�� ��ԧ� ]H�_�/�Es�����{��C��y�2),��C(�H���x#\�q]s{vfJ���P����E!:;��4�gB�1}C���uw74�}-���e�nWQ�$��ڳ��RFX��p���p���p�}���v�z}�*�8+a�$�VkN�<NF������Z
�4k�V-��yϻ�q������NN�%�wky)�-o�GIiR.����:�u�,}/U�ĵ%y� ����������`g�9�j�D&��ə���}�{ףqLgے�#D��
�~��{�]2T�n�d��v˪M��$U)j���H���z���	�$��"&��4�O��p�Ă����f����8���{d�:2V���"K�e�;�I��v9��5��l�����Q���w���'q���Qd�ԼX �\��n��I?�K�+K�U6"�so�H."|�/_����s�~#�˸q��˝��f�F �!هΟ?�5N�����%�������rBx��n���?����@��^|��b�j�wR PS4^��]U��y%��8Y.\8n���xJ�M��b�����#��0G6ªʮ\�����7�|�lg\����w�=M�kL�d.���Ft�B3ܾ�^z����t��$x饗U�XUD����>��ދj���=������y��s���VW���@9E�GWZ0����}q��א~A��Q^S�Ү�v���>x�5)���l���=y���x�Dz�~�g"�Ra<Hm�2�;���ݛU��S�z�j�|W� 6��7�	o�͏p"��ak]��6�aκ������x�lt��@ְ;�sk ���j��U�����4�$mz1���z=b����8�����|<55QF欥D��xv�=��q��E�^�I��$e隆��#i�z�n7TΩ����L��D��P�'�={�.�и7.@�(Ë������N���M�0��_��_՜`Ly�^r����ȍc4&�؜��?��g����=^ӓ�LM���~X[�.�^��,�ҽvXY[	'OI�3>��w�������{#��Y�R�h���C���U����!$n�υ7^z>�ﱇ�S?���ÛW/Р�8P������m4������iiM�R-�+"��\�7^{U��n\�'�τn�mA<���j�ژ��@^#�)�����ѭ�3�bO��8y��q��Q�#UD�:��v��:�sS)���S���/H�.�o���G/���t��.���mZ���� �W����x֬iH��O��,+fB�^%s�5[D��)iSu�w.]����t�+qä�N�Lt��9\��`�7���Aqnksg+!~�<��8=�38J^?,�%X��.S�E,���G6��K������S��T\0���~݇]k~��atz�SO�"�#����H�u����u����͉O<�t��_��=��g,�s��d	 �����i�KF d�InU´:��S�E�|YA�b*���Ee<��2���Am[�T����ޮ�682��� "ED@dNp]���*�E�Hբ�*��� _�r�Ze$��D��1a��J�z,�c�<�zQ��9�)��p(���@���Ý9��Kz&�[�N*'?���4%���CT�X�[*�n�A�����kuU�$nN��$����nm/�a}���&�l��3209�g�"�<�W�ؿ�D|Cg�����ߌ��2v��ADu�ak��8�;|�|���ra�;�7h�4����I�����9��Q�l��*(Re�O��A7\o��r�v�%|�?��?-50|��/�E�r��W�!yK�uq.6��ϧF��Ҩq@&�*�V�|<}h��z������"��v��'R����/��u.�7����Q�^��A����ݿ+�!��E:��lg;^��_����OZ�;�9�*|3T�{�V�]����'5Ǜ�eG JU`հ��'kc@���1�9�~ډ��u*u�0�&�eP��Cdg���q&��z���ӧ�W ?>A�Z�mu���0��*�E��.�
,�hA_ܠ_}�����-�����[sѫ&U������|5��}�:��_�Ui4��Ĺx���uE%욍@I��(7[��Ңo��n|/˲����=���}��t���mmN�����4�[�yCUV3��z�ܜ��� 9%��L���n�W�7�hy�����iUL���2����x�������G�=/��s��O	Te~��U�N�3k�9Ɓ��(9��;<j3xz����N�˫���l�8 ���`+}�G�Y��0��h��Q�&��;�_Ǿ�o7���������hK�}æ�9�sۍK1>8(/���� ҽuU��6���ղ��{��������5m�̮������&�b:4����.;G��x�E�u�5��1��]��"���vQ$_*q걛� V+��8�^�h�1�m��d���r�t{jf����B��S��.��g�¾��H����H?`ps�Ič��ç&,���Rg�M�F
ji��ԅO���������/s�֒���EY�(�2��gM.���D0D�.�x�?��" ٕF��#'6�ސh���{{�'@
F���$��v�0+��)�z@q���	�-�MF��	��-������Qo<�F��D���Ta`r�?"o�Y��W���O����=
��)���8<O�H�^x�<y�U�U��ذ����	�[���nk�>���{Y���j�\��1u=#JS�\<�=h�>Ǽ�=lJ�Ɵk&�@�=��+����#�Ǹ�*�6�/�Q"r���Ѝ��K��0��qj'����ٮ+�:��+��!��6�uT�z��!b6�*�F˞��{��5R}��@�܌������̞�fnv&<p��5���f����ώ�q}���'o\��� |�[*�P�y[T1a0�B���'�bސ�TӼ"t�����k�V��3�f>���N��Z� ��h?���uǚR�{���L_}�:֘��]���@Dx|r��%}z(G���~/�Qe �q�W�C�*�˅cFd^�@rrrZ �4��h�Q�u��3�8E��0�`nvN(�Y촆�&�C�x!jH����_J��-I���^�z�jx�g~&������e��n�l�;�C|'����:�s7j�G�*�&
��>�h��0�Gj�
-���P���h
*�� �����R��s�W[;[�_�� /v.
�%:{��y�� [8V׮�_��_����_輝��!�u�r���l�L���V(����dHy�®Y@���!ǌ9�l��XH���ѩ��^q�Ҙl�R��֚�w#���vjIT-�	��I�މԠ�&0mq\9⺢�\�}�0�=��W�}_�®�3�RM;�N�0Ut�H�G��譬���R�$���&ag�nY��,C=�tm�@�n�V{�K�9�vۦ���6&��wB���^O���r�)Ð��� ��ά]U ��2F�����>�Q�}h��O9^�W��m�J�{�P�?A�Æ���{I��(PS�����S�A����VT��ioN�$Y����)	:��(�ô�'U�&��׽7�#�9�q�^c�3~N�5�ݏ~���&b7�2A�U�	}�:�ȫ���t�Z�F������?e���y��8Q>;U+�����RF H�Mx�D6(������k̽E�Gt<:���$`�S}���ߌ�K� ��5���-Q��ʥ����ܙs� ��t'��w����ޔq���-��f�WV�y{
���xQzI;�h5�jc�ĿQ岿��V����L�L*�S���,����v�������ڱ���*ja?~n2���D-!|��R�c+η��ZV�L�b�HJ���/"�J����`�ɉ�݋G'@^k�@US��D|�D��#���<q:?qJ�kt<�$�+�����$�������9?��\��ݸv�$z�/cIB�fS�.����+�^�A�J�(nã�Jq,D�j{�>iq~��D�Q��ۊ8%"%�󱶱&29Ѷw=��2�}X�(/>ȏq<������W9r�2%��5����0��g�������X��:UBkYN�@�6�0��ۿ�B/��ɞ�r�r���l��X�w��q���^���c�)Z�:I���.��׼��L�m�Ͻ�Dn�]�W-$�j�P��كj�1�-�&�=~��"ͤ=�����wV�3_-��r�E�GR�`G�9?��k��`�����w��D�c��\�oٵQ<U�� ������@p2�@;��G��d�ĵ7$�N��0�m����nn�� u�eâbg��-]��?���||���'>��<��\�_~�Z����>G���J�7��`c ���hAR��`@`\�|�x�amG�㼔<��Pqz+�f��ϦD�*���'т����_�{0D9<�v�v�! �����a\h7KeT��I�BhZ_OBwVn̂]����T�im�hpM��W���C` ����`�{� �|����x�,L����Qv.A�G����wt�\s�{�HQP��*ROT*�č}cc5z�'D��Ce��c�������V�o��<�I ��Ӥ�@D�t�2A��v/E �b ���	��P�ë�5��n-���cDx(3����JJ������Lp��霤��#߯ƍ�IUϼ��E�&�81ی $�yw�2m�C�A[^_�o� Q0�҃�*�Z3ފU~P��h��D¬L�v��\��s�!�0�g=���8w�m��2�����x�;���1��]/��bx����|�x���g�h��� ܶ�'iy�*�E� �fU���G�n�{U��.�����N5ںK�<^~�����*g�{�y4y�]=��x�vܑ�;}�a�a��d~*�<��Wl�{F�N)8����p���#9��5����0��X�8�7�SL���MoY�D^պ%�G4�L�|9���+ꞎ���[UM��,�����M��2_�(�� 7ä�/6]����0Td���䷓0�l�g���~U�͡�{���yќ�lN��}�q�O��}�;��
_lg+�m�����H�P�!��XUr,�
Z�|��瑚jR�u�(��B���\7ě�£Z���Nk�I��ͪ����f�2d`�T��'�Cx�$F������*Z��n��/ {:ǣ1b��59 s��QB��]\�X�>  ��IDAT��WI����Q�H����~�f�@���-�'��]x���@���!E�\�qY^����8�����k�|;^���*-|:�=��^��_\�7��)�j�c<f�F�����O�#�q@��#W=��T��.��	�a^�>s��$�~�>�Ƞ���������(�r� &&&�t�3t!:O��;��}s��� �F��_����- ��?���\����|�z�����>����� |p^�z�?�ϝ9m����o�ZV7�O�3"�_���^�.)��Օpc��Ā���\(���d��v�Ʌcqc�7�h���/6�s����+W�l�lG��C�[5L�υ�~,�<s.��7���5�O��������RMk��*9@I�o�d�j3�*�j}BQ�n�����q$"�iNυ
���5D������JHWV7��ڕ�pr>���J��.k�S���Cv���^��q�������
z�T�~��g�y6���Q}���Ƕ'���[��$H_c��K<����e��#��b��)f��J�i=\�(�z�;�D��o8GpE�]�� I�qͼs��=�x��w���s���6�1$b�M{�	ȣ��r�y�s��î��̺����}�c"̼F�LQJ��Hz8t3����_�I��G?��r�����淢}���jSf�~�UF/��ě5SKH��Ǌ�$�:�Σ��T�_��`�o�U�������3�U[�r�6֍j��#�����g�h���?�41'ݝcE��DT����%rJ\��~�����87o\�4w��n`>ܷ�ރ�D���`��>�{�RZ��A��Ᲊ��6VU�8:���瑰V$�+�����)49�mUXC���C���Yմ�ySG���H�tb��9��S��z��h�������--W�eb2�}<|� l��!�w *@տ���،��T�G��T�g�x���S_�ғw�^X��"P=�G-C�m��v�S�݇���*?�kL��<b'.	[U��6;�jɹ�2i�6>C�Ɵ�ԍ�7"��(��A��z!<CΉX���g	a�>- N��T	 ����&�������-����n�p��PG�<���b0Q"0z�ʉ��]�]*��=��g�?�QX��R�ko^�<��6e��ޮ��MKGeZ��ͅ�SO�nآ[u|~��&���]�k�VhI�� �r���*��?vB����~J��������
�����[�vH�k:��ˠ�� T�M]��J�}��=���D�����K0!{T�'���Wt�N�{k���[]݌�f�:���p�"��Ź�L���ͺ���. ���o(
L%���������fh���<z����ZU_7SK�'J����s��믿�� MA��jŔZ�<��ZJ�x���Jr	�:NW�@9ώ!�����υE�ƍ�_+�nǍ������W����8jӿ�kF=��0*�6�6��^2�2z'v�5���n� �ƪ��w�(Br�M�g��Qu�^�k��1� ��S�P��(�j���n�����"i˸s����{��R�ֆ��Sϳv�J�<�!�&��T��zM뵟z���f��y{�9� 1Z�1��*-�~nuW�﫷U�8H8��o <)T��ף��/*�`t���O��=oh9J\󨇿ο�n���&����>,p 
��D�T�~���
���#�B1�l���'�Xޚ=	J���Jy�h�6�Vj����)�x0��/�$��QLr�¿i����$����<<�N�D����밅{9����������ٹ������ �)��:��,.�І.O �g��UY^��Lpr���ȅW����Ȁ^Ue@��%;��ٳ�J�0��uoml*�Eo��~��'�����?P��+H� O/�M�C�/��� �����_�%U��ab��+1����ɿ��D *H�4�c7����ߧ�?��K_�Rx����k j�50��ڈ��7^���pI�qc�ty�}U�E�(��*�Z[�ak��̍��"�y���q����A�#jS�H��y��n8�ԁ7��h�._���]"k��;6n//��@�yTQ��]��~Q1�H���^0ON,`eYR:V�^�/�M�2\I8T��k�����ܡh�9<M�24;���ߦ�h�������Ub��95�&�o^�������eW��K��K�n7����uj��Z��+L;>��[��~���ڛ��r�Bvd?�K�I�iC�CTG:�� rpՀNP�4��Wn�$�j���F-��v��]m��h� p����V���8{0��Q�������ΛG4��}s��P�!�Y�ۗ���԰�?w��̈́����ݶ�N'��6�g�_���sM�20�8�8"�'�t����P��Z��=�4���G#7�D�4���a`s�Շ.R'n�D�G�M`f���<m��v*�Op#���5�M@�Hq���2,ث���A�E�������|�����E#��_�p��^�����1�_H.*g}}�R)������rD�kKO"����caH*@��\T�7*^�&�	�K$�'0a�n
׆�rr�w��\5�^)fUCh� FѰ<�M�Ƥ|�����"�X���TP�]�.��/��0���~n4���s#�ey��񙬹q[����.."� �<�������P�Y=oL��D���;�/���*�B��1��͔�`b��v%���\����R�R׽�Zi` $��q����UK#�3�9 �'?�I�}��������SOic|�ᇤ�C�G�\ch��M:���?3��� ����4�����}H�I�9�g��j.�Wd^Y�[�j�����Rx�}OJQ��v��.����T=��R�^��oa� 6���D�k���7�T������ގ�kw��R��˕��zKE`(�p��5VT�ҟ8��plv!|੏���k����;j��g'����'�����*�Ž])3Ɓ�ʵ�*�(�_ZYז�����OM����.PQ�f}h䴑W&�8h��C�w�r\��Ao�˪�|m�ech��y�Ժ��=ި@#��=9�Y��.iq��J]e� ��֞5�$���yM\��
�@I"!]J=z&�w0x'@'?۝>=j�����6 igAE �[W�/S�����ߛWA�s�?@��v`Mw{i�_p, `ED?8LAހ+�����| !�|:[Û���p�xރ0(�	 _�*��`��:�'�#X;(S3�Q�w�Ph���6e3q�Z����N%��A��RJ+�Z�����MW-JT��7$4'(�H{�OV��pC�5FJ9�8����jU��2�v�Bw�275]�+U�\�)�-<�#��b��M+�󾵓5�'�b�C�⇊�^�!S�
��&��;�M؈��vD��>�$A������hj�����y��������c����x=��ۿmi���)�e�60b�߯���RQ�O���pZ����[��RFc:)\��~xA�j���� �&-��_:�����777嶼�����^���o�iI�B�a�y��� �!�G:�`$��_��_�q�C��#s��� ���v#؀[Cj��������?��T�.���,�S2ߵ�6k)\lUZ�����D��BoPVC0q����9�G��#?Ff��� _՚��b��_��ؑ�*�;�&��b�V�a���t��q���>"}q}�-򧼹Gd�F
*��7������ѫ�k���׶v6WT�������7��g���SsMTz�ոyj"<S�%�2����	��^oT���>E3*�XJ3�0��^R�ּ����q헶�FמּW��R!C!�V<����ˮ4^�4t�6�� `g<S���*�^��Rn��D�])\�񼵉��ĭu֓�A�-�QG�nM9�3� �v�yG#F��s�q�ɎGЎ�"e�wP�ӽ�~G��2��d��>�&��"�߾m�����?�$U��1ʹ��麟�VU��᫊tc?y䒲�?�B����86�S�Ӈ�o����ղ��ڪ�j�Ʊ�r^뇹T��~�n�f�U?NF�����A0�B��}5Ĭ�uTB>N�>��S�?(�9w���\X�۴2ݚ�p܇H���Q�\�/�I�D�U=U�u�`�7�x,��G6�^�6����-��y� S.y5��7�ggL��Fm\'�!}<��І��]UDV<<�xU�*�+��������:5���|$s#�UOp�H����ˁ^��#p�n�jr���E��W�_Pif���$�瀛"�A_�j����L?Q�pB���B"���G�����&���7��q�o�S}*|�ӟ��掄�!,���'>�ʆ[�˚/(QD&*߉
zD^�"�䥒��!��K��K)�8Ԑ������������	�?��^sO�����3p+�L�?�j|x�����!ZC����?�h����D�hrט3S3�Y�)j���4Wf��7���8����ͨ=�Ts&,�o��:~<)O��>�ĭp����y���� !<�lj1TU�l�oa �=��W}D2���k�Ў���g����p�ԉp��i����`mOj��$�OK� u®�QiT�q:HAW�C���n���P/\�&�仟�\lX�}���.$ 3�U�v��Rʊ��w8����ZyJ���"$�g�4U���y�u{�}%�S"l6�X���Hky4J�2����O�������X��㰣�|��;���8�qAV���	��"}�>s�w�ڪ��l���֩G}k%`���w�>{�	���y�Q�zҼ2u������m�T%��߫����s��h �Xa�>���Нh��D�s���Ғ�����df���{�R�e4���J���V�����q���\�jm�������ThL4��ǵ�7஍�'ٖ�?���H��d\�!���w�4ń���ޯ�����\g��o��������d��.��Mwck-|���
'N���|w^vF�D6����.)4�Lظ�V�;�n��[��n��7�<�3������g�^��5]6s�_��F=1�ʽ|����ѭ!ɑ���H�p~D�]�f����->���忮����.��(����
�/�1�p���$\���*}����-����8,�z��+_�4�:�O�^��T(Ŀ"������.{ϰa��3w������D�uY|'$�HU��\��� �H`i��He���g����4��6���ӘD���JA�i��*Vz�1湪�ҭe+�nw� _�Z5UzT�z�jw|O�1�v���՛�!��,�H;�o��`�a3{�9��u��E��ڪ8vw�����N��p<��3·�K֐��$O�l_%�ƃc��2��1`�T�Eeu�iH�|sE�J��J�U�.)����*�1{�[^;�,;���H�I���9�2ٵIk�s 2�1
Z������+-'��t����{u �Ϊ���sx4�σ���
��0�-��-��T�8%=��n%U!��6«8� зuIUh-�T;����﫟���94������f����Q��VJmTIU�Ӗ9�N.�X�+5�M��>�h���ʁ�jϣH�6
l�[��Q�I��llG;���bNk��2`��)����3I��6���;�b'o����hԌF���H6�x9�� 氅=n��u:-a���@U*}��0͋D����7&_(.�Φ���vI~��\��`U��шϨN�+YzO&�꿣��|3���{.*�j�E�(�[�Y���:�p}�4<�ΧSoTy�h9�=�m���_�zU�q�4�J\O�9.F��F^E� ƍ	��:m��T}�4b���G��!:轜|,�����BՓңj�X��UN�s���7��Z��q��7o[\k�B�ER��xq-�!�+�E���i�o)F��;ɷ�E&ê�*�����t#���Y�q=�@Rj׍X��ee���=L��-��0#߿���h���<��Fx�ۗ�9�v�%��ZadeB�����
,�J��#� f�B80�����{8�H��#�����q��>S��R�tT%� [񖵟��6n��]������1jw|.�Խ:��ͯ�¸u6��єV�䗃T%�Zv����������> '��=��N�4��{�$��=���'&E}<���@Х�(���� +v��~���W����k��}8 �j�4���c4�a����L����C����|�P�H�*�-�O�7��=
�>�p��RRM~�@�a��Qd�� �ߢ���8�=�<�2�|�Bs�&4���F����Jr�����U�R�������̸����Vd �����q����������G5Z�z�*,����4r|��ੳ�DTMe�D# -.��<��m�.
��4���r��8���&��ߗ.]*K�/N���	�y.�
�G�z��s_Y��^*�/� �%�΁1�#`�ɟA��x��Jx�!�9��|.���='�o��J�z��<��|�(����$ʂPǢ"V��X��LK��B)�/��n��3#��jT:����3>y*��z4t���O`���* 
Oɖkͯ�RUTIUH�V0>����K
Q<*�H�u��z^�*m0�ѣ�6�8}��@��5�_�*J�II��"�FT�Ѵ�S�I%�����0r3.:q0u} �6�|��b��{08���v^;���9|r������9����?
���	ؙ �����[+|��.�(ײ�>�#�ZEDJ��}�k_S�{�<�A���8���Mb{K����+��-������tR��"�$lQ^�?
iz���gn��ˏd,ҧ��ƁRSAGU�l�DM����������~���[�W��^V�Y�I~�q�=���^ݑ�����o޴N!pڶǁ��j,�!O͌�r��-
##�:F�|��I�iE0e�}x�<��M6U8��>�Օ�'�/F����5�v����7\E����P)���)@�7�c���b�y��bpȃI�">��H�����Zh�����.�Z0�
Wv���q�c�����9ޣRΊ�TyԆ��G/�H�5�ѹ/������Á^��(	�7��a�Q�1������yL��`��f~��6��*m�p���D� �w�ٹ����gÅsg���U��i "OL����Z*�C�<4(�N�흭Ͱ%!1����~/yy��3R��XV	w%5��o�U5Rg����ڥ��^M10	���I��^�1{�=���;�2ڊ�&Չ�6���F�)P�էH|/�2����j\�~08h��G����G�q�Q���k8���^����9g*�&R��:�~rt�f=J���ʹ������O��?	/��M�.l��i�g�GO���m?�閺]�0��"� 8{\-D�[��L_I�̼�1vi>9�#�����j\k�H���SR�Th��멜��+S_D���ZS���U4c�E�Nl��y�sNM���0#�Wi��G5=��~�����A�0z�qҷ׃r�xw_���=�dx���(�q(�)rb�d�.4'�=���%P�`�gc���ߟ9���c<(��! (�� vo�G�z���ǨS��������P>����@+�������)���?_ƀ�
��A�7r��H�Z/ߧܶ�~y.�Xa~=|���m��sr���8�8.���{\(~��4�5����@W���S��;9��*���8���|�4�;{�d�� �Cc:��ر�p�������S'�����**�����^5@ᐊ������kw���W��ڪ�dh�/�4}3���(N�(��nR���g
qb�.�o�Xߦ�6ϡcxt��
�ߣ�M;�8~L�"P�������j:�avzF��?�7+tYP��V\�4z߄b��5�ז [1%�@��ܸ�1�̌;���yp�c\tx�5�ߪ#����)2|?���1�[����?l\��?a�q�n������ ����_�;.�Ie%�۰�ਝ�l�Tt(O)bÁ��F$M5@ω�1%sA
lyyE\2O��~�U~��`���1`�R�b���k��h}�Q�5�M�˫���FToX�N��J���I���B�@��z�sP�}C��۝D�r�|M��ȥ�d�e�j�C�ᣎ��M(�Mcu-�ŉ�lT+%0�c,(����^���l�¯~!�w�7�F7��z1�$Jw���S���?Twg"����W��ra��+��f����X��R5>*�r��\�!_���z���4�Û����a%���sN��	��e���Wa_���I<S��X�����כ/����0q���w�i�Jc�?8�v�Ԑ�ν�NB�����D>'�B3H���㿹�j�5�T"�74P��2�c=��44�����;[a?�Z�U��;�z�1�Vn߸V�7Ń���PE���V5U1���Gӈ�{�=+�Jv��2�|�1��Q�-�0�|�)��ª0���p��&HMv�!y��DhR>���J)�Y�N��^�4�TQf���U-r�FU5.=�vK�ͧ�c圮�+��;EhF�^>���U 1.Mvص�8�7?��F�)��|��6��y���~6��o���*%!����S��r�RE��awh� 0)R��hѕ_|�T'
�Ml�P���ME��>��ۍ�7!�胕B�'τ��-��)�����ȕ�=򓷕Wi��G�T���LV��� ��ޕ-oH���*^E�Yk����O|�A�sw��ײ�]���q"5�c�����_����#S�O���B�K�mڬ�!R?
���0m�� �bb�S��jdY���:���	KCG~@��PC�z�ԣ��h	) �8�����z���j�����K����G1<��e��$Z��}�`�k��)�F*Fuv��b��ڿ�=���q�lU�QVث����z�G͍��<J�g�zF_?���by}I,���\m�q@NG}�o;}�d�����q��5-�)眚� ?�@dfN��'O�T�ec�v�v��LO���u�'պ����J�X�g+_��f�|��9���/�S��+oJϢ�m�TXc�����?h�7�|U��ME����,O7ȳE�t;�����0�c�)�<�M�؉��FK�����ĉ$�p&q<��1Ѩ�)���^�x���:�Q����FS</=�vE��e5	�y�V�o�h*��xn��5E�\������i�_��zX��y� iܼ�qw�G����A�ݪ��s�v��-$9�ݸqM*���J�8���KHϸ��ٟ��we_�&8'�Xe!Ju�$�����nQVt�X�vN	 ������d����xQ���;��9���5�T�HL�
d�S+����w�V��}Eq������������P�"���>�I��W+����N�͞�X��$��������p�Σ��_w�%���il�@%��)��W2C�Dda�C�����C��`!@��r�(�;~���sr��	�*��9*��tP~߮�P7�ᠺ�:*�1N��?�N"�Α?G�높S�o��w�ޜc3�����m�}n� ��t��E�����Q��&�=	.-�,#m�����zw�4/��������r��p,�Sq�����<���v7,�/D 7}i��1�&�ʃ���9QWt�^�&�����V�@Lp�#*SGCA�~���D�;���f��;�.E��$-��^;L�̈́O}�g���V�~�j	�	*�Wгf*�w7�,��ɋ���
�� �7φ2}I�-��g��e)����	3j��K�Ka��r���U�\�ډ�W����p�����,��͇��34��d�K� �jH�����pX��a��J�5���5f���Ǐî�;_�;R&lg�oڐ ���C"(nK=����.���w�N�P���wf�O8�p���^��ɮ�Z4��0��p]V�p���p��-�~�����;�E��'9��
H�VN�w�	��!�Ӹ�sk/�ZXιkn,~��v��<��J7�-=�{�yxϻ,;���1���w��M�4���e�+7%�"M{s%�(\��#��L'��+xK�<��W��� �v�+K��;(��$�h���r���z�
�{F#���>{��Q�Q uTd��d���CC��!;�7�֝��瑳a9~E�p�=����T�A�Gt��m�l��0�e���v�����8'��Z4:'�˜?A�d�v㺦�*ǚ��E�!�J���$0�K㖸��j=�B�T^Z��.�m�i�zM̈́��c��J	��AI(]��4*�2M�~1��T�2S�-$�����D���~:z�7��F�.��j��M)���Ʌ��Z�0E�x��"~SV�]X�jPS��6j�k�z1�ϙ���&mI{/LD y!啵u��g�B�7��Jw�lR/> ^�����gG���yϚj>Ze��nvn�/ѝ֞�� �������P�����N`hܚ|;�h47�t�z�gɵ�vwwĉ�ַ�%��¾�U����v��Eq���9s�m/�J��X�a�θ}AQ@�=3c%ݦ۶#���&���)���ҲhF�p| �D�I�԰â��A�oQ�Aմ`��Vx������/=rI@���� llmE�Ӗ.������~R85�I8(7g���C�!}�S��q火�0��<lB�L�$�Q.I�r��8�<�֋6M�lS�~5=�>R�&T���D� J8�t�����uɜ�p�K}�������?_�4��&���˅b���HD�3�s�۴=U�}\�!��1�[Ó�c!��u��<�d�����t��wܜw�9a�������K����;�8�TZ��9F�p�B�\���{}��� D>t/��x�{��x[�Nq�)H���f�������0�f��� �ʙK��ydls�j�j���#�:�\9�fkw?Д{bf^��k���?��&o!��z3��P)|�����Sn_�1�{��nr��4PЊ ��W_�s����f�9�]��x+�_�j�0�^!�IRuMEo�#���/���l�6�n���*���Y�
o\�".��~�g�ҭ��7��/="i�+��JSS��":�fB����M�&���5 S@5�K��u�s#/ ���^�����H�d�������۩�q2�R�9����x�<I�"��A��B�+΅4�b�9�7� t����9�C�WΉJJ�J�����)uŸ5�
[+A��+����pL$�`��oy�:��`��E��B�ِ,BTM9�����ًT�0H�S�͌\ɽ=�i�&�r�`ຒ��S)0�*$��öC*`���������������n��uo'���a1�n�N6B���S��Вz"��Z�$Y7\L>��c�^}�����B���A׎���Lv�*�r|q����(�^�YTz@��Lzx?�MC����!�q������8#u���������~J �~T��4.�e��+I�^������^s�5�#��3��ו{��_�����|)g4o �N��;se��q��Ǎy��q�1�ܚ&����g��mE$v�7Cg�
���g��t��I��oA:�^��LS���Ƅ�^�Ѐ��V���[a}�f�"��������n8�������я|D���o��x_�����N@`�YU�I�
ff�lF��gƭj�#��@��h�n<�F ��{3ǎ�������@+����q]��357m׍z�~������΅!]\� e�jX��l��j���~TE�n�4��ݏ=�2��[�����φ��v��~ѣ�>ff�Ub+�!~��]�=��0*خ�(.itRP���Cs�_����Q)��u�i�?��H��sۺ�H�;9�h�P�@a�Y�D�n�Һ�g���T��c^.��c�)a�v��� ���{Y�6�_$
��f�����'?�)ͻ����)SO�e�.^P3Hi�aH�"/��0r8v<��$��x���O�gjB�Q#�tڭp��uUKvz������R��B>vi���s�=W�e���N����`P��h�
"6|�z�6Y�\�ٺ��F������ѹ�G�A�h��jԭ2�
N4?ͻ��mFp�<������N�������}NJ�ttFY��26^r�?��5�$�`=�,J󱧞@"�����ͱ�d��}l�EirS�L�ύ�{|�9�3z���oIߍޗ<���#צ����i�X[h��C=�	ێF�r��W5LNN��|�Cѓ*��s�KT�I_ƞyG��{��2DшL�y�����+<vl.�o�G���̃.T?8917���y�9�^����"F;[aP1
�y�~=�ў@Ƞ�y�U�`����H����������Q�!��	����x֭�V�Y�l�&�U��wOQXz1�x�7�W�>�0�6��6�nj.򭰳��j�����O����*�d|�j`��2p��*Uk�g&5��V&5��hF�3� ad�j86��YSU�3�Ϋ�M�Ս�`R����q�ǿ�9���N�T��|H�-~�d��C��_��
�J���]�G���Դ~�����n���9�����UZ�]������Da����8 ؓ'�|R���򈏐��KAB��t�C5�e�֢
8��/^�W�LL�=�}�ƍEEH�
�&F��.�{�p��r *�3��DX�y\{N4����O@�~1��L��֯˭�(�\_]S:
YkQ6��+ɅY	�yR���L|/G�.��H0�v6g���crQ*��eɾp<o�ê�7� ��]p(W��E�/?�-n�j�mS,��+V���'��"��~�8 ��)ӥ��=K-��7����?�y�as�[��ߒK�{��8�1�n,z�ҥ2/��μ�|,�)�$ߣ��ǝ�^��֍z�3ӓ��YJ �#�Y7��D�[��U?��s`nH���tWr��#�?��,��L��H]��z���eՔ,�[:���R�ťE]��U�9{:��3^8qBDX��%|��VQ��)k+uоk�Ѕ{B��IGs�;E�B������p��7O��J����`5�K/�n�\�`��H�``뎴Q��]/t��g;5�zqЄ��j%y���V�sX�
3�W��3����ă���"�U��*�W���I�;�LRq��=�_����ܵ�@A��ޕ�	H�����5ͭ�J-2a{��T�y3W�AT������RZ~��J'��n��JY$��W^{���Az��_[�kG��wr�qǸ��8��N��w2Fw�.�){�o{�����ffg���x�O������<k�q�^���Y���:z���I�w�a�� q���E�J�ɿz������ H��w;�Į�o��i[�۩��Pv����r�Vi,
�ihY	��4J|���'-)k0�S�#G,ޱ���S�OR�������}/��*1��]�h0�R����%�".	��RD�I�J��������� GMtp$�em%�\u�V��	Kyٹ=�*�~�LJ�h�ukX���՞n��΍ab;�ƽu%�pp��W@�ww��q f�Ӓ���������;��}������0�5�t����>,�?�Uo�l��͍2��H ��η��[A؝"B�1���F����q��wS�r���Fpks+L�
�� b���>��(ޖ���{�̹Pt{J׬�9q��ZQ7��ݝ�E
��-Q�h��Z��as��r�1��M�[���F����ꠧ�5*��7�#bUVUB��Kc݋���6�}�H �9������!��סJ��������aeuS�U�7����R�<�d�c���3A�,^gC�!��j����
�8.S�L΄��v�V�٣Cr7��/++�D���k�g^����z"A���z�;�d�Y����b���݌B7�p��.@��q��O�׽oVw���Yo�E �(�Wt� yI��7��g�UzdH�L艔hD�FA:x������xӮ^~�'OUvcvJwW*p�c����2O~�9��=�c~\�GV���SW�'�?r�c��$b���¤��w���ҭ�p�Q7o��c�,8�Pf�f:�s6k�����Um4��''P@��=��s�k\B��;S��ǟk�	�g@�h�:Ч���]�4���gۿ\�9	��j}�T�愨���hw:�J���2��FJ�7��l݇k~\P3L���'�l���x�n��̒ �������k�Afж��C��<#60&&��{��sZ���r�V� Mr�<l�.
S��bJ=��m�D ��F��a�ȩ�����}ap��������bl���1�Q�,3�����ټ��,9z!]��?��Nݰ6�s��^	�lv�k�-S�.,xxM�=�\���~�ԝa��}a��}U�K��n��f�+�ki��7�Dk�2{a�R_�=jQA+�nWdX4f �������h8{~%���*������b8~�t�� g|:Ω�F�޲5�<u:���V�V���Zس{Wع}���!
D���XK�ֵ�N��W�N�ݻv(�5�޼����\��޻�R	,�y[q��1����~�5��7\�"���,�/�K�����HS��A{�ݻ���)�,�j��=6�ft�����D���4"���/�)�4>1)>������p�ةp��j��џ��:'cab˶���/�����r��^��~�'�0�}�;�9=���zVDl���(f����B,�im���T#�ݕ ��|�A\�R��Jkn��ȏ˥��t�:�R��?�P�s��{�g����}4���@���u*��~�O}��T���c���=��lwj�9�l }�������V����y8U������ysn�ߗ洜�Fe�<��K��ܙ�#EE��N\��ײU��-2�k�(2cEd'�H�����Z�2�kV�q�1�U'
��7O�tk:���p\��ə��@�����ޏ:"���i��Ɓ�M��<M����&��� !x�d�t/{��*����+��L0��� ��u�����u��2yD �d�ܽ?CȒ�Nm��ēH� @��1�'q�#� ������:r��!t����͎�WP��ʡ��o�����}?�cWO<�ŋ�d,�Z���O�+���@���
w�ٱ�&�Yu��s`y���\!�2?k��{{.�E�`��G���u^�yǣ�;�|j�1'� �b��&�'�jBO�М"��7|��!��"ѹqZ�cTR���c_$j+W���~�� �UW /��lK��p9o�׫�)��[�yY�LE�X\O �ݻwF��G��T]qN���Ⱥ�����lH����1��鬫 �p(�e��0�#��|α'�a���g1�>�ҍ�:~�Ǖj���^~�p��Ïh>�������]�q�'O��cSZ��/F�=v���"m<ç�~JQ��>/��"3��ٴ�/z�\��l��:|�f��X�C��/~Q�#�@������ǆx� �o|�ᡇ�y8����l6Cjy�^D�y?J������z��̳�h�v{�������c��/��~	����o�Nѩlb>�F_^*�å��s��щ09>�W{��KIȒ{�>�T�X������E��
j��ƍ��W����r���$�5��0�?(ߐy�{�P�5�Ô�k��H��un��F�Vj���F^����F�x��nݻ���dH�e"���U��=s�pn�ԴZv��>�T�#IT���G�8F�y�T�fσk�Z|!x�	�&��:[�&��΢pjb�K^�2F5̫�<T�c�w��=P�W�G���ҳmd����Iq/g,m����a`7^�q!���J�;@&�J%%��J���ϗX���_���I�̲��ď��ʍ)��A�<�@~��������c��=' �l5�ˇ^�xg
C�<���~!q�^��m!���8��=��D���8���h���Q\d���ީ�Óaqi=\������Q~�N�z+T��F���m��
S[�#؟�Mv�m��܉&n$.#����\��E[Ev�?Ls4LL��V�����ņ�f�j��=����kaqu=>׍�dmw���w%����p���U�jt���y��O� 8@-��K��n�0��amc]�xa|�5��&��뉺---���(b�Q~O)n�q����^�LD��z��+��?s�˽�7�͢���h�p�zߔ������͢=�EPݎ:���p��?��?O<�D��;|]�0�mpT\����^�����ǣ����Ri�� � u�#�F�6?�Q��e����Ƽ�w�N�l��xy9���7��Z �Y��^�?���Y�9�#��h*�)d��쑱qU=Zy��Eb��a?�G�._k����j�[�J��� ��H�,>����g�d6*��S����O?��Yun�	�
�)��qR�o�G)|��zC�T���F�$HOP��	��e����-�N&�x/��t�E]lA|�ܫ����H��_�Mpo'���c����"׿���MIe�^$\+�(�[i��[⦅46U(l�Eh�x�E ��>^���Z87����4�q �ߗxZ��W�e�>�'�E⒦���;	�� �b�*��79<h�6�� �I�9K/���R�?�����S{����s��4.L��ɹ���H�����F��-�]�
ے��ܣ�F�{)R�.z�B"������ �u�ʏ>*��Lˁ\���_Z��nm^癝���k�� (~�"7I�)� �ol�M��8�ӛŨUI��9��Q��c� ϗ1`�g�m��v4���B� -��{K���u�d��l���h���%#H�H�<�5��¥Eu#��i����שi��ؘ�8@mE:��}�йf"A��k�f滭�2)�����;K��*A7����Ű�4����Y��?s���l���eN����98��h������>à���������s'��|�������j��5��5�ln\�W.��k�F'��Ћ )	��fu,ְ���۷WU�>��7'��㥢��[�Y��o>�H��� @���2d�F2!�C^k ��t�"/|n钼/���(ke|̚�*��fSՓ8D�.�Y�(�yWNe❖��s�zmQ�U$
��pN�A���?�#G�������	�77&�}YW4yo�`0%-
�����r�9���Oe���A��V��'��R<]k�etL�@�l�\;�5�����%m<dOnҁN���+\��A���ah�o��x��"r��X�\ܻl�^��LOE����ڱc[\L�l��E�R�D=��[���r�,�J�'����'�ͷުRe���;�PK;�u�h�3��w@����!�MS�V&|�Jc���y��������o����9`<�T=O*Кug����Oy墪`�=�ϟ?�0�{��V��ZU%Tu��U��W��N"E�1F% ~�MBI%�͢V��ԑ����<��ŋ�.��N|FK ��ߏ���E��x)hRp. �M����� ������4)QTy�{�JW�@rv���	zT��W�� �i�*��I?�׉���j_6��U����H���p� ��HPv�8$A���׵(۳�����*����u�����k%�]����+�)�'ƝaHdO��т�#49���ıY$�J '��n�r'2�f���oy��v����#�3��Np�^��??������������/���A���[w<���M$�+:����1���������~^܁���q����f┑`C V��h��co]՚T�;|�tT�9�~�p2:q^�r�`�y��_��C����N�dC�pC���MN_s}c}5�	�Zs�S|��z?	�F�v�D��F�檷Ip`����!f�-d^��= ��\�<����Fҿ�l�9�)��͈�ξ�SYÌ�CϤ��H�I'�n1�]$QK��j��7�T����Bs���$"��_E���y6��r-�~�gX�l��,�V���`���f�	�O~���I��=N��X�_��QUv�*��D61�*T���L��F>C�۰E����-|�H����`���O����h�G�0$x�<��V�+o$ S��m�Z��{s��`d�0�����v��)'�"���r�u�MEH ==#Hy��J �ԥ�P$��j��^��o���NҺ�4&�к�[߾V���L!�)7���$���%�Y����0:��<�f��m�ƛ��ۨ�z	�s��9^|��p��%qf�'��1�I7�i��-��25-0�h���`�_��ܲ��[��f�L�"����RF�R���][�p4$�趡ѻ��Aͪ�ģ��KWDfpF���ʑ�O6gd�T�*� s��[�������/�F��uV��B_ck��q�<t��M_��y�!_�����)��x�u���>�Vox�j���������&���� G �<�"�>~àЏ�婬�����1)�����	��ԧ¶ċ�s��p�Ĕ�s�``����_�����ijN�`Np�&r~�I/�Y
�	{ f"U�xӍRǦ��R�ӄ��g΄�q�q��8AJ���!�����F�NtZv^�Btr��}ц���1���*�o��J���Du��Շ*���#Ű5���q�AGs�h�/~���p0$I��F����g*�(��\��77;�ji�H�6IPr��ʾ5���a&><&�w_%@�}r���4h�%u���T#Z$aū/TP=F�QP�5��
���|��<�.��b[{����&i�͙��Ώͪ�+|�����Ԟ��s]ј/��.��(�9,įcǎ*b���Y��Ty۸`7�a,����M���ؾC���K�ҳ���/�Yp��#A<�;v�^��BU�u�z��j��#�FĀȇ<p�i��a�ͳ'���Q��
3S[���u`�yi�y���pm��w����N
U5S�ڢ�ϭ��)K�sp��^���qn��L��/m���ݹ�vn��m��>�4��N�zK����o�u�ց�h��?x�@x���P�o���0	w*�H-,�D =�f��Ќ��l6F5V�WU
M��Q�+��]��uJ-�h��!% ��پuF�#��Jҋ�u��̅T���k��D2"s�D���$��m��}�*��+-��Z"%�$�p�~���D���m��i/E�B(�z����2x9;F�r|�|��u�Y�f8r�9�����瞜G��x�xFk���)��M,S�Xj����Zv���
�w¬��i��]a���Q��#2̼ ��\@6!W6�������ұ+���~���c����r�=������rffkp��<��;,#I+,��z���9ԡpf6��I�}�?��b��~�hkY?��88 ������>����w߭H�ѣG䜰w����D}L��X068����*B@�&9����9u-���f�o�k��n
?��%G��')�[��
��0�56��(�=�~�F+\kR�5��]T�O�ް{�l��7�P٤�l�ȑ#j� "S���`=r��6�p���S�O,��"��&���S��_���O|"슛苇^Ry��졑Pv�i�
m�����z�F�2���'�����U�A���fMh��Y4�l��#� |�D4�>�f���p�S�Ϲ���y�9���@p��X����;�j-����"e�Ja�w�lj#b� \�E��`<,bOK�/e�#�x����`:H��O~�j4D�$���6,�{�+$������d�er"����­q��lۮ��¼R*���/.Q�#�>�cE�X������|������/���`��^B�G�qy��±��e��W����!�&�H"��0L����h�&uR鳖�`��RU���)��<^[�6##�����@`|t2�>S���D�8)<�����aum���|`G���"����V�|@(�4/Ec+E�x���� �[�7��4�߹OE�R�H�%��qH�q^Єrb|ʸ*qX��0>^)q�f�0�iY������yD���}�:Iѐ"�JT��h�|��Jֶ�T���{�x:��I�)=���a�H�6���i�a��IO���g/OƖ��=����+������6=�U`��x�f.�����DP1�qB���{a�B�ɏ�TkHQ"`��?�TMC�")j����LD�A���5�fg/���J��(���V���W�����_iA �S|=���������vj+����{��c<$���k�Q�ַ�UɊ��3p쬵v������Ma|��,��變֭*�5�eJ{ )��^���̵��;�+�ó&��u�����Ǫ	_��E� F ��dK�r�p�pZX�ʲ�Z��H`�/��SV�L��L9�+�Y���U/\��Dj8<b�yB/a�(���T3E2�`[��e|�`���{���������������aRVg����a�=;���Q�v`���ϩh���ȫ�Y�Rbh��[i�����B�qQ./��ɍb�B� O���D
M�b�
�� �\���<8(!u|��sn�^�:
�5�� �C���C��o'�4{�gt�m��n�^��|�&]7��/��*tVV��j����pF�h
�aSm%�N�-+?�5� .����(P�tמp�M7s��<N�<���hcP�j�%��@�"�x�|�=w�����F/e�̴ �qM�S.-�7ܨ�D�Gz�O���`��_�ժ����2�@�@
}���]�dlS�;�VRN:X���6��+�j�[��4�ϩ�Jz���.�_gΟ[�Ϥt�	c5�am?��Ј�j�*���@ $j���؈x7��8��+��=�Ƙ�L�r�Z����
Ѯɩ�@��dm�N�k����j�4��*r��MkA��k�ָNg�h.Р�9A/�'��bDcgJ�e<OW@��x��cee]�*"t�O�̀Y:U��*�V(t�k� KG��(<�٫^kϪ�l4�5/�I� 1f����x�f�3�\	��9��'�x@���)�a��S.l��ۿ-��~"?{����ת�0��Y��[��{"&�ԇ�[�<��O<���2��a[w���v�[�;�~��:C̦N$ù� �+���3�m��Lvf,i��h-S��9��X�@Ý��A����IѸ�9����4|�[�WŁ��NI��ǿ�Y��hc��'M	����-I��UZbkp���6k��{+�0�Ƽ�������sN��N���.���I�?���g�;�6����4�"�U0���@λ���z�lm����	�i��Ÿ����5L�&�me���E�w������>�[Dj�,�)�Iaۢ"��&�$X.��B�����pzԁ	LO�^*�!�)����?,O�4�4)*"5���S<6��P�GTK)��rL�o�c��81�$FMR]`q3�?ayQ� !�����č�������xti�<Y~���]~kX�ӵ�y�>P8�0�J����l���\�Q͏���	x2��_�47`lL����m��v�����4��G�h���B�o<�J�'nҼ�òÕ D��pFǭW���AZ6
�-#�v��2�ϸt�>��|�"\z�<p�/�?��7=O-xw�>�����w�������[�%9t? ����Ak|������<�p^�b�"�Â����o4�p���	�Q��\�q�8i#T]u��f��v�3OaDC�x���H����4Up�;#��+N�ǥ�FX��w�h�:Z	��7!���/��\�~�"v/��⥍���Ƙ��y�	N�MK�rs �o��� Tv���}��Rq$޸��cEU����ǁAi��!smd�*�.W@�(���hVZ<��Q��ҟC%���M�f��_7N6��:�\�A������Jh�5�Y3h�KRf��t�s�r�	�	"��)6����Н���p~�n�2]����w����kw���sr�������hq�x��uU����}��.��6g�Cj��s^Ae)=�xS�T�	HNMm��6s�5@��*��0s��V۲|�{�(��v'���2��;/��OU�};��7�{��j�di��]&��*��:�{��:k�L��t:��-��,@��=xX� �����ܹ#eD��\�����Z�g��m��C9�pV��?e��kr�'��u/�LDI�8HQ4ƥ_w�Z1X��&���U=��	�B����`i�fI�^A(�Qo�=��h�9/�E���&��\q�IC��%˝���T����7&���K/��Tm@�̊ �����t��<.���ܳgoص{��D�������f��O}Z��{E�sz�� �f2��g?+���T&ӄ��� ���|Lsc6�����V�������g�բ� �x�MB���!��Y�u���KU)�y��q�<�����}G�TY����DZ���~��F9;;��qjjZϘ]d��Z�lb?�ᏢG���{$e��54�4':{ 7�@����>����?�3���'�+�����rR���"D�L�<�0�����?���w�+ :919��R/��瓓/�_�B��~*�
Wф�H�������@t
L���R��`�� $S�V�I^S��"J�J��ڪ^�uz2썀6�3R�6@�MQ���L��	�R/.-�ss��F˚�Q`=��T���l2�Yc:[U"
i��:�u��̱ ���5���tM�K�[����ZK95�D��8gqm��n�N�¥ѻ� ����"V�<,����N��y�����D���Ϡ*9�0ٵZ��jr~�p�)W=�S�{B>�n&g!�
��U��2.��$y���|>�x�Ǐ�rQT��C����^xb��6��D<i �9x�4��簯:��Cc����˧�9p0�2^`��i����OF��t�ɏ����ِ�N�H��!������0��:@R�e(��ϣׯ�k� c�!j�Q�_9aZ��ˊZ��6�8,�}�_����Ea� �җA�G�(���>�裏����< P��`�w짲��m�5M�۵�{��İ�4�%:Jˆ���j�]��JQ�s#:4�^����p�ʖm߾C���K�q��R��~*e�W�|-�5�$���K�����$T�2z�>6(� �!O@�O0WTd���x���EuL)�˻��qܐ�I����PX\�p�\x*��~�o���y_m��<`s��@W!o�����0�^)�����w�;|�㟰�n��ީ��4�L���k�/�`A��}��_��,��>_'�sm�=E�Ӯ&>��B��\�.ݮ=F�v��Q�L?��F��f��'�F�}�<��c�eC�@����Cjѻ����&��̧�3v �#n�x'������T���i��?�a%Z�u�(o�S�:�5�B����h�>��D1\;�Bz^ s��I�������8��)��ܣvP� ��4S�0�_�tF)�N4�Ȣ�����wv�|�]ی&Q����c��ha|��}��n��x�z��ȸz+!Z7{qA��5=3SD�p�� T�Y{�'�W,���i��#V�mZ𗤿1!����:��e2z�����So�2n�xJq��x�0�,4(9g���n���h�υO��(K���f�fg�W�^L����;�ڬ�<�ɷ	�yPoܪ���5 ��׈R����Z�5�8�>�^��)���cOv&�(6Q��TL��(�e�c;����o|��D}��f���sϽᮻ�
�V���¡�_?�R��qpf`���c�Ս9��V;�g�̝w�������^ #�0�uZ���v|fq:̵炋�r /�p�S���*)��[��ZJ����7�{�?��5m�������1����c)�WM�<�^h�����Ǔ�%�fq��qg��|�W�p��6��_����f�
k�cs~���j=$�#��'�	��h)����l��&_�(��(�<�	��K�}B�01pA�'�'��GN�j�RK��p��0h ��Ԡ�7<����76/Ε��qB,�p����*���X�ꄝ����m�ɉq9{��@���|������C�T�1"�+��� �����7��1���M���^|��r�����&*�ӄ%��&͸A:sq;�5��k��>����b�x�V!RT�ȹv���	T�������x.,��c�G㈔�0:�u��(���1-�Z��m�L�kh5jr.���������97�%�#��Q�s1�|�v������s�&�\����������Pj��������4WEb=5X��pO�t��rm���MӨA�!Uyy�vM������Rzi�����	�{��.h�0%�#P�N��e\l����[�������S����/�>�-��V��"�䆛��\0�	�.�`QM3�c�}��:�J��R[��_�(�}#%K��*&���	B$�tSC�8T{v�Pڃ��%�6B�X���O��C�K�&� �lxBDpٜ�Fv��nܫW����T�f��C_O>^8fD��������"���^;sQ��SJ	O�#������s1<��q�}�i�c�r$�J��ܹ�rl���'@��3z�ү�-E<��3�³�<g_ii7��^J��R=���]-\2<��K�[K�+�I�%�`d�)E
؈�wٱs%�_\pP�J�oW���5��I~�ߌC�!k$�����ý}_�y�D���U;��^�c�y����g�$����b`� ��̱��}^>��ƚ��\�w���^J�?1�;��]���|�b���A�R�F��禨M"�s=���YEDo!�$q���'ȧ�'\�㪃��PVި�h=;�5dH�(�^���Cu�P$�{�l|O�Sr�	� �xXlN���ŋa5>d8)�p��6��н��#2�Y����"|��ӧ��>��\�x�|�gA �җ��F�D��=��`���O���
�s/�8Bo{�[��aPn������������̼11_�|��BFř{f�`T�hV�^'���7y �64e/����p��k��kzn��\��{`y�@9@�V��x�BTF�-z��������;�(�1ϐ��JγP3��|Pa}�x|�7���C��,�ޘ����R������
����ڍ#�{D|$M���U����6m�0>^��Th���`��Dpo�!�
+3�؀�����\ߺ%ΕN�X'��%��-��'�v*uƃ�4N�"�M�"�D��%�N�~+7:Vc髛 �{�^���1 ��KiJ�\��mM�D��Q8l�x��P��4��c$���vR|��!�k�[53=�㭒p0��K���J�p��{�j4�����T�ӗ�}�u���Ep�O��Rj�exF�"����z��fN�fUI���*'&Ba�QEU�����r�pzc�6����'?>�L������s�#�\�����Z'� 9N���J�H�V����t��#k[��/��c3��j��f�6H*����uA�mt�e�R�=?#e0����T��=��kΰacSx�ݲ�D���J�\5y��֯"[n9��� >�s�ܹ�9�io$I��炱>W����%������"kF������;�%v�t�@�Q�����}R�=�e��D���G{�����������U�+4���*��=j�m���i�2��F\�4�$2���x&���S�L��q�@M!�Ա�(EU
�"�uMQw������I��[NxF$'�Bn���#�L��Z��Ҫ|��.��UK��7'����0���BrIv�L��fj��ws��� ��N
�|�׿����|YBF|>��/&/�F#�hH _�� Lpq\�OĻ8��˽<���#��}6��Ɔ���ឡ�Y�Ks������:'�tW���cNd��3f�#�<"��f7��-�߮�cQ�x�W�0?�"e��萵������aQw:[�
�Ŀm�z\�@wJ���F���8z�&o�0L��G�
��!
���ʄ;�3rc�Oyu�m`�A#��s}Kx���3挍������W_�|�4��
�];v�[�\AŴ����v ����k�ј����W�=�Ȣ?�69�߬?��d��	���¶5��tX!�_9"q�W��Ҫ@&��Lֽq��∾�-JѪ�/�)��7��������L7)��/i#�o���i2"�ީ{i!z��Oj� @�q�6��oS��cǎG@�vn�*9{R�c��[ٌ��:�6y�S�����thi%���������D<��,��?���ymn�y�y����+�@�9�;�0���:U��/���������O��+��Һ+'+��R�`1o����zÑ�5�j�h����ى�T�O;��ɱM�[�H�4r�o�l�l��TE��Qb?��	8�M& ��U�>����㓕��Q����z�$ʹ~~�/�}J�/�h_�����7,�{ƮqO���PjJ�� �=�>`������5���V�(����<5��#�k/d.p�C���a~P�f�E��87Д�G.�n��J�TFՐ
r�+S�ع��3�K���yR]�/X�AO�X�\�fQ���h,8����O�['�����������@v�]^cR�}��5���Q
�Q->O��v��t��Yy�^J� �	Ǘo���Á�sl�����9������SW�Ai�c����i<'�&KO�t�r�Gn���_�EU�v��W��&t�+	�&h��,9!9��;L~�<�n֌�?�C�#��z���7дH͸�$�C�U!FRc�Iz��IEX���z��^�r�*nFF*�@�
#D��;��N!�����N'�%`"���� `3۳gWضc&z�+��K]�����T����]��t[$�X�5G�i�#9�¹]��F?���~��E��=vyC(�c$s��������)�aC�4ޓSauyQ UϽ{v+Z���#�%��w�mǶp>�}tw������k�K"�ѳct�Z�7�[K^" ���M�I{�qR����&`�q�E[�P��JISR�u����� ��	��	q�1�R}S2@�:>���l6��:���� �N�S�5|��t�����[��3 nNPD����W5Ik�9}<����Rg���w�����Qg�n�)�;{^i<�dX�4Z�⽌�
˔W3/�[�A0�}?�*�J��40�7-�@�u��z^��5��eޠ������I��<�6s<: 3�3U+��q�J�5�� ���6�%q��䱯.�&o1�xY�8۸ ��+0��!��=2/�pO��CFA���3�;*��^J!-�E��1�VqԭH��) ���  C]םX�܌����'���Dh �D��3�]�ϭ��g�^�������}��_��m�s"���d\ҾH��;�fC�$��QQ9�G��B�&�3���ĉ��^�L��8[_�(���;�����l�O��sǖh��5���F�!P���&�虏�� ��
�*n�=�qL./-g����&���!��d&���&��2hl&xB|=�kx�DGL�nX�7�ph�|f�;����j���FB�Fxh,@,Kp邱����!�^�(�I(�#9���W8h0��0�V�=y�dn�����赑m�Y������p��G{x��9?~����`o�nyly3�~�쯓"k�����I�F��CDJ"<!�F����yi�(X)�En��������ؖ:-�F��]�#ǎȀ�߻W
��V)�6�^�2�x#z�7�-�ah��w���q�̍?��?����hL�>΁gh�o!w7B�"s��?���ɣTXل E&�C(��$Q��ܩ�J?1Y�#z�k�NE���+B c|�+���#���!C"2�9�Ҥr�^���#B��2���мA�`��p��4uf���[c�qvS���B���N;�ڬ�:��(��q�]x;�,}
�ׅEذ�C�ʨ]C!}5%���eݣ�kϼF��j+@���|��]�#��`����;�qWx��W©S'�f{S��l$�����޳/�ܽ��[� 0�����	�Y0*�t��^_3�2��9`bM��G���zH�kw�pP�e��eIJK�IB.��=&@�Z6.� �9K�k��b��Ɓ�I����u��m�/&�g^�������I�=f� �	`b>���?���P�u�W�W�/��:�����"�������*�h��Z�ubܴfЉr��*4o��+��:"l_���������w��yϧ�L<�#�LmQ�d��c|�� A����uD��k��a�Id��=vJkF��q���#�O�t��w�]N`ejj\����f|���/F�\I_������$���m5��?y4l�մ�p+"�A�b����G �u�{5#9�E�9w�ZW�Ԥ�������,��~��%7�w��/L҅�%=X+?MBE5;{�e;�D�rC�d��!_����º�����v���R��,�K`^��&Fƥ&L��~Y`O�8)�^?YU1x��zЅ�z��{�ʯՏ��+��U��uD�� �e�77�	�P�3��qfl�l:YK3dF�c�zȈhc�j=č!�\�bc���gr?T�(ebbZHReM����FJ[mQ��_�c�-��-�P�>u*��Cߌ���0z���>�%�����Z*��c�=e!���qR�s��Q����F���|wP
ঌ��D��	�.Iϡ�ׅ�S�Tڥ���ͪ�w|�T)0v�خ2i*�֣A�L���4���;j0�7%p���:F��Jj�P�(M7C���P)��7�&ӻW8x����<�ezk��߭���#���TʣUtR�n)e�e+�+Y&b��e����``˲�ЂJY���)�~��j�(-�����y��ih��Y=�M��0�Ui�M- z�`�/
~|����#ŷ5�N�16��o�w��z��YW�f>�u�;4�I������p���|�9K����`�����N �%u��Oa�/�*��_�x��i�*u;"0��f;��3׸� s �eNd���<�%�ȍ�$�{��:������B=����������n����*�*�zgC'*�$b7�J�,6�0��^��;w�c-���s:��ԓ�a�D�>�v�sm�����G�i����ga
�+��۫��Ir%���uL/AA��FH�B���(��S�_�x�<�帾&��:�~w$�(����c��ٹ��	�D[�VR�__��tZG#��蘘*���~�S�oO�;p�^�b��>s����e�WA�ͯ�QR��	�&���v���5{� Sr4�x�5M��͗��oa���Y�f)�D�c�i �T��!'�9��Gĩ�qP|��c#�d.$PdQ�$T��e��El�{�e�g8�#��B�Fniy�J/y�C���(M�F����=?g�+B��TFl8ܝ�`H 4�ݴ�rT}[Id�b��uI���Ȯ"��!��"��_~@�'B�6t>�'�8��]�S4Jm�̤(l�����t�+�CcIqe5,Do�\JME�Rj,��D����W�J�����l�w��g�[@��yC�Ϛ5�c�i%����H;bhy.t���7��;P�3�h��f�{�s�C8}[��T�ͼk�4�*Ӝ���\s�a
�  @�S��`Z��QX��4ef��R)D/m��+%�HM�����+U �xR~Kꤾ�uJ�]�~8s=�z���p5�#"��X�]w���J3�y�t@â3����z�t�Ф�n
\��o����x\7���I0�-����7�|&�H�ϥK��ZoJ�ʦ��"�3yҼv#UK���y�	lv�L$��2�{)��@����M<��F8q;S�����S֍6�5�rBc��'�7�����	AN�9�"�A�t0���[�9���W�Ϯ��X\XT����,bkK�TT"sDF���>�w1��'	ܗ�����*>�'@���q�/i~r��8 �N�g�0���N�ތ?���c�Y��-�,1�X��%#"��tQ��=���l��@�=y�t��y�+UK%��b���D��s�T�w����*;�~����zrBǪ�/�"�B��#��/,//�3��LM�q�PQhَ�z�Q1������9f+M7�3?����{�U.��h�|m����]��UI&�4Q�]\�������>�����Ŕ�]Ä<9��'l&�!�=ِ��	��7���j��	P*/�<q)�2�.�J��JX�1�>@L~6Z�� ���H���o^J��2j�����2$\evޛ�M�ӟ��^�{�C)���`q౐V��!m(\�{ �A�H���{��Yd���'���~�
C�������Ȼp��W�q�J����3��y��E^	�ʩ�y�O�N���7�~i}E�M �4��j\�}��`ˣ�P>��cJ3��➨�8wv6�����V；�uE��SC|�9�Rz�bO�a$��ސ83�~!h½�yr�E<�Ѣ��B��s�>�;�?����[�Z������ݒ/ǰ��9|`�6���Ң��FCq��u��AYe?oQ�df�θ�Ӭ��(�6�������RB�^�S�3i������Z$r�F�MA�ome] ��7U!EǺ<�հ���@����j���5A{U���z-͙�v�{ �#	�Y�5�0�z����RO"7)m�\�&��D<%�����n��~<�mG���a��T�ʜ �b�������_�D'�����8.ű^������ ��~ҡC/�% �����~��^�>�7].�ɚ�
2��tӦ\��0�8o�#�K�@�G�G4�O½"ɼ�OX��\��nMzBւ��1� UA&��)S�S\�#�s	 D�֎��A ��n(ZV�y���	������Q�\�РeD%h�LNʔ��eJ�z��ʢ�㥥y��P��M�
;�W��Q��L�A!��o��7V�7f��p���8/6�d�eZ��=@a���l- (F�N?��N���d�w���9�~�fU��F�h)6���X��hf"h<A�j��@|T4�>����1��(*Zhj޲(������٥���?J���q�6MLZU����\���HN~M�Ʉ���qM85�2}��$7G->g%�x ����k�����$�N&��X���T^j�yb�L�T]a�3M�a�(��!PEET��x��=��io��HyȶJ7&�E�L��7zH�x�Amr{�����'�9l�.��Ba#>'�QՔs� E�FOA�u�� u"C���#/�8�Bn�aȩ�)r""`�c�*�Mv*zgS"ZzGgB������gōarb���<�ȏ��?���y�F���y�H�O���T؍j~�b�
.ű�@X���왳�����ԓ���`سw�<�m�ħ_���jL�i_+��MS�'�/��/j�W�'���}�_�{�{"ùQ�������O~�&�A ��� K"�$ ·�|����z����ϫR����?zL�G�2�ܹK%2x1g�la�4n�_��N�>A�6}���ML�@.�̋+�QW�bd,��I������*�4Z��u4R�L3�Pэ�2e����J|&dl1�2|����K.� �'2��8�5S���Ƞ�Z�顢& ;b2Eg"'�
�����)m��Z��xNc���Sq�a<L�l(����ԩӡy�J���W�F����p"Οs�d'�D�m��Ckt2��@�IF�b"q�n}���SJ/!��[��Gx�4O�u:�o8r@� �AL+�:��.a��a8y}q��z��;_��u �! �����R<|��=�����_��}�s��<����9;���Y�2��셹p!�
*!'��G�'�z�
ꖞUQ9�C<�$��KUM��k�-���j 48;5�*zQ==oS�_��m��j�m�`�.�+��{�+�n8y™	�.~}*�md.d�MLLT?s~�ÅK+K��9�O}:�S��Ot��	E�=���ۮtq����FE��Npn_?E�s~Z��~��u7U'1��uL���u磽ZU��kwJ�FZ�Mkk�����HK�w�C8q�XX���h7 �c�Xx��w��XG��v�o�x%�$BX/3@�^NrdBa��k�WsM@���=?��j����
=0�^�l�����&�I��(���zFbg2���ƹ����j���`Z�kz.z��<�C��5����Tc)"DSe����%c��k��O*M^)��R��u4IS����Ĺȝ5�+�l�o��oDT�*i��!g� �Z�/��\��_�?nl ��ƽE���9�l����8	xd��Ȱx�:o�4A�fj���Eබ"ύp* ������ˢ` %�DY9���P��܁CB�a"^�E�^y吼���qf���8��Μ���M�"��zΏq.�8{S��vY����ɨ�R5�}�6��+�Υ0]���b+�G쯗������er*<�ԓ�=ςK��zX�+��xyfχn{C�gT:�޵K�zŠ5`X:����c�x!����[L�������t�Qr�KcYx&��fϦD�:Ik��	aCk�g�F��Q+�:��<u5��tX+�k��]��"��������M�uY,.�o��+������!��{�h�����g�׽Ѓh��q�w����I�?�ؓ�;F��Iz:�i'�d��=�l���O�E@ ����o��j�E5N�D�f��+�>"��܏|M{�#���v{K�����7�k���4������
�R/�X�D7 $�s��"i�řEE '��L�h���:H�k�oT�u�x�X�L�|��߯� ���E,횚j�Bp|b4������;�hn���� >����3��^E��#9�IR��1/��p��v��c�����ڪ{������g�}��3�ߧ倣��	��Ȩ��]e��L��u��yX�듗����H�FP&����6X���
�σ�����	�Ǣ�}+�W�i��_��+��f�O�Rx����ʮ�P��4ץK�U�ZMS���5߫7]����Sw��0�����'�|J�3L 0{���l	q����	��uba���������4iSn��y���zS�+�i��#���䒗��}��}cVIj�?J+�ׄa"�;�J�7;<_<�*� @�|D�؈�c���g�s�iq5늲<�=�~�EP&r# ���0�hJ�,F��5�����&��%~ltV�]��k�=q���������8IAyq�R�������L�XH)���9���B�	�tm������H���a�g^���ٔ\��Df������X16#|��IT�{�୻@�U�\zڬ����y��2ϼ5��~_z�P�8o��VEY�u��h�6⦍AE���B4&p�C���:R$*t5o\�o�ٜ� ��I�^�F僚-��m�*\��������F5FEQ��|��%
8�s�Ƀe�Y����f�ē1b][��|�*��;�5���S��x�� p��������D�p�Rx�����!4BzE��80$}G���G�ro6"�hA�d�u�ԛ���pj�L��f�]��9^^����`p85Z,,���}<7�^fD�Y�[�կ~5���?��@�w��\��t ��bK�	]s�D� :�,�u�H��E���{�	��v�"&�Ϟ�`���<�S�N�����y�;*��|0n��5�>>�Z>�'��9���9ZH)���*�n����&;�# %��y �\u��B}��[Q��s��%����S$�5��r�cQ�ʘO�69t���E�>I�F�Z�S�����Z<uI�JՂ=�0���V@� m,%�4WE���6_m]y��6'�0�H��_ZL\9�p-*[K�п8ɢ��H��.J�qM�t�a⺬�{�x����nڮ?��P�l����:����ob�����N7y�֣�&H�*��n�6����4Y��i�3�vx*o�Ƈt���1Bl���5�f��_�W`9��sՌ͓O<��b��^jV��8�؏�2����1�䲹V�>�ٜ1�xxe�h,�N*�g�c,�	pҋ�T?*���
�`��+�l�1U3�.�."vK*94͍Nػg��' ���~�|����|�o����O<S���
�YK�7�DJރ'{*��׌ �=��U����y�=db�1a��L}� �n�/C� ~�h��KVu��%F���ɐ�ȵ�	�Ӯ�&�H9~􈈐t:f������A�vB�b6!�rmUFJ����&i�T�Z$���=��Na%�sXqmaD	��^l10�|}��e�&f�3�^&���U�Ww��&��JQԩdI[O@9uo���9|���Ko{)�f�TM�)����n8v�d|v�T�x�P:�̙sz��o�V�'N��&5��w���)샎�ߓ�&�8}�X_�>�A�u�"8�.�*�7�z\������S����,�����O��miU��O�ƛ���/�#j�޸E�WU�ǆɵb����F�6e��b�"�G�T�M���;z�J�zI��q�Q�[Z7�vdo���/���o+r�l��ġG��E4o�6���v� c�f�m��������h�`;pz��d$�fRM�5��I��)5���ӑ��Ns�x�m�G]�5X]�L��+8=⃸!�ǚm�=MR��@��ʢ�����0�Z��<W�Ŋ�tq��k�뱦��*@��km������3YrUQ�W��|�X"����`���À	8a,�qP8��kiS>l�<<��#�i�")���%���J{��~?U�Z(K��1z�T�����^\����FJCC�:���(�@  ���a�~�ߌ����q�
�k|C"uv3�p9�`-�`�_u������b�{ۨ��0v]�����L��n�I�ҥ�����W9)>�M��T�3@W!P���yw���	c�a�s/$=�^�#�HR�����[��X�q�>6�x��ˤb
�@��D��I<B�O?��Ғ�������w뙐��e(�*5� m�C*����Y�^'e�l��O�Q4���*�uS;������kg43ґH�0�x�T���eyI�����#�D#�/��4�������W��P��d��$Rn<���@<��d|���8�������z^�ڑ�O8�r���1�^p�k�|��j%Xg��X�e��$XZ�J���dXYZ'O���ϱ5j>��e�S�Қ�W��!Z!2hn�r3���Ʊ<�����ˊ��-Y���Sl�|(K_s���|S�M��z�s��m�u���)�F��׾�UK7��ǉ0�eB"4D���h��o��j�ꛠk� ��L |]U5��r\#����k�R�Fy��j�D|���p��6����-��(���Ś�����/���@�H��XJ� m\
�Nsp���J�Ix��5���q��*~f��3Y��4��s<"���$��-"��kO1N|��T6N�R���W�,����+��7E�ft��p,�l��5#��r9	w����=���9�����J����	�IDa��@d!אZap.��9~L:H�#�'��b��Rt�^~��p��7�ߕ)[^�`�UW�n�|y�s���T�K9[��5 ���5*�D`ᐎ"?9:�&{4������m��'d	��6�1�RQ!y^�z��ɦKj�@�&�K����N�<��8 (s�p9�/"7�'ʹ-xD.�E�����
�S�-����~6����I���<��'6r7V�}�L�<�"���"6�/qO�\��ٟm��s=��O^���ė����*�f	�1]����>nl��fǋf�ąR��Si�X	��@.J���0[�J������+_�D� ��Vü
@ia�k���P�<���g��|�a|k��K�ݍ��O!�y�&���]~O�c�^w�����s̢��)mj�jۤ]��E�4<}��aRV%u��$1�u}���2�����ccV�Au!��&o�
<JE*�e*�}}�1�T����T�?eL�z7a\!�K� ����+�����1�$Ѓ!f���\%�cS�ԙ3���)���'����&�h�[�/J+urM�B�IK�4#m�U�5r?rM���Zw�&���Dy�SM�>b�w���#<�W#H����C����[��l�#�p;P5��)��!�'��j,J{ʺ�G�����! ����8��ܹs��!ΉU���fU�Q�6a���:>fv��3�~|,��]�M�k�E-���ic6���km�֍��IS HU�[���ّ�W��B�G�1!
˚��ĦNt�[�3��(-�� @u@o�W�Lz��N��1�k�s�2k�p2,�Q��v{-��'`!;#���@�4��(b���s)�i���5u���hcN8X�W�x�>?���n��H��5�oԵ<�������T����a`1r�G�ؾ7�N^���W���)2q�����]c]v'E�5��EKy��g8TG�������=�K���j�0��";L���$���' "�}=ܭ��ԋ�A�G�a���U�k�%c��2��/����(zo,~Gt��uo����u�Ϝ5DO�F<�F3)q����8�z�3C�)5���q~+9ܚ@Z��>IS#�J9ڑ��v\�s��L�:���ݹF6?�ZɹU��"�ς#_Oy&~��m�TQ<�����g�7\�Ȍ�I����h���/���|@�o�{o<S��_ "1!����Ĳ�/,F�!�FS�$���%�A4���#�il�r��ha�%@ލ�E
؜��]�^y5�VU�$�Y����IA��0� 	����T(�_U��S'����odd��)=��T���h6G�ױaMO���V	��T�*ҳ�^\��k^�kw��yZ,�N�8ԉfQ��:JM��K$�.�J��8�K+��K60�lڽ�L����VV.�W.[��M~p" ��r���7�u�&��xB�0�}��`��~��wy$�?�i���G�n�2�Q�����g�΂�K��G ��,�VH�[���r����j��b(��� ��@TQ�	��MU-J�l�������D�b6�����K�K�� kpϽwi� ŀm�`S��#{����%_�5�#��K������0�8V��
�順��4���i��i��Χ98�/"�D�ݩs��iH��`�3N��gXs;���^Q]���.�v����}���ܜ;o�#�p^)�a�[� �Șa�"�D�}����m����$�p���jrd\UU�ܬ�h��'�f��C�^�o����ؿ����Y�
�+䖚�yՐ��>��������S����eӓ����*K[P"UQe���M�F)$�S$��9F?��9���(O�d��_��?�6&k"���d�FF+��"׵���GG�4ج�� �xV,bW�㢞�"�o�Mk���-�r~�M7� ����R&Ͽ��Ϛg�Q4��es*/��"�P!Q��]|��� /\Q�`{�]w�SL��cy�ԉ��o|C����K�d�y
����T�c�ǂK	�ʬo�����j��R{R=�0p�=jDHޅ��	/�=�|s��{�-���F`IƸ���32�d����/���,	��J�1&=�Ր�RQi��y*@��M�΋Ѿ��0�u��1P}����j!��ܪ��U��;�;���;Z�x���7��*��5���m��_�?����<|oas�k4�8 glՋ�ԣ�v��n3�y6��([�ٛ)��߸�3kc$�x�p�6��׭�A�ze`3�����?���h���C*�f�z�f�]�����_���)����9� �O��OIk�u:-~x�l"���o[������pvx�KYv�R��}�~��K�-��R�ʤe����Tc���@�6 �����Ѵ����p��{�������� �����U��L�tV����'����\Wz)��]{����*U��>�w��±������Ĝ0�"ދ�*�
+\_��f�{���=£�n��k*�`��v�R��v�^�{�H�	ǔ �9��n����ލ���lX/UǮ'ef�_��"އ0$��F�U�2u|o���sؤ��jפ��0�J���1�cѺ��=H˃��)�;!.��ȑ�$��B>� 5�}k�`";۶���
��$7��0>;R�0MR�ҹg�$p1l(r � &'�n�_�Ro˥���8ɚC�q�Y�n���^Ό�#�
�fc��c:�7'�*�i�Ƥ'�;���ʉ��E0���sd�n��-���͆g�s�8�Z�ۚ@��ϟ�����X7��p��	��H����X0G�V���9(M�L���x�q^9X$&��t:�KZ�}�<��Q1����$�%�/�c�L\�Pn���݁9�'��<�=��]4#�
2U�UuC�����j�߳(�=�R�f�:KKz�Ti�H�oIa g��:yn�a��U��?7�R�[goo�g=����u��P�"O��F�p��$Ń"M;Y� Ct_��`���7ޠ���Sφ^xY��KD���N���Dt�mӶ1��TJ�p�{�g�ަD'NQ��诿���)��o�#^[[�ٵ��?{֗���
����F�\{<�3O��wH���=kA�u/���b���I�!�=z�A
���0�A��p����/����}X;��r�r9/���6��w4W����]w�����H�)�Y��4q��
�{���'�R��󪴤ꆔ��9��N�
��?��ͳT�S{���m�')��#Vm�!TvU��a®s�����LQԺ���3��U�N\��./0�u����	�YURC�(3��;K9`v>e7U�e3����K��10I������v�A���i��t�e'9c�z���d�o&���W�eu���gKq���a����qU@M��m"��'7�ȽE�~�
	�Kn M�Ϫ.��N��.��N�L���V=�,/��ox��ΜK��֖�C�>i�0#}���i������Տ�H���Y9�o�*�$�:Y��\� W�q���w]�Z8�H&�!J\d�ǘ�|�[�&CG��t3���E5�ȃ%��k���Aj������#0�er�&�h�Sx=�)��̙j��ǔ�w�"r����o�5�}�=z��W���~���`lI�8�|�k�Ss Y�)��UUUA<?׏)�g5�Z~x{����?׺ȣ��
�Y�T+�TM�*�����Q����VT�HsX9}�`��м�:�e?�M���W+u�EE��3*ե�2D�fj��-IP~����;ITU2*U�&� ]T{�i�G��9F7�m3�:��ܬ<c�������v���5���H�?GR�ue��6�M�ן{Q�S��w����ӟ�<����V� ��0Y�x�D1�����'�C������k怘C��0�H�R6'r^nC���a�#�{{^��_��0Ǐ��%윋�-ű����	�U됬x��2�86lF&!�6b6`H�j���m��&�/;���Ņ'��H��S1 
�(%��2G�+P�M����B������8�����U��S�J
���Y)�zf�9��a�����Z�����5�`7_�R8���̩S�����"NN�9�4	_��W�u��L�%l��h�"(��'�j�LJ���C�E%3���Q9��
:��+M�z�5D��4_Y��n/W�|�Zj�ı��6�eRפ��*�:�O��YK�R�'������v�V�{-�5=�:QXU�,�#Nb[O�+��w�f�,��͎�A*�����#FeCw�&�>����9}FaX��Z�QO$Ӥi�<��ƣ)R������Ar���c��A�9ha� ����}5��7�P+��ה_���1�� Y��?��q�)tĸX��9 ^b�8M'MZ<(�(���o4D*%�C�[��P�����Ź�b����E�^'���#f�=m��K�������}_�`!����@�n � �G��c��ظ0��T��,�3��r^Cm`jo�7*���j���qx�fd҆��=UJY�ż��1�K�a�)��V.�ЫGJ����I#Fݳf��q=���D��q9{�|��'VT9A��v�~"�7R4Ɉ�2�x���m��0����{��4��}m�8.0�<�ݕn�k�� B<�/��	6'�HwG�dd�����g�}&������5�Kz��%p��rݐ��狷C�ǲ&��9~#�S�� 8Y\�KL�쁿��@~���_��w��>��*�(
����f��#�D��|�|dݳ�)T �J��kq}" E6` (k��~���T)�V}�&��M7�$��x1���C���=k��i��)�z�H4�fC��qⳙĨ��wO�־�	�j.;n�y�*w옉��x.D�![Q�N����U�ZkX�6��H:VT�
� �SZ���w��eC�W�Q��|�3��ܞ�E�*��Ѩ."��}��[]On/�:U��<p�}�e�a�CU����Q��ͭ��׎�Y�m[g��3Ћ��=�إ��6$�g���"y�;�[�uɊ�tݚվ~ϻ��U'
r�J��Iy!���l����Is��I�{v.��h+Ul,iSd�j�͑Ok��_�y��дIa��!v}l��~�B�&�eC��9ɦ&LY���ޤ����J���T�Or�NR��J
^�e���)�������GΧ�k�{*��%�
�#�^�0��L��jyVn�=��¥���N'R���9�E���S�?_���W�����jm�\a$'3{�) �7�����<{7�<��0�S�ޣZl��qytn�o��<�������p
r����)52���׾�&��ƨ�^��^w�K��h)c5�.������a*�I+t���W5�鳾�J�t~�A#�:��� �FM��p�}�4�n����Q'?\Tl�yZH�^� WӨ7I�G��HD#%k��ʹ�ByY& n���h/��#�ו�
�L��K_���9�S�fι��J�%����^�z#M�Ϥx�fĩ��w��/҆#۲n:N�~H_}������%��Zg=���Y��p��JE��BܐuM�@�8 �X@��<��'��U
o��?�����_׉݃|?�_Rj����nP�7�%Y�1�y�����?n��6sGZ���h��Z����|M�غ����+��3�T~_EYS��_�����+#<��� ����Ohb�]��%_�L�=�~rA��z;���7E��~6,h �����䰢C�s6�/�"�U�o.�����ܮ��?|ւ�^2����� _��-��&����yh�+���X0,>6.�,~Ǥ44��ɣ�zx�v�&ѾQ5@�ܦ�Ѭ�ρ�N���R_5��G/y��P5��@LЄ�{�և0�n"�����M$Y8���g�N߃A#��x�������Ozy(�c8�m�:%�<D7�ߕ�y}r�Z���rx87����pȘ��������re�a����-�>_pXΝ=������JkNNh�]�0������Y>no������+\���6=�f e�TW��}T���������W��i2�����7�]����X>�y��vN�I�Ϲ�S!���� ��9�5�_+��J%�>��s�L�R� ��H
�t���$JCD�j=�xd|x}�i#u�_N@� ��Ȟh�Hk��z�"�|>�����2+�4����:�s�c
)�hbO<�܆"��� �^]� �w�~%6�Dvn��F5��p��ѩ����o�I%~�D^e����|ɿϟ�������;w��!,]�^�����<5�����M+ۡ�����'�S�_���ӉU�)ېx��$���v�E�����ɓl�w��S���-mU��ɛ��p���5k��sذ��l��B���P���J��e�.��ո�2f��@��M?�.��6|�y
�л�A�Q�]Ħ��f��W'�����=�~���1i&.F�g��d���H��G�{���]���D���v����p��߻��������s���7����0j}���]�-�:ґ�L85��?�?�����C�>>��d3��/2��w%��_ql�ְ���+͏���q9#:H������o�����(}�9J����EM$�"�}r |�z��FGQ��{��|c���x�{��k_k���gN�^�d��M�Sj�Mݲ�����+�2	9?�=΋r��;:�Zxx^�=���jB����׎W�2�)D�3�}����Gı��������p�u'��ޕ��ԑ*�km�H �z��+��7;��ȫ?����������:��j7���۷_vۣ.�N�a��T���Qq�u����|���mv����l�;U�/�CJ�T�ǒVP+eR�+9�8�]eYJ����[��ȵ>�ڧ�F�-G��y6s�jh7|��c$-j�N�(o�y4���䮄p7��en�J��H/32�%x Sa@7F�*^�qq~�#
��������x�����7��c�%,
�E���0N�8�v�g������ƤnEѬ��~�d��d��g�%�~��|�~ond|C�������G���O���`x���٠��ĵ>6�hl���^�F�v�~3�z�����@4�2�>��G)�|�^j�U�Ύo�o��ܚp�a8"�o>���Ⱦ#[����55"M���{?����F��Z 9V�QV��������Y|aW�����c��p���q.RM������s�T�p=Ncp}3�L�V���HU�����r��Wz.`$:^_iCo�1$�'���o�=��"�f�A�%]E�Ne�NΟu�l���y�ᛙg~�sˢg�5X^��J�ז���N����ܻ�Տ)!P}�FD����kv\��Ov���Qy,���'�|RQML�L"n�\+�I�D���7r����+g�o������n�z���äo4Sx�T�D?��� `������"��ۯ��h#���0������l*�`9���_�y�m�&��+��������sz9/ף)�8�Q�<�2��,d:�!����0�r�����s���7<6�;.Y�l�y��f�h���?{��e�U���}R��Q�� �$�2�Q����}��p���Ϲ������6l��m�D`D�%��;��9TwUW>��\��:�ϩ�Vw��K��U���\�9�wιД
�Ş���b�w��ۖ,����r����Sᇨ�|3�?�f	��$�"H���YS@������pΤ@�rN�MËuN�w���,u?\Y�iE�@H��[�_������j��L�EA��o84�%����Q|����V�7��t����O�;]+���Vw�g�	9V�jXj��/��85P)� Z""�����ɍ)��'��]��+�v�����\tx�þ,��r�abbȝ8y"�ù��	�b<��9724ↇB�"+�G�Λ�󛱈�:++��l�`�h94-BU��p��B�CH�=a�d�U��/�]9���N�AM�'+X hV��_Tn��H��js�:��Q�� �����`��;��̫Pr�L���"�, �&L�":`} @:?q�=���N�ZQh��u H۶lsgO���EbtQ���^\��L��.�v1�<%1[�����	4���]q����jZ-.�>W��kίԻ��*���V��k�.���V;�E���ʏnwΕ�h�X��4�cҍX�][.�4  �}��K�%GR�_ &�,����!�4%�}!Ũ_�i/�ͱ���Ҕ*Dz>�GI�Ȳ��uo��+*4m��� ���g}LD]$�lW�,K�C�]�����KmW�J���j�.���s��\6�m��(�S%��!�L3�yD#.&���z3��퐂C��CU+a�D�\���m�Z��<�+eR�9��R��r�D7Ցq��j;]I�R�l*8���aQ��4H���,�|��in�H[�����@M|���|���'?���9��m�&���L�Z�T���dZX����(�������P}��iw�ĉ�q�ٲ� ������~+��O�-֟��{�;&��i����v9n��l��i+.{���8��z���s�^����K��]�vl���{d�Fn�q�����{=Oz�bk�ߵ����^j�6�"�N��xN/��b@�W�{]G�/���4zݣ��6��_K�Mj!�R���^!g�Ø5y�PwE�u�<yt��.i
Hf*+���,�_)�����s4���a�:�"���""�xJ���UܧRȃ���v��l�$��c�ŕ��$�D��k��Y���Sq� �KB���)��P�>5��ჴP�.��Uy9�$�!:V�şg�gou�)t`�C�t�>��Q��	�LP��w�q�۰a��(�z��/~�����fgf-3/>lR���5����l� ?\R��w��`�;"}�_7�4�����m|��E�m����������^��A��f��h)WS/��F��^�4��E�8ϊ|� +\���<����h�,~^|�˙�KYz�r_]i[j��m9�������&�Z������I2Z��Rϕ^?X�Q��Sy��z#�v������W�޶Ħ)0�,���,%�4H�n���DC�Z��GY���;K\��@�������e�޹sG�4�>���G�6كywr��ZX/ê�D�*�S0�����R�{:�<'mj�d`�"���׫�_�� &�qj��	�S�.����-�Vl�"�F���)ڨ�)Y^�b���^�&L$��aN�GL�n�
(,[}@VI�'��J�j�]�f����I;��]g1b�
9aJn!F�����˺C^�3��c���幜k,�]�M�r7���^�s��ܧ�!��]��s��h�6��ci�`h2!.��MM�����y��X�{^.Z�bq9�Z��k)��Ry��ӊ��\N��Az1�i9�U\3�G�ތ{	�ś����5ckB����,�Q�C�,4!S���%0���J칔lN�Kl(�(�(�X]T��8񺏲�s�-[69b������%{����b���5C9����|۱��x�C�D��m��$�Bǹ\H��_7sT'�JTc�'����4�4��j(�]��f�\�v���7��8�YH�^J��Br��z�e�g#�&.2,0�7�$_��֨��Y��Й��F�F!��Y��Կ�����+�^��{i���.�-������j��������qW�5�Rm%�/]_i���y^����{��j�pW%�֘��ե@�����s��*+W�2�ෘU���@}��Z�R�V����~�z���}�$�=�('R}ܰ�#X�w�c	_?s��� ��ⳡ�G���Ŭ���)þ�a�gV�T�v�3)!j���=\��H��9h�p�cd�/ňX�x)����kñVZ)�?�L'D���t|~��j����R��U�լJ yZӂM���Ćx�sSlw�Rע�FHB C�䛞	�4���B̷ ������Z
y/�̨�u3�e�1���n�����{a�I-F&<�R�O��mF�aJF�u�~R�$���̲Nd,|�y�1�{�q�����-W��;�j>˕�+��NW��.wc����m=�S;Q�
�t:Q���t�����c��yn�Ǫy5���uH�@�����7�p���G>���>�:B@��$�Xn�n`m�u�� ��|����~ǽ�ҋ���Q2����jk�9c�VE������`��{391i���3z7�UJ�a ��k$� �nńG���J�������3�g������e�?�A�mݞ�tnu�Ҋ��Ժ�M���t G��h4��fD�� ׌?��UbJ���<7~"���B�j�_$1$�!Ƃ�h�N��\�jĭ�_9�7�L5E�Eɼ�&�����G5�抋t;����c� 9B�����m�n���A5�+�~I�մ�,%��3����z�ׯ��^?���BS�+�˱bȢ�߳�fR+I�� Q榄Y=���Z���$������S*��)��rν�cuLj�H�]��¿�<E׿˦�Yg���mW|�^��1�4��n��V+���}�
�J9�(��g�AKzȚ����r��+^I_@O �)̿�A�*��w���-2QS�Y�D]�T�f�q��[��3�*�H��έ����U{+F�9$�U���?'�Mk�]�wY�	 �(ȿ�к�͡�g�h�t!7�A�Cp��iV'��&D�hO�7 \��D�XG�;e�5��ʵ�78<hd,A�RK�x+]��hXpY\�u47L�VVkMV6@cum� �S@-dͬ����RV=�WQO]SUz�`K���r$�y���h�=�X Z~aD�����z	����_j�{Y,��r��gH��r4\����b%\aW�Ҿz��j�Mq���.;I�hj�Yh���:L粔ɓ^�^�s��奟²غ췖u����y�?O�v�ۖ3��@l1�H�.�z�	�E>c'�Ư�گ����#��U�U�����i��@۪������8�jL=�y� �[v��&˚�Xg[	킧��]�l�E����AGc�b���V��?��Ȩ�W��w�ܔqv�$�ZI]Ӱ�z�WC�[�G��dp׾TY�M�/����M�@��t,�.�6����SSD�2���W�H~0�A�%��U��	��Ispr�pLvL:Rk+J���`��cap��TRMNϛ��m X����?����'w�(��g���1[�-V��]yF>�=C��E9�LQP,&���Oˆ����I�JEp?�Y't^Zf��R��Q.�q��������Fm��l� �l��]�%9>DX�M&s9�)������Z���Z$�s�����-l`��z� �+�J�xK��b��%}eB޿�U�&��'MَQ�9��,Wy~%��:�z���ry.���m��k*�P��b�d�|�D%+�i{���艰9��u7y�+�C��9�Z-&jv��B��X$���T^tS%o�f*E/����������S~/w��v�EܒX�_4E�����ܝ;���q��%�3@� �Ui��Q�JK:X#�T�D:Z�S�6�"�*HC��@��w�^w���Mp�i�\0�\R�7K];�DKK7��F0jO�g�ݕ%���������m&��xaRS�c��Z������S.wW�������>T���@�o�M?KsѲ��[?�����-��yz���Z��7���K������K�HqS��&�+J��on�fi-w�~�	�z�o%�▒�[�2�&�K���c��p�Ά�Գ�����\�����K�%Xh(����g������	_��x��)��;��l�����$�IwUp���B�%�� �+�����3�	�����j������*yP/�?Ö������nط��~?!%ȅ���ɍ�YkѰG���g�6�=���4�*nr*d�?|��{���v{v�	�O�:ΞY�=	T`'�I�2��1e��s�t�V�����NQ�G&�M4�
�q��&�;pxd�@	(��UN��)�.��7��B�H��&N~��eJӄ���&N��h��$QU�b��Z�|���$Cf:�L1K- �3���P�V�"�4��2���i.	(Z=����~�r˕����r\?+�o��_�=���5�ۚ��z�_Qa���xP��֮4<�ӧ��x-��^ou�����L{�p�=��O~��]�z����i��������w��]�SR�/�;-��W*Y��k� :�m��fZNa���Z-TK�˂ު��� ��׎X�-WY�n�Y�7lX��-nj�W�G��:몵����?f������l.XA�`Xp������G����y3<��f�l��JͶ A<��ªd��M7=7c��s�c��r� Ը�N'� ��0�hQH�"��d�К�_�~�R�g����f�NV��~��$�9�<��y�V��y�G�t4�|I�G��*��2�ٵ\���X�(��Ȍ�Y��O/N����iFi|4��+3pj��uҗ�TqV}\��镙�86�<u��P���'�|���9���zi����������Z��=��nu	��do���JZ�"�fooT_���"����*�,=�ϴ�=��������yzn��]n_.e55��G�M�� �w�d���l�O1T^��E�ݖzϢ��h�������Fq��|����e\��ȑC����^�r'����hU��?Kٸ6�Q�P졋k�/ejz���D~�
�J Sf�ܹ�&�^w������/���9O�:�N�8�,���uk܆M�Mo��\R�Ύǜ3��d�x9 xց��U����~yt��9DѪ9!ٸ�B�ff9��=M�]2�#�\���C�4��k`�ڪ�tK (�;�|�on�P l`x�m�f��l(�5~~��3��{�M<��p@�
}��9	��pO�����K@�U�����R���Xo�Hw�������o}�+�uR4'�բR!08aU��;��"Ź�y,7\�Ź�_��)��d�/������?��<u�ɥ���I��	�﶐$&,���e^O���'���>�l)��E�&L� -���_�>i.:0)��gȣ���cE�K�oK����b_�[L��<��+q.u�^@t���x�帄�D�^ϝRM�Q�ߥ�����7�G隵5j�/-k��C
�	i���N�Z�<�3��5RE�\z�{}�-��n�a�>�xe�-�Y�A���<Ai�����^LQ*��S�Vħ�%��4Y,�z���-�O�bmS�R�m��^�d���V$R�E�6�6���|ݎC)gٰq�W�wXX7?Hz�>\Y/��;{��[��ϭnvn6�N+ ٺu��O�rξ�gX�xo����!͗�<('Te�7���_�gc�Oy�ų���@|�� 5�6�4乙���{�k��4.
�t��֯��n��V���@���8P�V�~��d8`�D�@������������z�����tYg�6�L�hUIEj��	��#?p�kF��q�FC����291)bM�<�M�� ��<��ȥF?�kF��zi�)0�����R��)oI�!�j*0�Pt���kZ�l�uR�T�+�+��"�Iڐ>��W����r5$T����_���=�x��/݄��1z�^�X�v��~#@�J�K:�����o�T��i. �����b�}�K��fQ��Q7ů߳A��[����)�t�N�K��&Y�����H�����S� !�`�^�S�|�Ҙ�.��8�rD �W�b?پΰ<���� 7@ȿ=��o��-. �RH���o|#/,�\sAr-<;�+d�G�K�r*� zH�G_��q�)�V�:�{˖�n߾}f���w�w�=(a?$�{��]��H)����'���֭�ܮ]�ZTR�d�:��o����ب?w��"n�j��5������E W���!Vݻ��a��v?G�����̾A�j�/���|�ƞ�tӴ��Ӝ�X_n������[Q@���'����Ī�U��ѣ�?���l�_����>�9B�W�^z�%FV����/�Z���-&)��s|�J�bY�u�LH�D�^V�g��W΋f����ܞV\@ʞ�Ki?��E�c YH���1����u�7*6ʹF��3���p�,VO�O���9���qܓ�g����p���.��'c��f[�M�N���W�,m�ѧK�~��Җ�퐫g!	sO7������g�No?m/�ҖnR����Ӯ&(X	�i����Z�i7�.�wo�f^/e��]#���<W7R���E� �<�9gC͝�ڒs 9%@R�T\���y��a�Q�n��59����5�$��c��`y�a8��E>J��hpóv=��m�Y��m�f5�x7Q�fm�� �^%pd��<1���`��Y�RX3��}9'��SKׄhm�����{�=�ޜ����������L�U7t2S@L B(���3���v��=����{��ߝ�3�Ӑ�<�t�7�����N?�}�Q���m�֭��=l$]�L��߇��3h��\���q���ǌ<<8X��Ç�ɋ�y�r4�9��hf���e�jD�ydV�>5���jo��9W)�ݮݻ�;m��+���[��b�F���$;L�dEE������Jl�����X��İ�$��M��B�����"ab!|����o���Ɓkâ8�??ᑰ��z����Ҟ����C�*n�ϙ�T�w��� ډ��%��i�M��H�̈́�q_*r���y>�쥅,SSn�M��=���W�W���1�xN�URC<��U�B�VN�������{Ϳ[��p������g͍��)H�I�rA�L�uĚJν�����*,e
��7/ޫ��XmEf+�tGb��e�)��t��������,�`c�������~��O�z�5���'r�"�?~�C(�(%3?��{���Ɲ�W{�8_e�H���v�m�#��{���n2J�F�"�e�ڕ���d�R}?���B�����G��qf:$-}���g�B�,��k\[J���r��P�T�"S9ߢ��g���ʃ>h�s�Yq�R�x��J�g�����n��Ɯ�������c�X���g�������p���������$SBc�s��}���T��������f,�iƀ��>2+=iJ�p��ĔW���=�}N]�9��n���#���޶��ôZv�f3�P���xvV��Č�{�;zܝ�J!R7db\Q��U�t�p��5/ �5kFX�~΢�f�*u�x�'�,ڐ����|�L,:�In&,����1�価�!R?~Բ0r��s���1Lp&����ě1�cp5�0 8|��5�!�)�J����>��B0��/B��@�7�pEB�~r^������R(;��cx����h�:C�z_�������l����~˵�N�=�xp� UZ�E!���P�V0K���W�ds]�d��/��^�AO�P̮�N[E��Ag�b�ZA��H�KjyJ�LzV�7�S�(�0�I���9L��X��fs��s���ʒ�KA_�'�p�,�I���o���*q������ҔA<'������K뤵WJn��G�_�)�����j%�1e�2�;��ce�;7u��Բ��UiK߃�%jő��Nl۶Չ�Q*u"�:�Y�C�����B#j�T��3YG<Ϟ={l�=��SF�����]�\���������
y�t�,d�u.Z�J��"�[�� �?��\��������=��)b��
�n$���X ��?�qw�wھ�;�x�Ҁ�T���v��m}������߃jN"E!�7��$2�(# ��q���2��
(�ϡ,��Yg �P�W^9�cAŮm֕������W�,<��F;7~��X߸�������K/�d}�Ն=�38�b��d���{���y�G�k ���/kg�O<i���[Fl���tU۪�tkK�i��fpL�Ml�X, %ą���ht�Jf�I,�%�0?�`�A�͡C�l���fHԲ�������;==7�`.k�:�JiI�bQ	ɴ<m�������8��l#$���CC�plؼ���;G����r���k �d�`�ǿ:�f�齅��A+kX�m�	ԃ���h��Bٶ}�ۼi�?��8@(��j�^y�Y��϶�,�񘚝�-0u/��3h�$�B`����</�Hn53�2������G���������pC�b�1� �y��k�_*[y��%�h=\�#@�����![�hc�<�崕�� X_����V�u�"?#��=Ns��t��[G [ �HHM-t��Aߥߧ\���GD�?�������d}�s��u�ꈇ�5 �V��e�ȓK�0r�<���!Z����,&e�7�y;3=��X���w@����\Σ(�?? bֶ����V�\R��ܫ�t���A��$²�O�����>
���D�
)��]�;�_`�BQ�q���&+�XO㫱3PX������o~�ޕ��&��R$5�J/�rw��]w����[���<�?AM�W�#7+��S��з(ՙq*#���[9�����{���>��Z%���Q���Wp^����qs�ubΛ�O	�ff��0��`�5[f��X�1������OG6��<`Ɂ�ɕJ��� U��R%�(�VW.�(�&mZ��4T��	�d>|����o�c�5o����ݨG��Q&���3�L0�1�י۩ef2��[�r�m��T�`��>��m|?�я��S6�+��EbN��&K������I��;)WN�#U��2�VPB>�	v�]��4>jE�+mEWT�穉�\7�Xp�0�rYh'_ho��\��	(@���0n5���j��7lXo���nu۷m��@k7���y���?q�N����=,�,Q��!hW�|ޒI��cm�5�ր	[$q��={��?�~#�	3����w�}v��s>����k�.I�KF���T��l��׻�B���~A���?6St;�R�����D? �Gꪹ:\G̬��f��Y�{�.!��G�>Z���E^UzLQ��BQ�p.�l�^.��Er��k����G����D�2?�-�3Y���A�b��#[8������1�.��@���Cw��Y���Ephh�o��xl��������Ѳ@ �����ݵ����o� Z[��<��S�y.��V�z# ��2�10P���������g���3�R����7m1�?������؊�E֕��-����2�5���^�̕e�D��"��A�=��� K:��~�U+6��\�d.�lPı"Nx��yx��'O����9~�D�7�x9v�;?~���I7���S~|FF��~Ϟ>c�"�s�g݄�(^��l�b\,H�nJt�2� .t�f&�{L��b�V�+^)X���d~+l��wm  ;�µU#�E�|�dZjҨ �+0�d�M�3)��@��Y���ɀ�9�5�[��ϝ�9�,�ˤ�p�汣��BR��s�u�ٵ�!l�dw�����q�O�����m�v;��OyP����<��Y�5�̤��j��Y����	&>���#� ��2��Fctbn�I���+"�Ol�!C0�H�T@K+��e&VuE8������SO?m�e��M��>��G>�v^���7�H�mzz�MJ�SU�W^9k�z�}�Z��ɉq�)�`����� �F�m�a���Y�E Z#���G�ouT�Ƈi����W~�W��w�ωl�)�(����mLS�} B���<��F���hw�?���W%�z����q�/|���i�|�;e����c�S��Ew��l��O��DqPrҿ���&���"�i�ռԸ�z�T�8.�0���˿l��q6F� ����6Wd�)�5�7φ_g������ �.�w�%ι(0�gO��OTh*O��Ș��'���q�Z�p��ow���w`��,�!+���LC>�/���F~ �f�/��d�!Bt����mMf�S�$M9�d4��詧�2w���V�$e[,�Տ�}7\g�� 	��M�[��4�I�w�Gy�dc��{���Bi���^!�eQֶZ����E
g0 ��	w���e.Y�ކ�� ��\���#̈́i*c�sc~?��Y�̋��͚���/��"p
�r���c(��L7��g�rS��^���z�iE�c�|4~�EAy:g �k�̵�@N�YeC��䩑uBr��L�Y
Z54����3�H <������y��ς�0F�0���O?c�QB���h︄��L	+���Lz�z�3�fQN��$R��V�+.3�&�*m���Ix�߿�����H4�]�U���D�-�͗�d)��(G�^V]?�,><7@ВbR��p�_�*������G�jR�U��-�MH dO�9��٣&_�R��9X�a�6�(�`�0o���Rҙ���A{.{Aff~f�0�����a��n�Z���������;�֭.%�=>�5^�����.��!�Z�^���;�ap�׾�5#�M�i�{��r�����M)��p�p���?�������.�H���,FD^	��J��x�~֟�E���˹��m�\7�>҈�sk���x��.��(�����y�N��Dgo��-��`�+@A)lMFk/8A�\$�dV�Q���r��_�:������N{��W�\W!`@
9�0c6�@v�yPt�{�{~���}�Փ��`<���&.�����"��\0�E /1�,���+n��?�������]o��D�Oy���s�&��r��ݻ�u/��;���7����N�,LdQN#�L�����,��;��S2�	^�F4$#�Y�P& y�ؤ
�~��sC�,�$�7�\�(m���c%
r8(�X�Q��@����Y�֕�'N�s���;�[PE��s���3�1nA�`S��y�Ty�q~h�=�m{���y�"�ؘ�q�����J(�����S#�DE��dѹ�O6ZI��ʫǊ�CC[�M�A��#�9q��f0�GgZ%�8�0�=X~�kA<�C=�5��y��30��G����$���\�S�^�ؐ�H�!�M��D@�����l�X�xР���@萞��JV�d>�)��	�Դ�[I� �p�47yA��4���f�\=d�y o�fQY���?;�x�I��бZ���L!���M/f!���0Vs�i�,��������ט�9hhy���h�= �g���2�(kwR�n�hM��=ѥ[�&w�>��{��@�$J������m܏9&�ų07��+��_�y�;�r]X����V|�^���9֚~�w��=���I��ŏE����g֩f��Ͷ�Z�D�չ"�*�G���9��PE�������=���O}��+��R�ԤԼ˃��;v�Q<�{������k򗵅L���_���\�u��B���@s&������@�;J�Zn�bC�ar�2�����"�j�΀�_��GC_TBT�?%o����v]��_?��PV�oX��c��,a\Z1����P[i!_��OE��BwrefϞ��rK独W��K&_8 � ��)ޒ�?d����R��K���{�c�E����q �qޝw�i�f,D�s@J��sV���
|H~pC����̸�U�=�>o{W����>�'��c%�MG��m�Y�i�#����j0�r]m�lU���Be�9���p&�E ��M�oZ�=s�m۾գ�!w��o<�7�7��߽�BҸ�ڋDQ��G�g�\4+�����4T>�f���p��a��ϒ��r���p�����3+g�:A��蹄�qK���H$R*xД(]ׅ��L^�1+�6Iݣ��#�=�B#L�Ze��BŢ D� �|m̨)����
�r�P�;kjj"'��k�(a�i�?C�!�U��3D�W)c�l�g��BЈp�5yH��XZ����93�_3��"� ���E��TX�@�����\��ć�ǻ|?�����X{ 6�up����3�#@xg,A�y�{�H�Ԏa�j���[�_S\/��Km��U�:�j��z����\\���"'��y��sNMtI�rIqZ�x��o޲��|�����1*6�+厢"�ȺDcWI�S�!��R�{`ú5�����;�� � @	���\g�`An߾�ޕ㙯����ᡱ>XAQ�aV�Y]��:���y `0*K;37�t������L�G�&�rGdhp�6�����z�%�����֔�Or�pJ�5;w�k�w  ����[��ܴ��r���b����t'��7��n��f���a=��6������~�oӹ!B�$}'+�z�����(*N� �j ��}���7�`��9�yXy��753��)U��'�j=��-�p��2W��Q"]K^�ï	������<:��~<��=��	�0\)�~��V<�[��PӢ�r�B��d5��B���b��^��Ӡ�p�	�ظa�]�����0ǌx���w��
 ��U� a^����:�A�0,r��Ǡ�Q��� �J���"^�H��BVc�, �UT�����,W�s��A��^B[�D�����q�r-�>ye�L�����D(�b'd�jZG
$���T/d6ر\���s7�[3f��a���{-o�2�I��5�b�м���u%M!fڔt��{a�7�䵣�Yt/�M�LBI5@$c(}��^yH� 6	���,vc�{�s��A�s,���a��>{��1S7���X,l�"eJ�ui�\��/G�_	>�J5��vTӲE�K�:�,<��C��O�zro�$�^���3�y�n9Z�L�g��O��A?�mnՎ�Z)�iܟ9���J8�&��O~�\��US�k���5�3'	)���<T ��;ޱ?X?���<��ߙ�RXo_�e.���2;3�m� ��#Yr���m�ͪ��8t��;u��i����L�@�	�r떭~�n��&�5�3ѳssQ���J�;����#�߾?(0��fCO�k�5��	w.(1ʯ6�U(XJ��0!��pN�h"O����T�l��@�1�"��R:�86Aq���B���%��z�<�E��{y�����\u���;~ꤳ�2����s*ƨ��u���H��+MV7�w������������ڸ~��/:��z��j�	���Bc�W��
�&�e�M�\0���}�1�S&�t㦍�Y�Y�������=�X����=�r<f���Y��_8r�5یJY�Ls����p�?{��!NFg0ndz���[�2l�->5��t>���� Hr�`a�)322���Ԥ9�%Ҋy Rӧ|�Ūܺ_QkN]�E�M ��1BM��?7�6l\�Gs&l1�C�����&Wۏ���{<du�xO|�'N�4���/p����y���?|�+.�Ul�WK��Ga����s�_��6�/:@�ރ�Zؤ��r<2�b�0b�b�@@sMex��yw�0��a�[��0�÷�J�p������/ɀZ������\�`�ea(�Yq����)~_lK���rO����{�t�H߳�R����:���K��AK���ɺ��\|�4�Q�uj���(�����jN�b�}/#T?����=��܎����F5Z�G���a����ꁳ弊�'����<e�A�@^7Rh4�^~�dю;�ƒ�E�,6dx!(;ܓ���S̲�is��h�X]�>����6�5�;7�[������?�w����p_�?���}��������m<ĠwEpYkp�k��ؗ��lC^�f�)�R�C���;}��]�sS��|
�@cIFI��\��C���ε�Ɛ�P^5@���C��Pc��5�U+y��||bj�d��,���O,4��3�/����I��c�Y�J�����X_�H`���T��=5c��>���g4Y�<�'��5�	߂p��"̽՚�#%�07mQTe���N� a���$�h�F���dQ�[�sY#�bGYhl�i^P��|��n������O���G�A��|L"e�E�t�`'Q-�\`5b�����I���R�u�Gn������V�&��3l~��0k�hА$$yO��_�����������e�1w_�����VZ�T�����٬���.S�-ラ�Z�aTj�Q�04S)�4�_$Yjz������-��n��O�qӠ���������j���n���Rp6�|���������P?�g�#cf�<nQk��`��R^�
����kĵ��*ԐkqM��x�t�jcx�q�0�T�JT�Qm�2�}��e�J�oDK�r�Z4=,���H����[�t�4Ǌ��^.���-���9z��иi���Z�r�
�bc��;m��=@�w����)��[���\��܄��q�M��7c�̷��-��[��=����컹�uJ�H���Y{(9�-��Xt�H��	���|��J\�_�lz���ͪIɅ����J�^��?gYvQN�y����ۧ���n��{ܭ߰���rclͨ�wg���uF��w{�34<��Y�^9�lwq�c��_9𒹈�u��)7@����FG����OPv��*�}�����}�}��_5��]���oS������]�|����>f�2���w0:��hEߥ ^�����8�&����%"�	�K{�2W]%&PdJ�7P3Y����M�n���
���u�P`�f�P��
����f+�-i�^f�i�
��Q��O�l�oD[��;�0��pYHh�EŢ`p	�>W7`39q�4�u�ָ��y����y�9z��1L �ev���Ewa��� |�h�f!j�bR.4��X���?�q�`�Tm�4=y:!�dNT$��L�� ,����#,/<��	�ǠQ�%'�͇�KX��:�EXL�����S]�J8�g
���[�-$AK����9�F����L�����?�gĽA���c�� ���`%C2}s��+�S���5#lH��0N܋��Ո�<�,k�j�R%'&���Q���2]�T/k���!�\	�R�_q޶,wĄ���I�3̽�i��"tId�֌O;�>,R�p�u�fkE�}�/-�{id��F�CK"�<N��?��γ���+s~�i[γ�$�33�0��d!�6����)w�jj�Y�UlR����MYA�8��@g��2����;�8q�m<�S���m���A�W.H� �i�.E���֐��d-����-Gr+�ly�Gp�l<v⸭ad�!:lRu ����,����'�ͷ�(��j
������rat4 (�n�k׆�.��H�z�X�H%Mǡ��[/f����Yo��� R���,זH���JR^ �$3��A�ŧ�����'2�zz�-����M&K�,�4<�ޅ�U;��]������"����#v;�fL�bO�~�jfU/�le�`��oH�G*�=���`屝���	JK�a;�9
-djzƍ��}�1Z�܎)Cf��Р��Lr�0yj�RA�1������a�4-����*��M�/r�P�z�b�3��y�s! ���5����jܐv����1�-s����)� z�_YK���?]B�wa��e��:�	+!��	4+�[ �w`���#D�y꙼�Z�O��Ϲ6��	��������P������s���$|h�&7wCL�o���FV#���|&�� @$��O�=嵳�ntl���I�Z�>�7ν��
��;0d�3K� �� ֵ�i�
!`9"�S�E! ?7�1�hA��n��2.7[��������V�A`�'zMu� 4�����B��" }3��s��)u�nq�R�P������D���]��Zt_��4K�ry5���wEZ�Kn��-Pjzv�����e�p�/�xW�u(e���z�֡e�n��e�-U�5�|�J��݊�Լh��*I���-Xxd5H#�Pn��X��h��"QQD����d>�0"��U4�W��t܃�t#�����kG�$�P�e�U/[֮3"���+e#i�{�5��� +_{�ɜ�X!z[TF-���%Vu�$�*��������wX�V)��	JI�$zq��d�3�l������:� �~Q����ȭ�J�q�\�Ƣ�Y(Q�0R��kY�F��K.�,�Y
QN_d<�Q��b�����G�K�����~L���بU��(�R��Y�c"�`��:Vж�_�Ui+FN�|��a�(}=������l��֯u�&@hΘ���a�&0�7WL�~���0A��e�����[�i��-�&' ����Y�g�fN���BJ&M6�9�V¡A�BP�� hH�-�)�����(4�����߻o|��L�^)O��֬�y�J�7C��f��R�+*(բ��{S�ރ�F���m�'�D�,��3�R� Z�R��M��1*�`�������mb�Y����o��k�=���̙���d��hm6[���}��}M� �(ñ��D�����,.s���'� h��{@_����3Ϙ�W"����5�d���r5[њ�z���EF�����u��]kC���k��f����K6`� 	���3%��+q�rAE;���Օu��ۮ{,R�EQI(ZfӍp�~.�E��"K��	���S)�
��nl��y@	@D7"w�z�gn3,�~s'(�<�3�/�L�>��f=(Նj��Ω�>۝�-�A׈�OJ�QN� A ��:r��~םyet�X ��jZvZ�$�@�,쮝[$ԇS3�hȠ��ĕ�{�5��g�5;�]��W.U�j�f�O�ݒ۩�M�\m��!���妁�rL�Ǽ��J��)�P��-�v(�����ܽ+�Գ��!��� c��:�W���8�M�R�Ω6�?v��,����x�,P˼ GB-�x����8]����
��#A����鿆�L&��I���V�t�U��(Y�\.��T��x⤀�D!gd>?�'M�b����j)Ʊ�0xlzd���7��B��![o
0�D����j�� �6\��4�dbT�IiQ�����,�I[��t��x�	�F�\s���)��-�:N���m�f�@ދň0�z#W��ǀ9X� .g,aS����=ǩR6�=YDj�p�-b˭ ߠ�V��F�5׌ij����?����*�f!ʩ,1���5�6`f�W�VK�b~�ȧܶy�D�����c�ffPx���PH��F(H���?��OGs:s��\Y��.��7�NA8���ڛŒ��3���k�9���|)��\ �D�W�/Q5E��g���L�9xg�E��; �������Qg�H��@���
sau)Q�4;L���M�	\�螒y�w�M������4��}�ӟ��q�Oi2I�/`֎ N����7m�h�T���W�:��\%ڜei6%������*f�s>��?s@���d��nqk��^����#D�_���Hf�Ͳ0�7��|�,5f(��55��;?7���z��Ȗ��1z���V���s�q�ۓV�{�@�{ʲ涺��J�].��l��I�T�p�&��H��k��R���r��8@��D(�=�}�a�Y���-�̌V�M��%}g��B�-M6m�`ܮ�vF,n�ږ5#Aj�?�f秬Og<����2 �����1��t���j���W%��~�i�QJ�("�tA�¿C�?��_<j�<	)s�ĉ\�|����'���1�D�)w�T��J3��I�:�Ҹ�Ş��:���j�I�I͊�0�����cC̎)��,!ư��͊�V��K�����i�������P���b+FE�;���b3ǌ��6��e
А�;�ɠ�t2D�U���>�pі^y�e����l����cC��������`a���'�w��w��I�N׭�h�w���sG��1"p�|�h��(�@�L��?��������g�}q1O(���C(ÆI�7(V�O(�6l5���~���H�1Gy��B��r�YݝH�.�@��ٛФm1^����zE&[8��Z�|"*�yNRL@4}̘|���5�
�Z�w���g?����Y[�����ȝ�Ts��"�`���îs�%����.~g�k����яr�j#M#�|0��F�|Zqn�/���q�Gc�˚���Q��_zY�Kf��y� �X͆�@-��]�z���;2E�'^��ҟ<]�1b��X�呣GM�!\�ό�,DA���x_\��X$҆��g���7�bK#����"����4��2������%K��欑%&���c]+,R�'�Gc&�M_"�)�.����>͔�V�X��z��	r�̹�,c[w�2�. ����R�d����-�-X�ݘ���˚6��pN����P����Pe�e��N�<�^;~ҍ���^���544j!�_5��.z�u��W-w�j��ʫ+�V�t��n��,���HXd��!�B�;.RM*U˕%���X6���w���A��M�2���>�Rv	Hг��TsS���4>�9�ؿ򕯘+�pE4χ�i�C�],�*E�44���d:r��i�iV��k���(��p(�Щn;�q5e�335�X�r%�)3=��,�a	�%��w�|�/�ϕ��"��g��v�8c�1�T@�������pfφ{��'�7g!��&������ީv�Ȩ��N��>����׾fdC6i=�y�q^�{���?h@�Y���X�7���2f\W�i~��"�d��պv/�Jj�W>��*KB�q&k���ۿ�۶��X>���Mu�B���v�=�mݺŬmaY�p°D��g?��l&�O��#��w앓�j�+מ���|[�A�%7�����
X�װ2/�A�g&� �{�y8��~ޯE���q���i+G�~j�S��R)�cX��7D��	n8�S��A�n���淾��gn�>v����o}�[fYPd���j~�P�������
��`�U��e~ ����Z�~���ć� j���i(t=��%��Ӟ#�ε)CA�C,�"s�o��!۽�c��
He��U��yV�yEp�)F�Pc$�ʙ�]�����e�@�� gb4Tc�"^�rٌ5�*�Y� )Xf����> V�ڵ����͒?�u���7܉��,WN��� `Łt<8P��Z�ϳjd��V<�I�Z.i'����E�@3�B���'���i6�/�Q�O-�<�3n,�d"�Mn�U�@��韅��\���|�͎v��ӿ�Yl'c5W��
o�¸���Jps͉H�S6Pq�X�~����~`��v��,,(���c� ������*�+M;Ur$Uq�ˢ�&�P7���;��܋�"\�a�Cf�p�𣢒�ϭF3qRe��W(k�ݩ��3)/���V�f���=�;���"�'��oUd]�%�}���a�5u��a�+H��y��͵��_)�4�z"�S�*���T��� �ƛ�*ӯ���j"Ƴ`��ź/�5V6.Y
��e�y �M�F��स�O��\�?ـI���	���FS��Y�z�_zmr] �� ��5Z6�������?��v?W�,�lz��Ysu�Grӏ�'�C� z����F�Y���>���LY�k>���K�>�B���5Z�D&��]��ts�֟�J9�@|��!�h#ȗ�^zŔ�xy9�*�e�4~�� "�I��n��`rc��5�G��RF�\~�VW�<���W� �?Xc�e�m���UxL���D�	���6��۽{�}���:�h%�Kye��*��y1�_�:�Nh}�S���ح��m�u�>���}j^N]c�#Ɵ�g�\��T¸��*V�y�i�v�%H�E����9_o�C�_�k��W��^ݞ3���3�p�_�ݶ�P(ir�;�V������Uw+f��GJy�_io�BR�u�S�4�JO��3��'(���v��ҹ��L���>c���eh��"�rZ���h��-��̏j�6+kZ(�-�.I��d0���2fY�	Yyf�6�`~O��e�,�~Ze�����M��B��WNìf",*�/�B�b��.Lf�X�m3c�a��~|�D ���%��0a�I�2�g;j�݋_���
D��Yl����Q�b�V:�Μ9k�&��7��$��k���Y�ٕc�.�g�Ν�5��s6�{:���'>a��-B�>�u�M!���ħR��#Q��/�����qM^�5R ��X'����.JM 0������̦öi�ލ2�2N��"ϊ�ϓ'b�ѭy4����r��3��R H���l���v��k\.85�N�#Y�R&�J�B�_T��$�/�Qr6mi��?�j�,�c%����.�8O
@�U��2��Y�E��H>w���q���h�re/�j��b��py$�����>&��Q�7�"b���L#e�'�ވ���M�|�f�w��o�v+O��[�D#V�1D�a��~�dǗ��f�V[d{�ɓGͭ�p�T�y	��,E_�-�~g�?5�eߟoJ�?t�5[���}fݦ�'�y������:{vܝ<u� �.�l����*�7C���?o����=����*λ����05[w�=��E�n޲�M�\p7޴ϲD#��7��-�Q6o���f�`�F��IB���T5v�E^Q�S�u����tjuP���`xA	�GAs1�c�K:O�w�,2���L6f�Ǆ�uh�\K�Q�N˂��'\�&���u���$�\�s����������fw���)�1+s��&��~�_4�k���:��t����HS���)p6y�s�(  ��IDAT4�/����OE��u�b0��X�>��4X�����ܕaW9F\�ui"ڄ�ЛjʹVKZS�Wo�@Qx�����@�����g��סi��|�&�K�waL����һߝG� ����wW��gC���f����4l�*��55>�+ �g���U�1�d[措_�T��j��%/�iC��F���=9>�f��{�0����菬�������4�?������U���=�	�fݪrqZ*$���m��_J�c{���M���d���r�9U��Y"'�dD��D�a��;�:s���Jm��I��0�q v�����?��YIq���r��L\&����"�D*��d$e
�"��"m�ʙ�����h�7Y��+Y����I�e�����)���R�Ԣ�:p(q��<y��a�"���O��o{��5w4}gբ�D)�<�rHqޕ������� ���'+�Rt���2w�/����b<�����E�	��K;�&4d�shR�%������e�Ҕ��l�n�V�N�oKp%0�Bd��k���j��Y�?~���w6w�o�"�#�-5;e�t��m��{��Z�^��"�M�(�f=�N��חX�Jڪ�I��$p@�L
���蘘,,2��ВY�L<m��K�ű�K�G�eQ�7"������BL��/�����g�LV�0��LT�-5���:�=C��C��Uy��X��/��7�t�ܹ#i����,(%�����2 Q���i(z�4,�s1QעV���.���N��ļh����<}bf��N� ��ʥM԰���I��2�2�pi�bb�E�}�J�K�p������ 6�7#|�"A�gb���#R�G+�4̘a�a��/��:�w����3�#�MY�_X��b�`�>�5Aڲ��G˿ܶ�=�#d��H�8��sCs@�J�1��q���Z���_�>���?�3[�^9���:nZ������(3Yd��s-��^V�b��t}�Z��V��%+n�Mg�g�q*���O�`U鬵��Y4\�l��/���I?�E�9K�ci��2o�/�0��k�c�	�E\T7n��c!-��M� @�����`r���y���Ӎ7Y�C,+(���Q�־\m�$6]�_�q	e���	f8v����N�:�[�x�P��d������'�(̶͒�O.|�!�2��������U��+.�T�z���2(�w� ��7
a^���0�{����pD+�K<��H2&ٌ��|c&�v�,�:�CRs@6���j���]xg����!W�*V9}f�b�hTB}���܍���Aa�h�V�p��E�'y�d����;A!�>��Ӷ�	�Y��j�Oit��1�!ۡ\>XV�Q2�I7�H�����E2$�p����5X�ڸ��+3.H���{�:ZV;N��f+��M�Ǝֈ0�<U+u�w�-��2��R��r�Z�!U%��㳳�&������5@�N�ꢕ&M
����V�w��1)�,N@BH����4m��M�lP���I�5Ӭ�&~qw�HHJ�	�YN�rnnU9
�����G����
��!�>�k��
ˉ�*�[��^�o��oyb ���E<��I@	T17�ՠd�84e�k���R�D�j�k_͖n��ӯ���Y&�LI�:.��	�R�D��u��ۥ�f�%�������srE�_�T�����MȈ礙����J�bD\��(��=�U�b9}���|�����[��Z|����ŜF����|����;�k0O�ΰ~�c�g�M\ɭ�:�H��k�ޏ~�E��ŋ�9GrB���˹`�^z�弴�@��{���=��Q�!��{y�Q��<!��q�7 Ǯ�)&��1��-[�^`V���e�~�c����/��� G��@�鷺��#�����J)W6�I
�Tr�������	�O|�~�� K�v Ѕ�T�kw�mgM�7�����F�n�n�#*��?�xP��+W)Jv_�-7��S-0�9�(g�y�-ls[6oqs�����S@-9_�a�4��ɩ3�OJV�ĩB��	��~�y��z�U��<}����ŵӲ�Qxn�Rks��R�c%ڊW馥��&��W�X8����� \PJZ��/�Z.U����n�جs�hGԫ$v��,��6�ܩ�� �,D&*[�P�9ݒ�x@�l�,
�y7�	��M(�ÓT,�|�l����	��)T ��^�N�<u���<߁*���e�$׊�����zrr����{�ɧ̌H�Q�M���؅��㸴��t�Y�RwA���
��s hqCQY�gY{(yS�0�U����Sk)�4ԛ��Ϟpo��fe �����, !6X���T1�l�4�P�Ky+c�b�n��k��� 0Y#���e�w�#�~��m�-	�����Zb��'u�hM��I�� Y�i���{�u˦�L`\�#��C���k��f�f�_��2��D��q��<C+���9�2�{'�[Jh�*�O�e�Y�)����p��{���lNV/ˬ�3��4�[Zq�"Q�bX'��4�C1�g���4@��Z	���=#2�ܹ3����W�^�1"�R�ZM��ѵ���`6�Y��]9�(ج$�c)����+�&^�_�;�g�d�1?��w���� j�	(u�? �9*~#?�+�j�ͤĩ<��-*-�4�Io�t"�q��'�I�Q,�hl������p �l@U�h{�GB^�7�=����䉓�x/���=�1���-���9�}�5�ݶ��e��y�\�+k�����-�lټٝ>{�H�!����~�B1w����ȭ4bpKE��>%���_P��T���4�(n�b�����6!l%1Y�A�_+u����^JC�mr�Y�y������  �E�9j)��w�B2�4�B�<&LbY�d��y,0�L~�L̵�Ry?\ X} %l�zN	\=K��6������\W��
�!d�Z��z�IK�������3}b�t�Z�YR�.���E��"���{k|X�$�<�ǈ �,�S�/Y��N��x�*���g��(F�`�(K��c�������<;��{=���9����ll����*���e.Jg���s��\��?O�F���.�|	�9�6�G�+ F�+����=����������ZD�¶'\X����
ի/*�4K���A��ep�rD��ϓ�%��匛�WaU��B��&026j�
���b�I6H�ѐ��p��И�or��G�J������ ��?�l�:=����%��]�)��z"�)A�:e\�g���3����#�n�X�T\�����s9^���Zp��(H9њV?�L���˳[A�M���;v�{��MI�%�q���={��$�\���Y����d�*�Ü�p���&0�����ܰo�|�A� ��Z󗒔��+�U�[(PH17`=D7��?GbQѣG��W�l��y2�G,���-d�SC�����}=08bJj �g�w�!����ts�
^�;���,u��`�V!�C@5sg']���r�%r.���ZmU95��c�, Lj68��1���� ӄ��M_*�~|m�9?&�R\Ĵ����R��%_j��A�����"��LlR|�ZR�S|�|�k1�#@J�8�ι��uot<0�  �J������ '�D�̜ς�?YH�m��+2 �	Nv�_|�]��4�����F�Θ�&��,�q�� ��`6!<��*lz�I@�C�������TXT�l�{Rr�`�	����v��1s��&�]���M��1��i
�g�{�=��syD��ud�2g�������1�/lЖ;)�(�I�\m`����[�\c)�7!悯���T�f�r��0�����dV�6#�V���['�k ��'�'�m>VwO��}�q��̲�]���~3^���������l��^�X|����]	"��ֿ���_~�E����n��u�K����*�u���:|�����^���{Oz���%H2�u�<�_s�:�[Q�����\Z�#��lce�"y%�y��9K�����kw]k��G�O�^k�����>P2�r`׮����w�O�?�48H���\�r� ��62m�_�J�B��J����Ĳ�F%Sr>u�3� �*Q�x/�nT�0
�Db1�!_,�n��x���O����[�O(	X@D�O��4J@�3+XV6�~MpO��[w�L��k˵�,��v#dQ�_w��$m����D�M��6�j�f�L6���N����A�{<z�`m��ۭȋʲJ��o��K���K�G6�ܟ�Σ��&a'�����\!XD}
���i��q���q�-�ڽ5b:\U�eUH�O'������)#N�������.� ��.�i&zG?�#Iw������e��5�G ȥc�߼��>��;����w>��m p�n����"��1T�C֙��y���9��<��)��}�JZ��$�k�܅`��a�,� ��N���*����+A��~4�;s�Y�к"�/���74e�"����Ģn��?qu^*�j�	�X\VE���i/�G%�{W�]��zY=�g���oޭ`	���.di.Ǆ`m�P�^������r:�*u��B��w��}�2��\�p>������4��R�sn��,�q+dSMy8|/�Z���l�[�&�l؏��/�W��!�������5P���S'��S'�2w��Qw��q����DCїd�%��ƚ� B�.i�0�:h�\�;nd*@B�x �7�\1q=o߾����kw{�.��lڴ���h�R(�lk�\���v�3�2o�学��Ĕ��zt� '��pwx �8'�#��c�!C|66ȡ�A̹f3D�7h#d��۳�l̥(�4'Ұv���I� �M:���,CV�-衯_�O�^5���{��~�D:ܕzCnxY�:�^�!n}a��mN�ޝ{��1����Q��h	��{�����D-싑�
(��d�(�xqKY�mL@k!ٶ&<�b-��,�-֒W"�=�x]Vv�j���ۻ;F5ڈs��5+�V�H���G,i� ����U�+gIr�K�-�9���7��"�-�P�7^/��]����H�I�n'�1�G�N������EC���QM�\�@�Z/`��SK�%��D((�c0��	 ����/�ȷ�>��%O��H0��`�	e &��sގE  J��^m����fn����aC�pt��*'��hZ^��i_�V�9�z�Ϲa�Ƽ�0�G�)Y�I&�qڐ��K Q�����ȉ!�<Ҭp�X�vP�&���q�̺�~����f,��m1��J�^�е�\J��&�Y�%���!�w����Қ�ض��~��߆����}��~�w�H���e����1�������'>�kH��mڲ�һ;q���_w_��tO?���!�L4��ZjsJ# ӵV�J@+�<C��M�]���˯߼�x�b� i<��s�o�� �M��3�V\�|I�J���r��d7�$�,�lc����Q>df����n�&S2KݐZxN�D�g�Ò����? 
���1d`Ğ�ˎ�N��-�丩�s�M��I��v^�����g�����xT� .H��Ϲ�5k�"1���7�.�?���92X�m2b�-�ܑQ����H~�3���i��s�Pe�,Ƹ�_|�� ��G�{0_��� kǏ���R�2/�]�۩ҩ�|�e��ܺ��\�y�α���ȧ�G�\&�Rm�|��S�N/i[mK��5	�i\ޭP���D �J��w�65[�!�&u�S�d1�*��V\�Y�/T���.�S�3�� ��QVq��ZqP�j�i�g�Z�pB��^EA����׏�e�d�n�u�Pz��.��v�*L��u��{����	835����'јȃ���*�evg2�0�}��\�6g��ɜ=s�,�?���;�0�ѳxx����'y��l ���^iiɷl�PO�X��`�z 
��]���Y�|?���^z�_琁+�u�J��Y�ɛ����0�^s�6K�W�Bu��S^X��{bh,���cG���܅�s��)�LQ��Hy���9ӄ4��R
��2�BM3��l�٩�yH�],�TʳY��k-�y�5 @�I ���;@�6V���v�)l�d��yA��k���[���U{�¤;��Q�����s�}�3��;���3@cF��7§������#���Y�Y�Ҡ1�(>���K���KrWY�i�]�Ew��̦�2EaF���X1�16�{ n�n���?IQY�/�M����l�j����T�ŰzZ�
DYY��r��4�;�f��:b�$��>k�a|5Z��6�!��M�����c�>�R�.an4�2�h�CFr$��'ܷ.<������LA"����d_H!A�r�ϲJ��������Ĥ���;,����u���Vh��x ������ܬ�eb9	U��Ұ��͇<$a�)2a����2�2}�"&�{���� ��9����x�EXF	l4붾hը`a�D�֨U�g�����X;�s}��O3�,�#PB�����4q�e�$��͇2	��a���
Q�E���Ԣ��6���r��K	�v�y��J��ي]Tr/�b��GO���tĊ�{�"s/GR� -������P4���HsX"�:��kYB5���B�4G#������9 
�`�L������,��Ù�^Sy�� �@[����eW��b)FM[J��n9.Ѱ�L-�gq�)�z�bg������,5�����Ѧ��LK�Y�5^���c��	pU2V1N�gҮL�+u�7�4
ʹ�Z%��)�6�b�'�V�[��޽�M�  �RO �B���9\�x�=�׹m�\�>���k,,7����Nw�6����z�k���-���>�������p�v���*�~۱s�mt;��0�+�u��"틫�M@.�:
Q�d�p0FZҨ{�y�ֵ�hQ�14�,7Ay
	5�����M���|�ݰw���pj��[��o�@��7���O=���Tg���9�H�ɛ�L�eY��5�"6� ��v
��"�����ۢ��g��5nzf2'淚w��Ixj�K$i������U��<ePA���5��U������f�Z��W�~j�z�	����?�=���n�����5�����k�u��ZRF��ϰ��܉�Gݹ��Q\{��4�~`�3�\��xN����,A���Z����
ht�\��$ �ʝ%�%�h�u�֭�����lJ�}���L+M�G�%�{����h�^�Xx� ��.�j�/+v�� �������E�֛�.��]y� Ϊ�	��˿�����z����K��#:U���8>�zl��g��;7��Nmi��[�$T�V�!�����Q}�1��	1���Ԍ��lҥ��� L�ݻ7_�)�&]\��)u��4i�Wd<�m���+�� �
.�
����E�n՝:}ֈh��m�9�ZΏi"�L�,v����������(�6=3kZ��t�ADX���>�.Ң���3R)���24\�����J(h� E?�t�f�����ٳǢ�f<���p	S$���/u����:3�q�qoT+���u��"�]j���t��P%#�+�a�z=<2fiX�o��m�A����P������O����_�/7=u��}��pC���θ�TT����}�q�Z&O���5�ן��qr�F��%�!���=�5
��Ƈ���]-/?y�����vך+�gڗ�gh�����k�81�F�ݮ���=��s����t��y���&�����0K��s�&ற�B@�<�l���_� k�\�"�[�0_� �O�d���'IVzр�����sSd�o���4˓��[��0�C;l��C5�o�r�X�����ϩѴ�s�-7�5=���JΙ#~���n)�:�kR�`}(�X�&/�?�$c���U�V�N����i�B��V;�[��ڭ����ԙ'
�O]�aTr`Ę(�*/ϐz 5霑��-��#�)�*׷"��R��Zq���<W�S�h����^\�m۶�+������E?-���$�i�z4���^M���pj�Z[���i��$9��h��=��(4����,{�I7���$�H0]�� ��KRA6M��AD�6G%�!���
��F�a2��f�~����nfiR1~1�B��B�9Јfc���C��0�[VݛBg��� ӱ-&B�=�@�-/VI����E���u��qL�k�f���v�F;W�噙 rʭ���R�� D�!L�O¿��"A�j���ͥS�T�iA�d���:���f5�rN�K�i���Zrn�c��M<,V�F�:t�=��)D����>���mx53���'���������=p�}�?w��e�u]	��x6�+�}��D)�iQ��%3=�^�<3k���h�ì�����"E��͖��!˪B��J��{�{���2+�J�}��2�e�0��{�>��#���u{��H�VΝ���_��%���,;pp?Q;&�Y�X�F�yB*"�qT�q�R�z�n(�b����E*��;�� �������6S�hVj�X[M�.囧�1����$�>i��Y��:5�����p��Z�M��w�Q�H�~�0kf��_�~,�0�G�7U�=ҹa�?�ӆ^	�h�ɻu�KR�ș�&�)4>44=�s1������rk|;j��ZFS��0W�ҽu����#{���t�g�9;�;{�(�-�������M.�]�����8��N_R�}6�a%hC��A�/D���؎ ��yc6k����X������1��0T}[s�έdWBe�iv$�t��1��rMI��9�~���a�:]~��������,-.��yj���U��v��Us<҆���Z���cT��ڗ��	�[M��?���l�����l����cSFyB�����37�ഀ|���/}��5p�82nދ��e��wȧ�G*(���
���o�6��^�iCv�Y�tx�����8G�jjj��k�Ev�IQ�}*�m�;�q�Ԇd���YW��.7�N9a�fu�� x3}�k ��
�i$SE����.����k-oR)7�[�R�\p�ۇUN6�u���y��-$m�݇��G�ؚ���ü�
6�1R��s��t+�jQXՃ�=�J�U�;�q���{���˓O<.����H�T�]�tE��%�:^��+r��M��o�W��&v��i�pP/m�M���$�w�T5(�֑w�y�kD%�"ߟ���Y%���ȹ�A�
�+�<�A�ߞ�F��h�G��r�"�p�>��6�UY"��mDʩ�%���sF��HJ��G��T�'(L9��+^��h&8&X#|_�U���R삀�AB�8&�.x%��#���ٻo7Ӄp`�=�Cn>Q��762����� wĽw�95G�p�ܹͬ=˾m#�5�]�)�t�ݗ����q7�g�D�Ԍ)mT��YI�P^�Y'�1���_���Q�
����bv�'�dQ�᭷����?�е3E�Q1��]Sc��D��y��1h�����J.�zQ�Ll&��?�8�v4shB�6���X�A1D������1%���w�>��{��&�G���E4j�����\� ���X��?��ȣ�y<�f�ݣ�����6�ɛo4`tl�^@�]�Q�6ܔ�3���m��y��g��aa���7�6�׶�v׹�i�3P�:|/�Z�ښ*���=sfcs,��%�&��F%���g�k�*ܤ����C�vN�s�{����a2�d�@r�3B�΂"�H���5H��)�^�u��2�������RPv�f�J�^eO>�QR�K/��\}ydJ�V��]ب���ӗ^���%3�����nxU��O�t�����?.��n�d�ep�fv�iw���X-Re�m·nݔ_��KVع#��5lL�t�F4iG(�B�s�}�w�
�A#4��C[I�*.�6����>�Mȧɐj�t�
S<CGFќ��xk��{�9�O{�v]4�Tŏ̩�v
$��"��Kȋ
S'��=�g#bM�'���D4�*lD�o�<��ٯ=�g�.��ezf�ܘz�����5� 1���6���E�Qe�����5)�O&귲���_s8�ť9��̳�a���U�*Y� ���_��s��`�|�h`R !��Hi�qfc��!P�r2P+0�n��]��W��2h ��!Mj)/����n�&7�Y�3�;���:D�`͑	)��Lbj�>��ye�jй��;���}(�sH5{.l2�+=���x$NM9��?�
�|C��h�oZ9R��2�ʟ�/{e�?��88���A��uQ+Z���ܹs�F�yԡ�1�L�#JF�����Dk�o�G����?�p�g&:��n�wHǆn���칹{�>B�)I\����6�;�6 ���ZB|�� "]U��S����,D�U�<��0Hk�]��a���)��독�i��J�wF�'6�Pr<4l�[����Т.+��¨�H$�k��!��is^6vޱw��!�	���Wo�I� U+Q�U7�Y��(�S���q Ҭ�۸?woߐ�?��{rgu��=H��D���={��qn�px!����.�<��{ݞ�f���������6��r��EV� �2>>B���}?n�pr]SP�FԎ�΂��_;�(�f�Ǡ�b�1͎���3�c�������̣�����'Y��
�a��L^�����J�8G��
����,�sV�yi+]O}�6�D�
;�H��qhdJ�;$���S'�ȱ�d�i�8�X>�|�LXz�*�S]OC�2�Q��,&Ǧ9�u�$jS��i�XLΌ2���{P����{L�5rf���r:4�����ӡI=���9��}&Dʄ_غ����H�b>Co�=�o���A�{�=hX���l8�j1�� �P89%�(p�kQ���ôw�O.�8�)�����dp|U��X'z)ju�����x�Ǝ*
��
��c��LO0�>+�F�(`��H�/���ǻ��e/D�W%�zJ��8Aª6�L�^F\3�4�82�R�B1���K�|3I��mۢ0��d�4�zJ��g���ά�\��I�n�s�����$s�n��G�f7�N���Ȱ4���`~Y�8�%�\��,�A�%����ϡ7�Y��NMAo!�pN��)�bc���SM]�>-Unk��S����qo`�L)�ѐM�cy{s��6�q�g�i!�i��ǎ��afe���p���p��u���s��S�����'7�=#�<��IY�;+�?�"�* �un�mх�(�r��r��� e�6P���M~��V�2�ÑC�d��)[X�&��W�ni����s����z������Z�6��:$��{f�|�s���'��æ�6��gA��
0"���a�[2�8/�˺D*p?��
�3�
$��_�H�>�7���G��z,�9�1�nO�t hK�Z�24�SϜ����q��9ٻo������s�tiu�*�G��W�Χ�e~��c ��7�4_pzZ)�QmΉ��*�?1	�����&���{,�G8���DZ��w.ڋ���wn�f��Z����d=��l/�����=�+�k�4��l���~�큍 J��������$����:�߱W�&���S(H�m��>?r~����k��*#���?h/)�s�H�;.�rA�O��FZ��r�3��gŖ�2q�D>�v��c����6[�a�oZ�ݍ���?]�����85a5���������O��<����1���&S���
A�<���"�4`�|nܺ)�/\`C<�u[��Y�6��U���y��9v���ٻG���%c��i6k��1�'�}ץ箓?��M ��c�ꜛ{�����Y�y�so��������l��T�ɝ�>`I��GVe4�4�1�i��>�]~�?�Q_�F�J����A�}��ޕ۷n)'#jz���61�e'w��\��G��'��.2�5�J0��{�s��Ͻ�9��L3*�s��۔k29����ҝk2Rs�;u�6눪�V�<����*�\�Clt��躍�1"��|J:."�[Z���0�#�/�%���t��o}ޝ�y~��6B��W��{IO��˸�|@Ɔs�]��w*��4��yP�w����f�<�;���*�F��ȈZ�9�iqE���Z�tj�� n�ϲ�q^!�9 �����xc ݂>Q���Ω��=��r��a0�.ʠ[��������
J� IՀU3H��a���yE�`��hɔ�u)����o�.(M��0p᪼����We�]����8Z���5E���G��Y	�v$/P8#���9ek8�(�(#����x�w�ܕ{w�@��3�j�5��
K��3�tq�Dk����mT�Q��"�����$���>����J'}�ʟ2QE��i8vD|�9�Rk�����_m��=8�E�G�2S��Bo�2B^Ȁ��qI08��FY�5��?���l��|�Q�X��f���B�H�9�`����z{�mjs259-'O��'�=.gΞ"ApttH�F.J�yG�]K]	��l����L?��4Um4G�gVcZa�3`��X^n����0���}�]�{g^*uq�����iAaPk�*7��u��r��1S���ʂ۽��������Zs����XZZd��믿F10hm�1��orBi���;��*���������5G_���15��c�q9}������Yn|���|��{&˲g�n�tlz�
�HW,�4e�ݛ�Z"�H܎���ͼJ�"�Ľ�r��THU��T��w��癩iՃ��&�OP��}��e���t{e����y��_pÛ�������ƙ"@?2(���-ڑ��W5��Vid�:�=N��{��a��<@0���UP��Q�'�ޡ�0�5�n�+��і H�bT�U_48u{d�@��Q6�%�T����S@]�ǇdffB&�����df�(˲%��L�I��82 ��y⟥����&D�
��b�#��Â�b� <8�	=�ؑ��]��ڥ$����w���ܳ|����WX)�gQQN^�xG2�A���t�!GJ�V��6m����@�i�;��򾱼Z@}R5]4���{��@!�h�A�ڔ�hߗ����5�]��f1M"C٬��a�es�<?�BU�|��R`��Ӣ-�P�Y���G�~�?O�1�o� ;:vĩ���]u����\��b���,����E��k�x�9D3~B�%��ª��}����G[�r*�}�95&��K��*����RK� ݓ�� x����Ľ����}Z:좺�4��f$��;\45l�گ&�����'�e��qʽ���/�j�H��=�Έ��/g;��9�sk^.~���;-��J�/,.�W���3(55��qK;���Xf���L]�p�D�@������edf9�幱��h�.nӽ����b�8#	3�$Obt�i������#�r��r\�@M�tjfJFn�С[^��n{�1NOM0��()E:���͑�$ޑ��TEi��qĞ|\ ��!k�Gn�t�J\s�:�Oʺs��i˝g���7��pm���޵+�*���@�r�JȇmY�G���9�sq:pݴ�L�HSxG�i��-4t������5����'.Q�OS3@e���n� �:�W����u����H�yԔ�c���\ﳃ�3���d�+5V�`�V\tШw	���5s츢�cC2�g\*��HOj�VB94%�4�5i���s*�Ty�����p��T9ߠU-�(-b�8W�RYWB"o�9��NEV�$���O��ĺ|�;H?������tM*A�O.J\���j�V5��<H�p �چ��-��n�æ���V����Q8�����-VV��i,�w{�l�c���Q�p��9/�`��T8�����M��$ 0���#<��\�Nh�<�6�c�8e^`��]O�X6��G1�S>��Ҳ�}o�6�"-`�2`;��ߠ�B���ܶ;
���&�3�&��B.G� ��Kym6�0b'|�h)##�؜���X�E��UN�V{�����agpG�g�����3O��k� oKk�����Iw|����e,��8"���D�"�XwSFIǉLL9C�뤜Z��ʕ[Rry�&�/]���e��;'�s�E�/67�����}��o\L����8#��Tt�7?O�742�64~kɘ�w%�Eg%�P+FeԱ#Ge�mW(���t�<�/*9�½���1�A�a�'���g�0���c���=9�N��x^���H��]E��0_������l$���qE7�X.s�_�a�ę�E^�<�qt;���λ�ܲ���HRSa8V�4jl��$�3��w\t}�����
#R,�v�ؠ�#$Z9,ݗ��� [�	�˻Ｃ��]�e6�4�;6y��m��l�+���8)kn�?��4ܑ�Ś�{�Jg#ͳ>���q�@:�*kj�q��|G	����F���Oɹ����f�/:��a~I<7"b(O1L8�V�s��!e�`uW�%�����Ы�5�衤�-� ,��q&�b/��#$��Vwn-\W&33���/}^{�ӊ?��+�x��	$��f��Hz��p
�
���3�{�� ����X�)e���ޱ)9|��<�ē219#��-�v��s�ޓ.]f��i���}{�Rx��vPwC^�1�þ���p�	�/~fS}�C�=w��te��Ϗ�rv�m����a�Zq^ǥ<����X��鲄�~n�|�{v;���n�y�kʓb3���rglN̓ޯ���ll6�KAm�t���d�dl�4�ݽǈ�n�d���Ϊ����#��5._�����G����2:�"�˾#z�����О?���ȭh)�
F�j%��X�LE��4�ԥ3(��������ߑ7�x�El���4�ؖ��%7�rv����^w����J���J���\PHq762��fN� �	��8B����ߣ4�a��?�u`���ꫬ��NK�5AhL3ꎘ蠂�;��������_|�r0?�2��D���\��1F�
a�{wn��5>B�&��\��E��^��E�!��!��bn��}r�;Cp�2d�-���]���U�������رc26:^�Ě�R��~���m68�|_;I��#�W+\��fU���q^�Q��L�$���#��>y��aVT.)�r��M��������!���U�uٷo�:�_>���e|�鎽FG�טZ���i5�ۙ�7��K�sr�YA�b��`SX1��DU<tm��'��ךo�2�kE��i7�ݼ�y�sL[:{���c���3E����n�o3����n�uǐ�uE�Y�HA��(kya�3���B5_��޻grR~��������ĉ�$C��[;G��)���ȹ��6���^�ӊ5��f���8Ap��l�#��И
����0[m����9��`5�(
�GI��:���矐���&$܅��<&�[���TH�,z�}�@���ѝ�V��m������'�a#���ZY[����:'搜:}�E��K���*�ٿ�"mNT�o���P����-�`�l�i��3�f�~W��2=="_��g������o���-�����=�e����Ù������?p2�wM1���e�v�1�4�!���n$SG�ȓO>!?��,ux�Ϲ7{WF����߁�e����V�}O�
�;k�i,�S���`sU�Ƞz	�Z��N X�cmbsE�$�&&�����jSI�M8��6�zC%�+�â@�Z7ʥ��=��l1R^&�c���#�+|���á��'�9��7�l��k�<�3����IˇF�8_���
�t�}����<h���p��a��<�s��u�i��LE$yA�עmt&��c�s�{�E���y��3r���=6o��3�#�󪦛�~���$ռ�=�\�U�~67v�δ�����G�p���%�aJ�N7H\zIu�ω���-뷕�TV�t���$�̝M��`�cS���~_���&�������-	�����^���2�Þ�7�<J��yq]8IΡ8v�|��_��h4�)�q���3O?#W�^��i� l46�%Ԑ�ln���X#�NԦ1l^:-��V-:�4yO^e;{T߾�+t׳�s���>!�#�#aXyr��Ҁ^Ė�Y�F�a��P<,Gg��D�{{�ޚ����F�}4�l?+�v��qs���5a�2Zg��޽)G�tQ�s��/�(�O��zg�'=��B�b�B�����"i�%�J�}Cf� �	6�J����x�^?�^�s��q�o��slޓ�{+���L>6�u笽�W,O*u���} U��8y�۸��ݷ��ϑ���=�ksN�yV�59��!����r���c� ��'��J�T��*H�EsRg�����	4j�9x�2���*�3�4��)(��6�&R�H<�jd� GI?ȇ��J�w�q���!������Jt/�Bf�U�r?�-�y�=:,M��ˮ=,ɶM�ܣ��F��q8/&�O�O��6���fk5���FlH�Q�N�Fh�t�nŹ���F�e%v+��f���+���wO��_N�:*�>�K����M�+ޚ�#��5�;�ڿ*�0��T5sf]�3��,���vr��p�5�!��Q����2�W�@ҩ�c���Vg���7��{;c��uw���b�����7��}�=�~��/�|�U�l ��tiŗf��D���b?��P4-�V��S�?p�< SSl'���)�a�FF�����Ct)�(=1<���Ͳ�cu�<������qj�ug8��BcU�&/R���[EiB�2|S8���H5εq�?��H��D�A9�P��"$]�Q�Zk�?�)�O����oT���
*�����G��Q��o��.��>EZ]Tq��|��{��$�M
^@W�z�q�����<��Ӳg�4]�����(M��Ѝ(�)jr,���Q��A�;B�35�:���F���0��`lg�w��u���W�]������:K22>$�a-S^^[&���s��I����^OH@�A�3���T̵I�CW�N�R1�|IN�9C���Ī��K������c @��[ٺ?�[�/_&��s ����L�$��+���0�P8�j�^��:J�[��FƟ��P�t������6�&N�d�$ֹ�D��\�{�
��߻�%��n��7�����}�63�&�Xv.�M�y�L�@�t0/�6������w��%C�U�k�����Fg� a��+����>rHN�:�
��G������^%7G��
�R�HSt�m�̊�$��w�XTap���v�y�k�^u��jK��W����lԛ��|�m�y���]:k�Ч�Z��<���[C$�� }k��F��-y>�j��^E��)i�2#����gezf���+?��,..w��\ӛln��Q!ʈ�"PT��{6p�������{ #3'8��߳s����r�k4�<4�.�Q7�76B��el'����g���t�hd谥�~�f3�;܏Y t�;K��q�`�L�uIi��9�1�=Ck�_C�Tz�Q ?S�-��y�5LG�95�' n�3����S����<���C3H,4���k��Z=���9&���3ȝ���!9v��ɟ~C~�7�v���%���FI=�K7gC��C\�*����M�Q\��̹�X�'��(��5��噽��L'��8�F��zW���]qFw�ݓ1�V��*���Q��Fz�.�p_���>��G端��8�ð�v�.7Z8��n��e����7V���G��ܧi�Q3��擑��4�C$�_��(�D�ÒQ��L5Jpy0����Ħ��7TN?X_t���t����ٗ�Jק5=�#E@b`/LC&�6;WC����v��G�Є�)�=eG� �o�n0w��Vʺ^]=�W2.����0�f��Иٷw�shN������5-{�L�9�t���4>�\+�=��)�+D�3�� ��%w������8�$��D����t���A*-c1���*E81Zk�L���AM�-��u�Rp�:/�FI�Gzxf��FQ�,䲩��j)���q��9'�����іR�+���W�dl���)��"�߰���1�[�p�����A��o��?��ŁC��̠����w���>c �ι�� ��e���ɞ�!�Ɨ)�!P5���!2d�Ҳe�f�S?�{���{�c�畨��������)49�A�P��D_��@�ǋ��6C0
,�QxO��vxbPbjlx���D_$�*ة���]�V���tB�V�S�:�>�Q!�Ni�q���QY�1�<��9����sy��s����e�ڢ�4�E����>�mF�(�Pb)n����4��+���(Q�.���Ѿ=F��=	�M��ǁ��	У�����w���_���a��^r�ˢ�NL�n��iMq�tƾ�C��*�>@�p��+�y�,-�05::��Xw/ )��.�ko�#.^fi�=C8T����u
�Y:n���� ��P7$�!���+�jp�$M��7�"q�)�k�������6��dG��V7Y� �@Q�����p�( ��&�~�jj�X�|�����.��u�Y"�	*���ks���XT[6�9#�G���c0M@�m� ��H"�A�ō�W��Ga�'���@�x��I9qꘛ�1�\����9�P%�{(���Ԉ����R�V���������sh���_X&B��:t�-;�� "���ngQVW��*5��1lp�M�PU���!��&��έ�{kU�����#c295*Q3fe+������x%��d�<��?��ߗ7����Z1�(�x1�R�|X�SǳG�:7"e�����p��U�u���[��6�^���ݿ�9Q��+��_�W
t�3�W8YO>�$�,!��C��P=4%�rC������L1���CN�6u���H$,�i�� ���2|��d��7��;F�S�$E�5p3�(���r�lt���������0'&�����&;�(
��-���6�AƲ�kz$�?�KLX�}(D���b��é��ߺ}�����W����r��Sn�/���(�)�fj� %f��e7������K�}z�P$g��JH��l���m@��sק����pE��#_^��?�+U�0Y��ԝ|�3�dbzB����\�z���*��{c�l-�{57����w�*��*F�)��oذ��]�rE~�����*U8M	�i�q~Rc����	���t¼�n��N�b�c�#�F�L�����kf��Ǯנ@Z��*��U��3�l����oЦZ�s�9��[�Mn��a�ҫYYY%��Db6��ѡ4�k�� (�X���ЌO��f�q����}�9�"z��H\�55a�e)
4�ܻo�&��3�<'�����|��kM��lM�>Wl�M��,��t�j-�ض$�8�Ҕ��6N��^K�s�ž��9�ܤ��.+:�3;�kZY���Rg��W�#Ֆv�B�t�^p��D����h�}߯�E}�LT���ɣ�G�o�#2"����t�;^az6H�5�b�E�y��Z���r��r%f�����]��+�Hchԝo�O����L+	��{a�]�kz9h�h|�*��b�	�
tɚ c��f�̓� .^qn�Yz�#�x���z���h�#���g�P4,�����Iy����������wb�)RO���$�l��s�8v(�0(�n/F�qr�6�u�5t���x���2!�b���/��?�ӧO�({YU?#�x��ا2/|%�	�-[��qY�ɲ��Ŧ|v9��Ry�B�MAu�B�$�"7K݋\	ɚ��95���;I��\��E�t�*�����?q�}fS~�ßȕ�����e��j�\�z��_���������%A�ސ���KK@b�p^�(���LQ�D�8HW�_��mg�|�� ��$F��(D���y��wɣA[42��g?K��o�Rjͺ<q�qj��n���&�D:�42C��Zd^����%F�uG,u�g�y ����;$��27;���1��G�"M�׌�k�R�|�#������o��k�N�q>����^
�G�e�d�6heI49��$z�9��<����.������ge����}�#��{�S�K}��$�N7f�h~�#K]:8�����>H�4}��C
��Wh%�}½�MB�hj*�trǭ����Q��;��Fܦ��C�dt�NN\��{�qt~�|�ˏ?"_��o�p�ʏB�s(`��k��K��(*��hqM*��w?��*+HeVjDoܸ%Qr����R�ԐJKc���/I�'��ɛN�Fs.���9�aY7'�X��� �[�i#�W����!	���<x���$:o<��������z5;���"4UL\44. ZO����
SP��9*$.形���� r� �f�[oNO�s(t�>��h��6�{�Դ[*60pFVﭐL�o�������s�GsJH���(L�)B#T�Dp��1��j,Ţ]r�YYʙFl,��N
�E܅ʰ{���*Җ�r�FDp��w�<,��yђNDt���4�4�=+p��G����*r��!]�f_�s�aV���qw~���� /�#4�S7j���v	Hvh�;�cs�V�T3]XXt�k�4��_�9�b��C`����';��{�w�S����"��ԩS����j�i}e�����>��H��ҹ$ϒޖ�X,m�
�(7�
E#��2��t��V�3I]��I;��Z����w��q�� ���ޑ�_~Y.\�������L<�4ب��"6���6�-?����K��C$b�J���Lm&��?���D.Q�}��~9y�4�U�k �`^k�kU��asN]��幺�q��"���g�1y6 p�(�C��H���#%�g�q�1������b,�$ͯ(B�̀�8�����|�96� E�^��@�!׎�$=�fDUN�>��o���m笯���z���������d|,8�$ӣ5�ۧ��[p�C�q�� ���4ih���2?�q������>X7$H����&A��|�2���i7U��V�>M�������W�M�N&���"iQ��e���0^A��F�D(�U�Vب�r8b׆]hCX�0\Rb7�N ߗ*sh
$�a�M��FD�4�-B3�jdcB��~��6��O<&���?��������ύ��:�-���~��ܻ�ʣ4�wE�J���M��Q煹j�e�!�T�C�H!_.*b�&)�x~�\&�oWz9s�xH�ڔT���k��h�N�b�Q��n�>�gy��U��"?TW�k����иa�ñ���Fq-��v��K�+uƵ�6�3{���\����l�Ps�Z��f�׉m�|V~�N>^M��Pi]._�ĞH����K�]81����{�	9|�0���r��]�}��{$ʹ/K�nR�89E��@���O�ƣo*�3ѵ�y�u��b���4xiwE�M09p�v�����-�E��1��g�7~���pb�!�	���.\'^nƙ��QZ`+�[Ao���Z�����S��2��y�-O%w(hZ���~<����g������r�����AA�����h�TT�&�����n��hM�T�.�
�!�Dt�RW��U�_:$��Ϯ��R��w6<Ǯ�4Cr+� ��zC�l�|^�����%��T����A0ҹ�0�	 ��}&6X���˱��z�����o�����IFsЇ��rQ���+z��u�i���pA�[(�9���sO��o9�iy�ه�~�vD�{�`3g8>����(	x�|Ur�<P������T��s#DG�o/!�C�@U���~��G���0�#Ej������c⫕Y�P��l�y?��J�eܗ������ O�x_�%Oy�Qރ8B��G _��cX��{���64��=�QI��DUi��r��1��W� ���g��bKl>hZ��*Gި�W,��e�����	}O�����t�d�[W�.F�H���}_)Ӵɼ��PJ�t�lmH�MɄ����+��FQ��~Yv��9�"@\h�j�{>2R�3g�K�%�E"3k+��pg����W�l���+O �OOO��NLMK��e��"� ~M=����83��Q>� �8LU6��NVBhn׮]�]31A���Q��J�E�o���\�x��$lD�ڽ�7����E���A�u�r�F�q�X�qF��#��e�WP���_��΢��c����i����V���D�P^|��MV�=vX�������{����/�/��g����\����9��SU!Y�|��x0D���	߃Qv���VL9�.�g��y���/�j��O�'����3�o�n�3{���#�����qV�Ũrʕh�r	�(�|����X�ծ{��h�h�&����JMSF��@,�6m
ȼ�᳖;W�Yf��5��V�N���
�`\�Z�T���6�t~��|[�Ֆ4�C��T�.� TǾT�83��*I�HG�vN�g^xQn޸#Ks+n^�;�Ƌ�_�	��<��U��RC�x|bR8Ȋ�5�V�q����E�	@&���~���7qf��1�MUx�|����F�6ΧRt�����	L���UT�?��r�X�����.��{���^�; ;�u6!�~?�}!:g|������>M+�ʯU�����{��g����9��3� QT\h�R�_ ����˘o֎�0lP��l\�r�\{�E}n�ȯz'������n�0�@y:l�1/8/U��M��D.��{	��6����Hi��`E�l2�\;��{+�</w�Qq�Z��f�=p~�"|#Z�E��2��� ���7ȱֵ��i�[�)����� �{��a�q�[&\�~�N��\��Q=8��+˲���ݶܾu�ݛ{2ToJ�=���9�8���vΩ��&�Jӳx�/�zi��ml��2�M�.�ɜsj���笵x�M�Ӵ�~���舩X^[9�:��̠˼s���z�*7��7�v�{���H�<�M <F!Q0�a�3�i��8t����V6v2m$
ߙ�Ɵ{�i���%YZY��G��}{��6T��Hڹ	f�\w،�g��^�����e�4�Y�fБz4�����V�f���>��@@]��uB�h�����ny�^k��QLhi��hg�n$��EI;H��K.�^s�wS�D?|?�R�:7����k��򥧟b����w��lʚ��`F�-���W������V�H�_�V ���	�ף�<��a>yrh�ڼO��٠3�c"9�c�95!��X��,���	㉁�s�(=��>�A#��ߛ��pf���d��������]����b�/���a�}�)g𞑩�I_r[S]�v�;)�Ѻ61͔놣=�b?�+��N�>/���(��' {�o�i�?v�ze�pVi��T�ũ�au��J�R��!萠1]���"Yq�B�3�#J��oU�mw|l��]4�Ziݫ�O�,o�M����ciQ�G8چ0��@4
�	#����>ϭ�C�0��qR
���
/�ћo�R����� CZ�ѵ5�Ⱥ��՟�F�
� %���rK�{�8wG�nK��c81�7��xNGEK�)����+6ָ6/����L�H��Ϛ������/w��!ܽ����Mxz=	t�F���ɢ�3Rgx��|)6�^�~�����g��僞��hs^ 5V݂Ʃ��<y�	�1W��F�s�n�t�g�7	և�8Q��=e���:ǡ��`B9cQ3�Ϳ1���j7��ժ1��؈�Z�86�M�-�<P�qv
�u���@Z��M�b 
�P��CQ� �N )��}�FF�lw�ק�_qo}7Z�TW����e9��;���[�[�w�Ԥ��)�R 1��(L�h�z�ݢ��F�s��\ ��k��y��#xGY����Q���y��L����H6y������G~�-�g*��P/��:�gl���Tl5E��a9̍����s䏒^(C�V��i����++�D�>��i�*�i֑'�|\�~�i9r��w�J�v��@N��k.6�ſ�8�TyLoQ�8�>��&�ڎ�Po�T���A�5҂Q%/RZ� �KR[���H���[Q�F�"J��}!���5��!���4��}��v�=-g`���H�ԩӼ��(��'�SC�H$^_/������	g�� �9�SP����?��"������*�w�&ڦ-��KF�"��?�ͬ�`E�޺~Mf��v{]W*��S��6T͙X�C�TMY�@�������.���k2���U�F8R(?�fx��9������� �Z��ڞ��$��c؋�:���2诅yc$�2�ϞÃ����5c�Q�ĉ�r��)j.� -�g����&�;�n�Q|ő�5���)��DS֜ӏ��4]r�B�%ӕzBn��zB;��?�����*�U��7�u-.����0WWT���-�{2�&��B���D+7���髈���[_W5�؝�w�G��U�ћ�ܷ؝�[Z�t��3��o9ǄUA�b�(m�]�M�ٞ�9��/i[�%��p��Z-�4}���<�a�x�g66��|�a�ocr R��c�8�8t��N69����e�KG��RѰ2aP��F��}T��F��h���W�?��F�����jc�����f����������cGQ��y�t2ODc�&�L��	��P��ȷ	���|[����U�:�3��Q���C�t@#�t���O�N�{�f"qn��.����yBU.�w����%�"��x�:�G,Wg0�Qh�&�dv�Br��:�U48�g�����+�aJ
��A��ݩE��@!������HF���ay睷�+�F��K �$1����n�����A�	�S�$�n�E�]�;��9�rJ�GT�&����G�1��̅��|xkV�������Lm����a����S��V�E�)�剴%�i<mdස�rL��y�F�9P�Ч&B�ͭm<tv�R3R3�>fff䩧αS���2���q��4U����AI��\�>*V< �u����i�=�v��b�����P���G�}rk��N_���0o�m ����*����*�װ�Յqo��@(�*K���uU�؈mQa�ZOem�C�֬z{�'�_����i?6|�zkQ��ߧ�A�3��
���i��h��N�u�f���qP$�><dT6<�V�8m�f�ӥ�ЉO�UDE"5��0���kU�j�Wqjn��U;�scd,l�&6�����yh��(zd^w9w^���,mg�>�y����BQs�ۉSG�F5�6#���麶���
�J���jK;�N�M��,�mg��R6�C�:�n�j��G�Vu��T�56aw`t�F�U7���9?���T��x�C�HN��.űv�N�\*� ��D_z�g٩a5D�Θ潕C g�>�~X'\'yrjr��f@�G�a��ʕ+�@��o���QI��t�x�"w��F�8�z���@Y�[o�E����z�ݏ�r��U:;���b�E�U���0�shvv�Ɲ�� �v�!���R�	�+-CX���g�)���|鲴��Yz�>���5�\w��9~��LNM���jq���4@�׀�	������ꫯ]��Ӈ�:{P Tn��~�X�� �)�ϡ-�=�Q�; 1p�'��fש�ǯIr��ب4���9v���Cg�7J��g�`}Z�P�8� ����k25=)S3��mxm��i�4�x�ͯAO�F�xFۃ4r���ކsnF�Qf>���vdeE$��5φ�iԑ
ФX�0�dlK�N��#b�Z�_�S�"�pې~���<��7��;��p��vؒ 
쀭���XE���JIخ�R��9�0Fx��w�{fym�����h�E�A���r/����ǎ$�l���axͅ���ۉ�v��#��itQA�>EW������w؟���.������z���Q�x8u��Z�,�(N��H���p�f��]d�:VW��0-"�Y@vL��"��NxZ��l?RC�+�b���,!��(�7�I��_G�h�I���c�祯�2�"HH���Qu����0K��/1��d�:-Ha@��N��M��|���w��qG��" ��;ߑcǎ�Z!���ŋ�������j�Ь�|Y�=?p�3V�&�ڲ����"~�Mh|@�]I����<#���4����m�AUT�l"��/%/ݺ�!�\nQC*��Yd���7�7���B���3��<��Î��;�����ɺ+W��W�Xv�B4�"U�E
�	)��g�2����8��'�GdxdX�g�8���Y��Q5z
u�xH����f���њL�t�1��î�Ze[l��>u�JEϕҞoZ�H�'N%��2�'��v~H�2u�9�r��nYY\��W�ʝ;s��OȄ�)��1wU]\C"Mkk��*��=�.����AcAєs�>�ϐn�PB$���j͖-@E�͉��˯��'6g��yd�I,�����10q�lRDQO�(d��7n���,
'`�����iex<X�) ��cb�!���fj�����ݻ�-�	6���c��J���+	��]��0�S�Ϝ(��zm�˵�s!��N�3(]��Y=��8G��{�� �_|�H�K⌚4��G*���@�Z^���|5�=�F<O@z�Ah�#�_wm�sۻo�e��?�-+.���X�p-�Ďә.ޖϙ�cdL+n:[�}?M�|��\����?�<���W^�y�8KB5Դ;�f�����V
O?���Թ��t_�t���5w//�{|�E�k+K�{�Z�scbt��{HC<�W�="7�]��s�<�.�Kը&S��|��'d||B~�ӗ����㿳"i��^z��N�r�[޼�6#t��1!
~�c�4x0-��"Z��o��9�J�pW	�k�5"T��:t����ML���(�D1�.�w���}�).�K�r
�6@� �m�Pˆ�.Q���:4C#5-���{0yDTۖ��.�9����i�[Eb���O��RF!@��#Ք�GO���"�g.�?��|����v�ǣ���N4*���9�h�edlD�޼'+s��}�<A��f�}��s����/����<�[ٟ>�^�q��)4�k �;�p��M���
���ｏ�M��J_D�a����H����$��iFl>��.�U�r>��k�i+�8�>,�N�"�0��lP����+����<�!�F4�N��r�R��j9 ޱ��ؿ�B*{�d]��Y�ZH/1��i}<)�5%��h,����H��&� �nP��ɰc�{{ԼkX	�i�P1b�%�i�{���UB�TH~#��{��)��/j�p�[����"�r���(�3X(�����{:@9�7M�w��o`Xט#��;x`�|�+_�/����>��x�y��Y�C�޻+W._����_���T�(h�|~zfJ����Ǟ��{wˏ_��|�[���P��8<C)q����f=ĐJ�t�ɮ؀�1�I�
���9��)�y�!{fi�뺼�6N��0�ᜎ�G���SgX,���0�<�ow�Z�=_s׮����y�BE봤[,M��C�)"�=@~��Gݿ���Xbf��H���[��:6\�l�h�8��:�q�s�ϊ������Y��FE&�q:�@�VV;.���`�A�v��}`k�:���@��T{����S7.���c�xWpj�~��b?
�Yy~�Sm6��>�:�6�_���8ޣ�?�3��)�l]s�fC�Ԋ6>I�F��ؑ�S��muK��� q�R�A�se�Vx�A��i���Sk�z�,�/�A����-�9�=�v�$<2<L�G���F
���r���"���+�j�`����¯4z��'Y����K�A��=�N�ώص٧<D�C�#���<��)E�N�'�K�Sch����4X�)�F"�����dH�k�\�q��CDq� `���+$7*�(P#}�SS�V|Z��p�,a���b�cj�6%a����<�jI����������<*�v2��j(�j��ޥ�3��K�/����������>uJ�K���r���K����RXғ7���88<��tR �1� h��Q�T~���:��#�Y�����~�,�Ovs������z�8y�(RR�> ����S-��R��̿R�0��r��
�k�9��^��G��&:tb*,0�@��yi�k,ʍ���G��& &%�cj�#��;�Z�s~A��V�Y�c�Ω�|��'[�Ug����IJ�y�ʺ��\�^&v6�c#T^�_�9ñ��4ge��*�cf���^b�{�R��>�܉�������Ge��XL��NS��<�`'����I���jX�l3Tpj�� ��<�� ���a3	ǃ&�����^�r�	��������Ȣ�_�j�ˁ���R�UO����&]_86b�oՈ �ƽ�i�fL跎�5�G���t:|�u�t�oJ����K���ywCl��̞ED>�$��lE�(k4��Bo/��,	��[Y�zqW��z�A"k����E��Fp���c�Wsȭ)���ӯ��@[��yfcU&�Z��g�yV���`#Epa��YXX��>C��rN#�/��V�����?3=�{�.y湧�ĩc$pg�ܗ�C�)aԆ�dHZ���5cA�Fe�e���g�����~n�6�
�ϸצ��bx/�N�Ds�V1�F��L�O������j��aYZ�����C�I�/�"_u�Q�I��2U��,U�|�3rN�����9Urf�EC��@	p|�����1��e5�:WE�h�H���g�\�ᅣC�}���*�����Ep͊[�p�ZRk��*��pm����+�� ���6_E�N���-�v�%>,7o�"�ʸ2�}J��(�2��)�-����e�|>��[�}����o��x�k�g< m��&Z�6�c�s��{����1E�p�����/�=stA�K����'+�L�A"Be�nп��A��Q��>�6Q�lh��5�؊@+��s���۰a������V^�Է�~J$��y��z�M�:��T�U��o� ��f��D%I`|�H=���5��埗���J��Rn_�U�ް��z��i�L�+�Li�
+��Te��1?�*��K��!F�6��5:d6V��(W����z����Ӝ����/�ҡ]�W;�ZH��?�?r��i�i<h�|���e
�r������~K�y�ٵk��<uV�9!��śr���{��iwھT���Bf�B�6z
� זQݲ Y����7{��n��)���m9z7��6M��
��������-.�Ȫs�'&&��VΩIX[����Rn6�,��ԙ�D���+V�*�'����o��/��0I�k�#PI�Lk�x��l��<�'&�d���GE�y��
��xd����@&!?�����cwr�D�+�h!U�]�덈b�@g����2JQ"m�W,˘.�*1簹D��+�r��q�p��~�4�5�W<B��4�I�w{��4қDo}pΝ�Q��|
L�ò�f���0ȩ�p�fÊ�ŏY	[�`YG[�T���D�|����[	ky���Ӹ�ا;|��53��͈y�F��eCg?�h#��6'sR�Sl�͆�R���<ꥴU���Qb��-0�
FG��b�p���3�k�|�%�!j��+it�����J�B�	I�$��a@�vW����#%�����!
㋇�q��ľSw�7���o#�X��R .�1�'@hʩ[s�2+=Q�\��@�`Y��r������9Fs�x��
��z���r�=�3:6F.�R@�\][���~W���o�׷h�5���a# �����r��eY\\�Nɍ�י�B92�d�X樄�J��η3����4ct���������ő
�RkCgBGIov��-�dqi�m��d���222D[p��5��:ʸ=)�7�P�&#�X?�*�
��sr Q�DL7!���VsS�Ƶ���*ڧ�Ӌ�ܨ��0��s�)�H�,����U+�P+�P~�MƊ���32g�o�ʌ��N����;4��KO�v�3��=B �0Ҙ��C�Ĺ'�C9�q�T]S{xѝ+P��ڇ�5���@0���8m���-¿3C��,� 6�����G��?/��P�&�K���(Lo�ײY�P��@�����io46�6�K��$8:�ѶVX,m��a�n������ԙ3���3233��&��Q<<��^Q����)�]9�Vc]h=T	Mǀӡ+�"%Q�]�֜Փ���D�7:o'I��8��{`pz^�������K?�-b���ֿ��(�.6�ơ���*�c�2+*J)���a�^ՙTΉ���::6�qA���0G�!�hsF��r��V�����,z�`m/�*�?��ׯ����,����${���;�����euy�m.O�y�MW�o�kK� �6�е��Y��R��[Ȼ)�>v��A�2e)����)N�S,{N Jֱ���Q��� r�򰒫�0@����I^�k��4�F�5^�+>�-l��`p���!"�\�q��m�gY��7���qI����Rb��C��������5T�P"νV���cJ;r��Oi�i����z����^t#Dh�^���3�A����3�����\�zE�f�"����e:���-��vbl�(���"��ocH�VF�o�=(��-���RQڳ�G�,��t���qj��F?�R�vǎ5�S*��a�|8mi��1�Jz�9E�}���d2= ���!X����+	�_F��ѣT/���1.b)��3D��s�
�F�������$�2��AK���]�Ԭ�����JY2eI��K��c���E���k��v�fG�&,���-\���_@�� M�<=ˆ����\��:CDv��8�K�C�n����l��y�떆�
�ۘ���8إ!s.�ͥK���ŋ��9ϰۑ�ɭ۷����{j$B%��)��/�LNϙ�κ�De�:I����c�S����������,i^�`��qY��T���s���e�Z��cs78<Ҡ(�Gc�ju�s����]���f��K���OP��^i	�������s���vQͅ�Y�!r��D��[�a����8�D�'�zN>��3S]��u�%u��=�b��qʼ&rx���r�dZjK����V�v�J�U�1��G���O�Z'2�k����w�#/&	�Ju��Bݽ�*zkvb;N�f���c�����e�{���=:�r���K?7�-�5O?�΅�m:���cl��@ك�=˟Y~[ɏo�����	��K��U��(�r��SӔ{����r���Ќ*��ɤ�o`�	!��5���Ŝ�U��תM��&?)�,��'6��;^3��vf|��FZ�:88��kD {~�VF$�C�}E��I���qξt3�qsh򼷈X�8Mx�������r���l1��T���P/���:B	`mnr����O���6CF���9"l�6	L2�	V1E~��[M��f��E� -6�*�Vg�WqU�T*�]�ʩ(��22�q�N��ѷ�,thm1�ki�/8Y���	�J����)-�)r���t׮���Z���Z��y��"i��'�g�UQ1�	)t��HSq�|:	H1��cU=���M⹹�Gg5���&j�Rƈ��T���u_I�z�)�
��*Kc^�!��Gk�R\+_��M�-T��i|S������z�eV�bN��̞�d�.��O���Z��OO���
�G�|l��n����-��ȩy��:D�Ѝ9����K��ts�k�?��s�D�0����0���N� ����<��2v��>��&QU�]{XUcF�$�a�ee�_�V�����i1@���z�t�(�HA�ҋ�|j
h~�El�JM�q�����j�����I!�R|F�6��@�+�4>O�v�pZnڐ�t��I]��MU������T�w�fY{k���k
�@���)Ɏ�?�ո���Yٳ{��_ߑׇA�&I�|1������	\�G���m%�nx�fMK"���|h1u��
�I,����d�$
|��	*���*By��Xp��g*3���0M�5�/ꝣݿث^�F�i_I�4��{:U�R�X�֓锚����%����>��s7�oD�5*��,x�{s�T�м�}T@�P�>���F�{��D��#�����؃yL\�&U�a�u��z��+*o
�&.�Qx+���Ę��!��"�헓'O���8+��{6�D{�H�/�S�� �sH>�&CE۞�޹{��)�7t6�0l4>I�O�*�'�9l���n�����WL�H>��ȝ�ܧ�0	�1郎#)"st�ɥ�}�5tr���2���<�s���cX�׺3t0���z�~��25��m���&&�I1;7�'�z�[�8V��d�6h:�y�r�c�jBG@�@q}�"5<?�zП��\4��;�:+�.:�� �Jg=e%����2'��s�20̓��x؛Qb���Ý���:ߛ{�/��u��k#��aM�T���<鯈���W�v�w7y�4�	����`�:�Q�[�Lb�G�0�@j��s�(�E�sR^a*sqtlT������I-�	�ii���u���Cg������&1�7!A�����\�m�ƈ��0�k+k�-��I�x�9��sl���~����R�'�Y��mR�eE��(��@����\���k���)U�RНJ;�%m��k��P���y[:iK+�ؼ�֤���ކ� �9^<V$W[����{�����������"6�	�R��)D���#���Y]����С�2�kJ�]��w�~��ӳw�y�/ȑ#� ���#	��gF��[��?���W~&w��c��=����/��{а{����p�o�� 5w�,�֙1���&��5��ˋ�'1vDQ،?^��Hv=�F�o
f��&�l������D0C���~߾}r��9���� ��S��ܹs�J�Pv�,u�=u(��~~��i9s�1>�~Fk�+�G�Weym�Pڍ2AtC,��E\t0��x��jd��B|I�(���j2�+�V��U�UU�n��0 d+���7m:U
�N�pZ�ԣ4Q)��{��Ջ��s���(����?4k0���eyy�G��c�H=*l�칆/��Hvz<��-�r��~VX?ߓ� @�s/��X7�̧O3_}���m�� t��q	�g��V���I��lw��������k��z�-k�����o�Y��FV�i6�Ϛ^Z��Ҹ���3�G� �޽��t:k>r���g���^��w9�U�*z�+��Τ>��Ƒ�(���'U�Bi��"������t~���P�?�/<��*�|���^m�"�?[�\%�乤t����<�kȌ���,X�PSϱ)^�>��\ܽ{�?V"S��t@�y��\��y:�H'��g���^�����ѣ���t�6;S�	�winQ��C2?;O;N�J<ت �l�>h?�5?h�l|^&��}����r��m9x�@�xB�s�#5�0,R0��p1��J�R)D�0�B�B�)��?�wuRm�7eH	��W����?���b���xY#>%Sg��}�}�����<��LGe�S�Sna��~��Ta��\�zj-���y.FVW���
��X��p���� x�7�_uJ��9am�i�e%Uz�qḠ��-�Μ�j�S5)TJ�}B$FKKcS�4��;+�y_�9v
��pW��B�!��7X+�z�wܘnC�
_�˃��?�0�xF�y>[���FFۿn���2!����=��ݲ]d���� �y{�����=_��K��h����gr�B���(:�ݜ��Rr�>�p���	8�o�{���c���{YaC�?a6�R�k�Ho��C�<��
�띻��N�=���r
^[X=hT���0�+�w<�C�3��u�cÑ�$�\���Vd��Dو��.䞓�e~z�Zkx�.�+����/Z���m�1���Y�n��E�/>�eR4���%J�5g3�ۯ���3`��tb����t���!��~[��_~Ȫ2�3RL�zR�����3�>+����<���S����]5y���g?{U~��/d}u�/�����ʨ�V����E(�A`D�Q�$��LiΩD/8�f�O�^��y;�(.�0�BI��4�̄���r�縙>�VG%����	�җ�$��,�?�<�77���(�ܺ����ʆ�����$���h��ӧ�+Ιy���(Q��;Lu_DЧ�|��W_r��WE����PYr���|�36ph������{ �9�D�m�B������B�PEu)r�Ez���{'����)�<@VP�&iO!���C���1�����f�HQ��*����a�=E��z����ʨ�{��i�mC)ʛ���`?��̩���u}e �B,	����]�֜�Mx�9�c�c����6�[�x�p� g��J�@���4�B��R
���l��dB��|/Bb�Hؗ�͘��f�Q�H.Ҡ��:h��z��lp桉��r5��z�R��*Ң�S�Bl6 �R��G�PܒG�i��kKeqG:t8EDН9k9���t��^�$g���,��~"�� �,e�%w��N��V/��i�t:x5}k:�=���F�4p��U$�΍dm�V���g�yF�Ϳ�7��o���/��/� ������(�yem�����DrP��t���V"�O�Q�y��g<���������cu�r�D]S���c�AX7�W=�I����p9olZ5*\�)��&�=\���`�܄�r�v��x�	���>���Qa���V����c��_��_�L�@{N�:%�կ��>�9n�$�����Z�w�p3Q��,��XY�֌�L�ۜ �6G)��Yj�����+ h@��Qo:G+�K��y'Φw[�v��"�XE�^��n�m8�m���VxRt(��/�9 ���=�49���>�i��o���yԪH�y�z��p�_�#��$񩫘U[I��A�Q�lo����A�݆��6���r���?ƍ��_�钘�ҊhV����l�x���q|S~����W� �A>罌�k"9>��۰��)V2��і��w1,0k���w�y�{�繟c�"��fi�c�%�� C��6��\���"ee�7��t":��p�y�V�=DQ�8"��NG)R���i�c�2SG������{�/:5�@��D�*��m�<sAZ�%z�ePѡ���6���D���h`��Q2Q}���n�"��Ֆ�PS����\�]�PΟ�����#GH~��/\� ?|�%y��W����[t\����~M�\0t�����C�����ٳ�����a�V��e�T
� ��M|zY|#�8�ԫ���$Ǝ95agnU���`5J��Q(�1�*TW��6"��4��È�7�ֱ�:n����%F\�3�!J����c�~���k4|H_a�@9����j��X�-Q��l�d1��Nq?4^ӈ)�s��s��aK��������
��`��&���N*Z��P�B{ʓ�Y$a(Ld��4����R�#��H6!������e2��3ơ�7R4qYx\�O��h/*u��򻢇�<ɷJ�5��i�Iz3��jE�9�8�E�]�{e�������?��[մ�h��0}s@��x��ji��E�k�V��g?C���g�1ǀ �<uB������y7������ˏ~��,���'��@��V\�k�.V�����1��� �Y���uޓB�ŏ�#B��V��s˅eGo���gv����N��#���b0��,=�V���
)����p����3Pb�\Af�J�"'�S>�� Q`��i�軕ה�w���x�6�i7.En�q�C㝊(/9����	�����41�L �
+m�{��g��y�Ε��)��i�J��o�$s����ن6��t*�s˒vn�<�mn���,��3��|���}W[ A hV9�:�J:�Y����O{�{��Ύ�h%��3"(� <�h�]���{.s��ō��e�j4@tq'��z�/_�5_D|��d[EfOMI_+�c���o��O���%�u󷺲���\�tŁ?f4���^0�-�M��{��ͭ��e�=��:�1����� �}f|�*���z!kS�k����/> �	��؀X�UL��h������B��Q����>�(��<Ѳ	��%^"�d��#��?�y��!@�E���[�������J ������dzz����[o����LLMȋ�:V���VgN����f�����t4y�K/�����rΪ/p}
/B�)Bc(h�s��R�/H�L�N4���ْğ�xO��qF��;�x����o����.܊����z��zc�Yܧ�W|�;��h]�?�zbb\6[:Tý���Џ��L��l�}��>��=�-t���;���n�ͼl���鞮�������/��9g��zR���u��菞<�u<<<"�Ν��_]�������a����������%͖B���~�������?�L��bF���������pr,?ʠ�[�*V6��أj�{�2��1���`������J��`�%�4��yy��Ze�~d�h�I(�z<�A��<m�[��\�ן$���HP��T�q�-4�`@��[��<��>=¯<��u�U�9��$MI	���J�%i�ױI�⚶�73�KP9��m��z�`dgg�CH�vdkk]�77�a*5߃���X>�yS<��g���Qo����1� @�˸����[�����G��R�)��EI�-�����������f?�dYV63&ӊ���?b�d�^�n��"�ӎ/J	��&�wy[=n�?~,�w'���c��8�<x����*�k422*kk�rϝ��GqS��_������ߔK�/����K�9@/���c�c�iCH�>6�L x�Έs#����]�Šw3�DE^ ��si��Ի����B�τ&�OA�O�2 �U<�^RY����)�D�a&3sp�� `�Zg���aܑ�9;3��Դ�k:IRO�֪����iA�����='t�M�q���ݸ'�kVc�.2)�ZU�J/C�ユ�������7rq�"�d�������������o�#�}�>�9²����r�C���-@淾�M�p�\�0'������?t�60Yp���'�T,s���/	�6��~���k5� �I��}�(�v���=���noU�j 5����6	�Z�ۣ{�30P�������_Q�&�s�C⁇y��o�n\�S�B�u�u��y�ES �d�=�&v�=���b/zq��H���V����$�䱊�8���AM�yg,�w|���.��=��֖�d{k�r��(� T�e�<mP�LE=s;!Q��G��p,d�����2�l���hk!Ͻ���Fe��2�'x�X�n)���V�w�ƕ�����9B^���6��s���� DʺOU5A�e����5�CH	_*��L�>�?w���O��OrinN��d{{����{���T���j^�[V��e�����9�{�y��zۻo��I
�D��%h��$����g$bqp����A�������B�݃��J`c�/+�^�H�Z�b��q�i��L	(3N���� ��V5C�*`+ J�n�c�A��G;	��ӎB�^��'�� ��J�ϪT*�,U�A�R�=��?�#*�����;9{�,��,�u�C��?Ҕ���?��*?���e`��^�+�/���Su͒ q�|������m��ܤw![�7�_,c2����@͞�Q�Q��Z��h"��q���v�ؓ)�ZdY�=�S�	�����T���������-*Y+��P���b�7�X�-�3$!Y6�L����^��A�{X��sZb�#����>�{@���H0���������X�<1�TJ����ߓ���D�iY�8P�D�OK�a��2YZ^$_����Ś�u]T���c�J>>�ZU��^`����Lɓ�ۡ��B�է��5gF+�s�E�N�`�xpX�2
�\:vq��Y� ��(4��������<T����AAZA�~@���d!+7��~@�cָ���h�)�`��8�20أ��$��	e�R@�ߋ�B�E�C�[��RB�2^c�I�>�=!g�B�C��K���D�h�l�EK�@�tZh�@͢��A�05�wb�!߶/1w��%�j����.tVԀ֦�|�-(��+f�YƊrTFXϵj����g�k8���C v�g ���B�����48������ݯ9�N����Lv�E����(���ŵ�����������ȟ���A�}�fF�����#_�9�Æ�P�X��ߗ���3���Nn�>-�m�h�, T���i��!������t�2p�9�,L<C�{oH��{k^jG��ۍ�f�a�����{��5㰂���zup�� ���*Z1�B�=�N�s����ZE��h���͸!�|;(w5(���#�e�_1��2����t����`����ӻVg�������v�v��"��R^�%!�q��S42հ�l���$B������l�P�Ȏ$yہ������:Ƅ�B��}X�f�w�m��5����#A� w�
�z�y#d�0x�N�>O$��x5F�c.����{��n���L��)�n��_����i� 8�t����(uw-�j��0����[�RF����I�tMf,T$	 û��ҷk�%����d@#����TH�Z�25�[�!<;�R"Ilr��@*�]�yI����K��D��U�4X
E��F-�
G]��S,X�xލ�Q�
�%�e��d�B3���/��{=؅��� X#p�����E�>8����HU	Ԙ��˴w�q=�@�c��ƍ��ʕ�Ϧ�n� c�Wa5�w�~G�z�248 ��5zݵ�E`^?8��`�Q?�}���ɭ۷h�]��Pm�{�A�<B�|��_�����=c,�),������p�w���	�,�w|G���Ғ���ȭ .���d��W�9�1f#E�96��`��m�8��:}���&��i��;�/�|
m�ށ��}�zz���/�XM(_�7)J&�6��Qy�I����� &���ˢ��f�ty[!Uh��D��SȞ4�B]h
��yW���,'��~���*���V}T��9���C���~º�>������X�<[/4�1^����a�8��=������Q�fp�$"I����{q�J�'����=5��Ū��jju��bQ��ɱ��2�-ȍ�I��YSef��>�i�qB;[�8H�ns
7�ű2�q/��/f�[����6��E/��~Om�yz��1��IxV�&����Hyj����n�pf_eޅ\�ꢔΎ>-ew4���/	��.#��AL�=S�6�� ƾ�૕5�qȊ~�zU�=<G{gak4�7m%�Y"�����U�;V-x'{���套^�o��,��*�n��7�uw� �%�y��cP�h4���бr����ZK M�J�*��i�����D�FۋS�N�~�C*k���K��\��$V��F�W���d�x7�l����ȗ[�P��R��<���3����XP��<� 8 A���<;@���������^�p�Ҵ���-�dX)��i;�C�9���f�%E
8�����(O�i�� T߯Q��Ұq��$~4�Q�kQ��df����I�6�kt^�S0�%�g��%La�x��<�ńkڙ��myX>4 :M�zf�A���~��-o`�v�����ᾬ,������rez��5eF��3{k�t� ����ш`k��:N�t�r�:�i��������5.��3�O>o�(o�l��H�V��@�s5�.��~O�b��ܴ�����e��)��n��i��q�<Bd.-���q[���D2��q��f�!%�@�}_AIg����x@�#xe"7p%X;��LI��c?O1�IG���Rxt��|�B. V1l���|��J����+�EV�q��{К�ښt��:�Yc?��| ���U�i������#�$�ߌ����$��J�N�a�:׮]ن�e0Z��w�0Pm�Рv� m�<v-3�(���3���!>�a���m�gz�+_a��vٜm6D� �L�m5���x-������/���w�{2���_�:_��ƃ1�����5�c^�ثw���\�&	�Bd6Nƥ��z>��Y&����v�����Y�"�b�T����y���=z�ǆpXM*��-6$�'4)����ߓ�"��_h��Pi�ǲ/�b'�=l�b����į�w��ؘQ/�X���٪��7�?,�hgP���Z���O����=ّ��eY]^�+t�Gr}��y��dk�B|Y暭��a:��#�eZ΢ �k1E=e��b�DTl��ih	�756�M�5l�&�)���#kY�gS��T}�����]I�?�*{}�kt7fW�W������ �����j����B @qj�о#�@	.x�-�/K8nm��w�St�͵��vvIHT��R��6���(O&b<���h/䑐�F�)�i�^�4�ķ�<�c�)�<����`5���Q�NR�����|�r
7ԬY]��U�@W�׸4fi�|�<�#�l����{��{����42+R�>B�@A�w��@ ֘y����i"��������yVw��Ҏ�p
���q.~FQ(��c/�Si������=C�nS3{�p��3���j)e�ߛ�m�c0�g~��7�3�U }8␏Yש-6��S�e���J~��kޚ�ke�,|����V��P�Y^��oڄ{��)e&]�[���u���a *�� �����(��,qEE=�>Te ����Ռ�����Gy�
M��������Z�/�xO��ZG)��O���J&F�ޞ~�}�Zo��oHFF4��sr��i�+ WQ{;���e���+*E8^G�Kd9a-b]r�kZC��e\���^>���g5�>�g?Gk�����Z>_ǆ�S���$� 5jA�X���aM��������ݼ*q6C�Apt��0�q���w����TbT��e�}�"4���1��B "�{��EֲA]�=�WK+�V(���{*�=�X�����#�8Q�#��M]4Ɏ�"E�iaY��	� �J�+n���iVW!��!hghK}�����:�7�@s�mkwC�N(��Nk

���Lغ��lOi>���a���@�����Y�C�O�T0�++�.�
����"c�<�
 �����#t ��޻���k����q�ߡt��ϭy�Y��{�٫C�=a<�;s��%(pE:{�7ʠ��=��ҭ�j6YV	��!������e��>_G(��ٳ�a�P�����K4@,�����yp:��<�0E��dI;	K�=�a,�p�$��;�	Ȭ��U�&������¡7R�3	�����4���y!=b.��ǍCG �s\��)`Ql
�K!7���v/�=C��]|�ɕ��sd�^�8�F�:�A��7��J�0&�]����&���9���U�ʽ)�H��n�;B� r��h{��g��z'�V�^3�=>ϲ��� ��O[�q�~�̱�O��
��R��*��%��y��9N �)	���چ��V@+vqǡ�n
��R�7s[�a�� �="�N7�{��>����%�����f����[�&��Ĉ�^b���������G?��|�;�����w4Tcڦ���M�Rug!5zT�i�,:7̠YU��2`�96�"�W��tB%+1�[����YѸ���
�i��
@��ƕ�{EB�X�������2�x~�N� �`��7a�������P��+
t�x=��>'n1��r��-�˿�eyyŃ�$�eL�Y���XH�<T��R�3m@�	UW}UTf����==�w;����SO�I|GTre(�}֕�Wh�=�@Ϗ����ȍ7�`�����{E�N��+@s����3�
�/-IQ�w���{x�0w|�A���P��k_�K/���0V ��B��<���"�ʯ����U�;�Ⱏ�I��3fmq��䢮N�o�	����^d&خl�o8 �S���UY�9�-��.{�7�a�Bq9eK:��?���]�(�ν������y�8�}m��� �!͖���܏OR)cM��i!~��-��=-w�<��u�;�Г~�]_W.]��_zY� �p��zQ�Aŗ��(��8�y�({�hH�O���͒P��FA��=B1�y��:����%��I���\[�T+�%<YM8�k�=f��@Rĕ-vmO욵�\�}V<1�n���%,G�B0ww9����n�S{�>�X�)��n�ܺy[�}?������)���*�}����|��$��|�2�	�ߡ�a-����.�F�V�%�r�7XbO+�$G�^$L�{v:���+��r����Mt��䱳�\��\�lbޚ�<=������3{Ro@�W( ��]�6)
�ފb5V':�~>�Y����� �� o�t��I�H��Y���uwr�dr ���N��~u�{h��}���߰�Z���P���U�s�԰�`��}�40��\H��^t���L�ּ�<� ���� �ˏ�WY�u �e�]zk���R���BJe����dH������� 0�s4���,+����;� ����< H�񃆊�:�;�C��P:�:R�#��O�k�;���H��L�P�}/gg�-�$���|��lP)�3��.[ԍ�ɺ7��q����\E3���	�x�8���-���=���J-�vͣ��%#O������L��ؗe�� �`�2�Ly9�X�@q}6�MU&4��"��{�	��oY ���=A҃��.�B� D��W�&�Ϟf7jd��8<:6J��V5L��=�k ��TI*A��\[�1�0��s6G�p�s
�cW�P�§�v�)��3�|̠x��E/G�]%�W��`jF�	"�ȋM4Z�gDN�x�
<Pf�:)�S�k����r��7qy�#��Qk���󼇊�c��YT5*J�6�|��n@ȔG�eX_��!xB�{����������u��q?�@�����PK���I}Zɑ����tc�5:Z`���=Z<�r,Pkt�γ��J,:����ޏ��b��TJ��=�Q��f6���e�,/G���x�fRyE�pk�ѱ1Z�=�4�g�l�[��ܣ*���R�,��==�`ތgR��������S}����I�-Zx��=Z��*a��Z��?F��ڕ�2}�LϜvz�{fdxP��5r4��/8�쌑�=qk���>S	�n��d|��	�K�k��@NY[E؉�j˾B���J���fsឌ����;%ۓ��k�S�f�x���V͡S�-���dh���}Z��l>��I��Aΐ�^�zE~�~$cc���$*�h�����Dr�4��\=�������ր����3����2��"��c��:�����5��̓۟�[rp�!�#��(O�#շ��6*EC[�G
�7��rj}+{x?,|"�s�rtdR���:���gb�w�!k��4|�Q`��o�ltN��h��D�0YZZ��I�G��l�*0�^����޹#?��Od~��'u6�D(�;���LOM����LL��&�
F�0Oxo!��i���x�A�����+gu��A�u�@_��N���#�a�'��C&���-t#t�o�n�A<S�pԧ���~]���&��ܸ���{����}�0��<�[�q�ψ��3K�&����T�(��5����g���ä_�t)�u���W�iT��UI��u������yB�m�*����3+pmߵ$O^V?�x-d����?f=�/����*�����;J�����5ZDN�q0�P�n��'1^	�ƈ������Yd��Wx�\ʺ�#�I��K�CI�������yh��k$卤��<�K�����˛<CkNlyO^5xф`��sY�UC�
Ja)Xw'u��#�p B�"�Jo�ƏH�N�{����+ҽmldH.]����S2{���8���R�34��?Y��:��«�zNA�u��� @69�ϊC|�)<�Ø���M7o���k"�/Ke��Yh���;`5�;�䉻���4���V��ڊ츹����r/W�+�q��O��څ284��1\��� �H=���"��3y�J@����B��F��Ph'���9(_TG�ڵ���I7>{�����{@o�a}Xkՠ�y�CCW)�~kE)=1���	�m��Ib�u�����8
ח���e:C�i�{���ǩ�p%&+o�s��g�鵵��ݗKsWYia{�YN�`�3Pш�8~���9`�.4������r�������;��N���Qp������m��!�2�5�7����`��j�/��;b�����Ą\�0G�=���j��N���/]�C��Z�4<��t��W���Z�i�{k�}��m�n,\y�^�k�`dW#	��5 `��B��x�n�̻����.�1�T_D��+WH
���_�z �D��F��{�G�>K�x2��v��:�SQ�,f�O4�S T	 �X�����_�%	� 2���
�8�ES�w�%��?He���#�KK�'d�o@4f]a-�$Zj�>�Xv���y��-��ͳ]����Y��ʃG������/�������.�ctt�c %{��u_���ֺ�r�;ײ*���Y!�NO��Qd�y��V�/����"�wccS�H}�u�D���NH�O��I��O9���o~�	�aY\\�����ζ\�rI��@����˃�p� �t�Y�@��_5��2�J��h���*�ăV��,��p�A8<M9t�~̝3����5�M�%q`�=2���.״djbFZ5r�����]z�z}�Ӯ����vB�i�!��{�"���r�C��F�lػ���R��}A=$,/-�3���^C����PT�[hQq��p{��������È++k�� �J��{f/�FM�������p$j��T"�F�A��GW��Vj��0ˀ��ܔ>��ky�s��ųқ�^:��C�V������x�֢s0??/���/	��U�{������)�����8'�Ȁ�9i����3?Zx�}h��.�7_��d���<!M-[�Bم=�ޯ~�r���Ǚw��g���p�ᑑ�C��G�'d����;�������,�9�i�v�=�Q`)/�Cy�����xn��L��an{C�8L�[%F#���J�L�8�sqlcX�8�v^~�ev���n9��Oa�] xo^|�EZ=�G����Og���Y�0WL"�x���jƂ�����DV�R�D=X�X�h�����w�wT��׸Ά-DO5�7������ {~�	qT 퓞��OE�V%Ra�wpb������D���C�����\Z,��|�A:4+͟��iyU��'ѧygҹ�g���Feh�)xz����I ��֪_���voը"lӓQ��M��}m�It#��Gh2��A��������Y��]�3�(99>)_{�uy��7���xr�v�={F��^XZ\�GN�C	���J���u
�ZC���R�@�$Ƣz��\�htY��R,h��Q��1*R�Z(Ne@���0#M����qdbU�^�RBe�1 S'd�j�������^{�Y�3�{PT���R7oސ���+,\�pm䚶��z_r ��2���)�{(y�x�]�ay���is��2������B��34��w��S'7�/L0���!��'���l.�
ù�֝���'%t�.R�����?��17��K�>,�H۳A�%� ����|~B�Rr��}hND�C�W��Yb&Z^�"��B��Pml���\�v���:�2^�3NG��_�D��kr��
?Cw��C����O�o�����6]V�׺�D���y�����ߥ�QT/&���+�t`��V��*O����^����3�,d�s_�xɽ>E`L�s�c�]��g���q�_�����UH~�#�z3³d�׋�����X�u&h�'[�����e�W$VʘLlت'V�2�]G��-���m�
��I54n �
k�}@ �|xu0�?��O����ef�!�n�AF�B)6��ƣ�wwE���!�0F�t �!4�*�n��g4���B�~����mO.lx+��6Y�{�=g���t����A2#�sa�5��I4��� D��	ɠ�1�E�Չc`%=* ����B���^vC�R���`���D+��z^]ݠ%w$BT�5�� ���h�~@q�\�9k-�ڋ'��'��q�= t@�d�	I���.�����y���&�C�����P�C��8e���rl F 0�	��A����}�?��� ��4X�A���9�ƩK�Y#)��-�V	�mqV�zG0/]���
�Bػ��w���_\Z��n�=�<�+
@���P0M���4��	���	Nŷ�0ml5�c@k79�D����R�S�WW������7��0KJË��c�w���_t��X��3�ܥWa�vގ��0 �n���w�(y*��	z�!�˒�&;�0SG�)�f��a������� ��R��wd�-->�epi�'�~w{`q�` �,Tf�a�����#y��1=cxNˀD�!ۛ�ܖ;w�++�Hn���sՇ�`\҄������Z��xc6���Zl�:��ʴ�I���c?��C껗_~I^}�5�|�*+y�VQ�'�`�o�o8Y�JP�&���0��|��BF����E��[�� ອ��x<��S1�%�	����ݨ5�Ȗő�@����;0�sssLq��C� �@����� /q&���0W$���Hm� �����yAvN9�ό���f5���æ��n!)S�xt(���)�n�>��^��AD� I���i��p��>tBptxL�6 �vd�Ym��(���s��W�y��� O�
H�1[ʔڂ(��T� 4�`+�cĂ�N5܃E��Hr+���Y��rk�2Ys�fks�)�!*��ų�l�`\�X����e�����g�wp�[���zӧ�����;X� ���ܿ�P~��_�͏o�}<4���>���`�09==�}�j7�q{l|�^��J�SQ��!؝��3�D�T#� 2���D��t�3�i��2�lX��,eF�{����0�mx��� aۭ�^�tς�y����c���*v �+�e��U��?u�:�ԛH ����6Z����m��Kf��+؉�e	H#�7�L�f_!7��P��Z"=�L-x(Cz��8��><M�NI/�\���9כ4�L��M
�Z�=���f�xR�_<Q1�߲�Wȕ��b�g�xx#&+R��j�� �)�V���ˆ,..;yx���%�P�Q& |�JUAmoOe��;��8��� �ై��h�Ъ+�Nkn�6��9�b���^H����hr+���"~�&sz>%-�g����q����_U^u�x5�vv�;��$��K/�86 a�-�TI]2<P0��<�x�by�kS�^G���3��K����)y-S&8<��D�'
�k��xk�a,ؐ�� 8��`��8LT���s�;<����ϐ:� +@�P�t�{J���g��h��&ݾ�����ok��tZd�:.$�_Z̭/���k���9q4mxv��������� ������OT���6���~�"�����ɩ1i�BI� v�ѽ��PPZq0��30T@�"���,�.=vA�tJB�/��B��O�ݝ�#�z�; KH�*'Ny5(\!��j�)u��ņ��	�[0j,���-�PrU_[$��z�~����'Ř��k�}����2=}�tuB��s�s�h8� d�<�*�m"C�L��r�I�w��� ����M�3l�=�����ʆKƟ͞qhR�f�/��W��rZBaN���]��.=Ȩ�6_n||�Jbp���ꕪz�����sn��?��|���P���l:K�N"x��ŴҦG��l���q;�M��ɑ��?:���E�*6#m����YS�(�iU�J�B��X^^����t���5�9�e1�c���=���f�'�����Ь)M����s.b�B�N\�>��
�� ʨ�8����b{�$o�l+=���	�N ��/O/D���1�f��d ��P�#�~��r��)&�h�(J����G�>�a� 2�n\{j;dV|R�N	F|��m�i6�r�+_�����˔;0�����������]��ޣ�]��X�����[,e�y<��x���y��W��w�ɬ`��M�o��R
��������}�0���B� )�č}�ǉ�1PV��#�BhaP�1$	�yY�����-��@�͌X!- �+�e����l|��tF���"Y�p 4Ă��w�0)<F��'�����n�ި�b�z:�O���9S�Ze(͍g�[#��|���J���R	7桬�m0���TZ^!�V�>,���]nBɻ�/�
�ҽgT���&�b�Kwg�+��X�F�K(&�n�Y�;o�
����Fv�k����N2��Ј�T{�k����~_���gX�J)*�/Q� �S��$�M@�ѭ��zt	��=Y|�,���5���o���� �v�nkΨ�+,D��^d�����Ã}�,�u�&V�[�~b��R�Zة��<,*Tw<���\tV/Z�x�����
�}�j5H����q��H4�|銓g��&�&=Xo%7H��W�F����lmm�Uq|�)��Zy��"S�dC�W2F� �5da)p~����FSj�Y;4�ܞr�e���;�[r������	'b20��$��ػ�)V�0�1�CAIUkF�Z��K�V�{b��zR:?�f:�PRz�}U�y�+���[�L"���g9�@����=���9�0�[�����<}�,�v��d��x5�r+e���ۅ,�p�����"Ǜ�r�����t��z������#5��,��&��^;F(�����u^}�UF/v��H���7�����D��FBp���}:�^G�IC�������:�{�=6�f��`i�f��J-x3,,d���u�ü=������?�gV4&�Da|�wM�@�Б]�d!}� �@��7��2pj,U���Y���_F��R�H,����p�� �aI��{�&D
'���>)��;�73��5�I�ĸ��WB�V�瘴g� *@տ��zA�~GGauHv��Up�� 5�BKI�%���r��%��/;�hh��98[�n>��fgN�CӬ7	D=zB>���IX����Г����8�9�l#���� �}�a��{���#�����?��D[��߾����=�u�X>Ƨ��p��t�/`ݎ�RB�'����,�g�fF� ���S8�tγ�jƘ� a�z��s��}P!usU.~�C*�T6�w0(��kz9<K��T+�:%�⁣�������#��Y<c:,	���������elt�O�y��g�׎0��z?&��EٖW����i�L�_�\:_�2�A�<p��nxxT��&i�@1�wr��]y����{�Ј͘}^��%}-�4K|����&�rn�pO+�y[�9�._��*AӁE�Pq^���P�^Fd�*Q��B���;w)�a���Y�|d��-x�%Q-@+n�}�%y���G�8��t�'�Z�[�˦����y���ѓG��'�7u����� h���o1^�&L���!Sɩ�p_C���Cg ����Ȏ��θ�6X�V�ޝX�՝Yy���Oj��@��42�
�����,��*�Іn�ׇ�������P,\�J��w�{�{�xh,EG@�R(,`'gg5� 7$��a���������=��R|V�L���� Z6kԬ8� 1�&��@�����6�ˢuk��T{�d���N��K�W����ϐu>G��>�����b�K��6FǍC�V���ퟲ�HG6I��F0��������olʨS��3���U��i��P�oM�J����Έ��U���,
�یZ�����Ư�U�p�-j�ư�' ]�
��Y9s�4�ݱ8�h�ܧ^2�!�)A��^����p���S1�sQ��^�����(���i̙�9��o�a -z�w��Ӣ{�>	@�c����M����S�5�����W�����~�mڭ���a\�Jb�5�	�*����L� ~=����Zi�>�'�+/0����Q��=ׁ����d�uYh=%f�V�dE�R��+wF�<����,<��{NF\�r�\��,�P�\��@�X�g�J�^b(7�1����P��A"ў���G�I$�#�I�\���3@���ɹ��MVY��ø�y�	�6�v(a }�1���Cv����$؜�2lQt4�y�1�E���#ˌ��2*��� ����E����Oȩ�^c�U_Ҏ#p�|1`N?��N��ȇ^C�לu`�[G�m-Z6�Qo��k<��Rz����q"�'�\K�f��X�U�a 5n{�n�PH�r����@�4Zp�_@����e�S����O��L��ŀE �.~�Ed$f���"��&ܺq*�[��G	��^1x~#�½���A �"��_bx�������G9���l���,�˙3�9��	�ă�<���ب^�و���<>�{�#���]�#���j��!�S�[�_|�*���f@ �	�`�I���zoarL]��c�IV� �D��Pψ���㳄&��#&���!���ݖ7��g�*�cP:}�Y�N�=Zx"�[���-�T���6y$�T�����hZ�T��6Kf���2%�黁E)�_�A�gZ(v�v����!�������(rZ� 8�|�Urj��ի���B��?��u����TQ`ZI5]�#iow��W���r�qG������^�G�7D(}�=����sӐ�`�F1���h��hz�8���N�=�2K�����ܲV��%�-n���P�<�S>�����S�lg�2��X7�ȍ�3~�q������$������ǜ���	�#p����1������� ,C������h�as<I���CsA�]ڟ+
7�6��eVR���@whk��I���޾+�k��/�B��	�q_�ṣcL�����������[O.� x�P��ό�rI�__`0�w>.��ibaf��}wr2���Y41	���Z�x�ʲ
����5�wv<u�jld�Y��`�rA`��NO˩�gB�Nw_��\H��OS�ᭁp�{�F�E�����ڧ�S��[���G�Ѝi�Zب�l�����6u�����T�Õ��;���{�9��m�q_[���(X��shI�I�HvZ����,�������Z���̈I�1x�l�ȅnx���i�i��3���.�;�2<8L/{X�fu��`.�q�O��p���z�׬���x���/����G���n������+n힢��q ��
���>����e�+��)�v�A8������Q�zR#f�{S�j��1������JS�|RX��%� ^&Yؽ��ݾn6�> i�� ���۬nJ+T��� ���V���{Bh}V�aS���E����P�����ǚ�u�?ʩI�i����c/_Y^�皕x���8>;3K9N��
f�7|G�&�u}]A�,������������_���X���i�fPI$����2x����^���_�����J�gH9*/왓����y�S���ʂ�~��_�!�?��k����$�"�iU������zdx���έ;Π�,�R��H���n�%�z�-�ੱ��b���� �:b�{}�(t�߭A_�Ϝ���[����ȡAݦ�c��t���~6�00��,~�]��z���X���d���c�gq]3+}�X�a%�ϒa_P5R��ծ~��w����Y60��eA~�+��f��.z
;��K͊
\��au�����ΰ?��Ԥ/h�)�?Mɰ�P���|�h�w����pj>�aa&|o��yx���RӦi9c�G�U ���8��u�����c�sg��ijz��V�^ ��!�6^�	���!�\�0Cx-�7�;�Y�
�y�
��+	u"�r84���Te����¶X�kp%��� ��	� ��BHS�"��6`Ӄ�]k�:�Q��:?��[L�Ƃf���N~��ߒ�g����=vw���0�/H�z�9�7����������!	�)�EYF=�*��'�>�RL?�k���,�+Lr�	�i6dc{��rd�_�Ν��jŗ�P��b��V�vs���G�>������+S�SU��C?b� �Pї���W���fC�W�O�����q��j����G��'�'�Cف�g^[�cd�#�'C����o���5>59�ٲܾu��?<��x��8�U"xu"-)�?�LhL&t���:eFl��K|>n��yߩ��v�F�� � 4�js{_ J�;O���r�^�u��<x��uC�0rhLy����y�g����>ij_���͉�q���!|@��q\+h�� ����u���Yn3��U�U�\hs�㹱F&������q�2��^2�\ ��'�	j�T�w��=��q"��JI����\����E�Ύ4Xv(\��}@�Է�|K.;����S|���\� G������U�7��ׯ���x���~Q
�������5��,���z�������w�#��0 �;��ᙙ�$ Z][��Mxh�:pB��-֮)Z
��[/��UT��iL��[C�����
�]D+�I* K� 2J6�T�A�� ��&2~P�;*�*�r�^� `���!,`T{��^:#W}[�]R��@l~]`&���q� i�X�*(�Zr
5Y��A��Z�[Ӷ���c�Yw��9�/C�tEl�!���:,�U�%f���A�)AN �]��i�6�(�I�e��#3� ,��1/��+���������}Q��^�=7Z࠸�eC6�����}֒zK��b�\�88D��zh}�l`�U/��-� >��q3K��DPG��`�g��q3�>��e�V��fgdmc�s���ގ���{T��ϟ%YUC���=�F:8$~c[=�}o޹���c��й�=��s�w�#?�#��PcF\������C�C g��$�w�q��p{,p-��>�;xvo��&�����UVȳ�1�	D�Y�y{�,�`�^� ��ƵL���?�~�@���z�����0����}g~�*�s6�68�r��c�@冀${�"�&Q=]��:Q�Yf*"����4�����4�Ԕ	�q�#q/��I�@��8c��o{�@5��4�>֕�cf������h�VV}ff���f ��J����8���řc��u3/[� /����4�
���f��qߗ.]r׫����ܹ}��ˆ��Z���ߠ1|�/�N�����C�k�8�i6�VX���!��TMt*ފ��ف<����]y�L��)@����!��Kwc}��B5i���n�z4��]�ŚI�	��6��u~\��u�٬O�Dǚ��^��'�<���$����J~	�-��m�[�IůՄ��fe:��bSp����Q�ד�3�q�ٵJ�t�P&��	�=}5�ޜ����^�b9�z"V���k\����SaT8o ��������niA6���z%�9��0�,.�v��� w��=4���V�TC� �Mr߿���33���euk�`' ;R�Q�����1n�L��݆��w8�95�tȄw�tz^�Z�r�N�M^�@:�2i���GH� ǡ����1I�7���ۚ{�G������`��>�i����1�^�z���P�T��pO��"���|V�T��8�C ��sR�O#.�dxbT�ഹ{z�����j��,.!��*�|��PJ�O�܋x`�x�JBr1t�Cw�u'����̹�����Ζ��J��?�3�`�3��iN�b�SZ���<�(Ƴ'��M�� ��$G+���a���u�=*��ra�"�Hم�q{dKZ�4��➟�P��<�T�lnnh�+w=�0��)�g����1��Z"�tYXeb�8�R�����4>�Xo���Ӳ�6���*��W���&)�oy��G��;�*�M����2�J���g����zb&�Ǩ�S�7�e�U�Y!l�����ߑ����CC�����e�.hX��n=޾}K��ʗ9�X����*�pɧ!t:<2j ��� �I�zB� �J�����[hx��[��d�x������P�ğ�5����	[T|�����(a+�d�!P���ăAu���ҫB)x�P �x��K�e�"e�6�
`�s@T ���k�3�XE�"�y��Sn�.m|�*>��3���C�W������KL6�s����/v��R�n�ƕ�]'��3('��^	�.�T�l��0�4}yI���^���u���m��ñ	)5F��BEa��/��<��]`��
�l��t��xZ]������|�I�]�� �����=�kPqυ�3�6BQ�Æ4[�3��S�LЏ>�($�X?��{��>|�\���i��nƬ�Ҕ�&,� @�9D��{w�K�j�ɮ1�Kx�n߽��MT�xh!��<�0������-�?�#u�Ɇ�u�]���vjz�	&��x��'���}��b!*
h���x/�	'֥;F�t�F�*qP9���V9�Y����n8,HĻgf��`�������#P�#(��+\шI7�t����C�7oݖ9`���1�ʬ��i��Ś�R�K�#�>�	�b��!)��^�S���h� ����B�yv��C�U�{��17w�u<H��ƗYPI���$]	���1�/ydR���y^�_w�Id�F��9rff������m�g�f38t޾x��pB	�n��5��D��ZAa��EEW(+�F��C��\�_-�����h_�a�Ҏb~][�¨�?LSD�(�dMkD��|r� -L�&��)"�����Z�_'��p�$I��J���p�`�b�����Т�]��κ,D'4�h$�{��\�};������N����I�@�;����]�i� Q�:\�(f�/##�����$� ��������b��jϠ[ب�\�1=Xb��xO����i#��ִ	m�.�8 ���\�it��>G��^�N���0*����0ü��r���r:�;$YܺuGCQNn��E�?B�$� %��8<��O㾨�J�adU�5f�$�C��J�0T%��C�~W��)����d��e�a�ϝ;�靛��a �.�H)2e�)���0�������tZQ��5�P���q܈����/�$��N�-_������|�����5�xT�y���<<�h⊐����ӛ��������Ed����W�ཞ�(��8V�?��Ĉ���r�AQG��$rYŃj�9�G�����,��K��N�#�|�ɉ)�Y��Pr�Q��h�u}(kkLDR����C�b���T�E]UO��X��qN(�j�cQ�uaqO|�勗�:�  1���7|�azg��'���{Rs����$"ߺu�@���K��IBQ�[��m/ނ	���q�4Y�c���؛K�Ȉ��֤㻉4o����2��G@�C����Ǝ��]��B����KN�͹u�G�2?�@W=<XX'������{�+r�W���.Z,۪���m�cJ��\��|�g�l99>��/�a�=t|f̪�z��Y��^�d|��Y����[24��`��U֪��>�ܰNL[S�!�4MX��2
1eiųMH���G+��#"-��;�t�C�z3�f�����#óS�q �q.����c9{��V!ȄAm,x���U#/��WұOUn�0�C�z49�ѷr���e9`� (��M�{�2�Jڃ�P���A�&��0�`�':�L�k;:wCqa}�*��ĬS����n~a��(��iV��x���7x<�)���vV���'4
��ڤ^���s�\W0i'M ��A���eyuC�V�X� ��ԩ32�������ߒ5g�b�����Q�#�:�0��ݿ�M>������q��<��zƩ��s]����n:��h��
�Gc���Gmzv�!��%y�_���i�l��� .C��ťE�����:{������`���%��a��z(Y��P�>��_Q�ـ���Bma�rRǉ�t�g,&�#���F�UF�y�|d�t����`�qѯ~����{��y�
��2�q\��>������M�'΂�vgg��R��
S���£y��)�R�֣�[]���κV�����7��8��FV�<� 8#sB�C�&(��Ni:�.��/���|���l�q��tC���Ϊ���zMX���D��fE�<b�4	��j�ũ����h�q�t;�9�JE/ s_������i5r���n�W�]��877��:A�
 :U�޼y�������W�8V��4�w�o�_�>����ҥK\���<�.�g��O;�YGǝWO���]��d����X�	�q��2Z��S(�F]6ݺ?��+j� Ԋ"m$�$w�죳����̈����ZiZ=x�e1�@ۯ�ܻqRB�B��V-<�7���s��N�K��{���9MI�*S�����H��I	���@CXDj�5�մ�"��}Ӳ0D�ze����,��
�i��uM��x7��Y��a)E��:�C����C�� �:�w��M>�����W�@I���I�w�.t�F�Dp�N�9�Nс����0�x�\YO��;��e_��hwk��7�˄�ܙ�+�~)θF�r��4.��weߧ�OLL��ӧ��F̒��Wa�T����g/0y��?�� �,����Ÿ��:�Fp���u�O�vj?�p-_��sS�g���!?т��=gx=�S�gdjvV.$	���{�]>�%g�M�u�y�#uU��7��w�Pƣc9zá�-�~+ ݻw�}�@����/��Rl4��J?�m\�$+�a$7���g�w_��\��v�$��ܸ5&@�E{U3��=�(�Y���%�:X�C�5.Z�Hb,�����j�a�{�� f�9�!��*X8K�n8�3ໍ�}=>m<��/.����LI٦�ƖxK��2 ��s`���O�Sv-�9����XC�Ρ�g�������/ʃ�w݂^�{w���9<�'��x3v�͸q�"Al��`�sc���hY��Nb�1�_�ӈ%ԦHY��`�eVcœ`Wem��^9�+������ǽ�hPf�#�	�����7)�P*���!<FE���aG�2�s�m�>���Y��w�2���ӭ��a}��ぴnT=�C_'%�B�����s�Բ�ƪ� >�k�����aۙ�`$ǢƌG8����tU�!���hH�o���`��u1�Xo$.75S��ך��Ux����
� �R�����(3����Qo�X���ԔC�+�e��O�q5��P7ޛg�N>n>��.bE�Mƴ�V��*n�Jx7�,�@�f�<�7�+k{o���8{��#bG֘qQ�
����}�vbE6dA�V`"��n?��k�	�}�������@x</����|x�r�+����^���Y֢��<~��U�7	h��y��X px&|ǘ4�I�K@=�����`�%�_������2�N��{��SV�vi+q�����)�\F�A����N��9g�f8��Pr�#ʰ�E������=h��&�L �Y^6�r���ӎ��R$$�)�X#H;��!���4<N��e�S'�.#�6����y�ג�A��aa����fzjZf�O�I(?�φx��h����G�`�o9!vϽ7<�XA�x�"ɥ�æ�4j��	Y�ߏ=çOc�����gX_+/7��6.<4F �b~�7B]k���_�9'��?�/[N��QD}��9^@u,�0%)�ȌBFH�ie�Ӣ[�7��ET< �	�&)6r�ҰQ��JE��;Sa7�ih p*�e�76�������ry�i}!zhC�	ld��������?���:I�GR�YƉ�g��> `M�jM;CA�7����O�� �Z�����
Zb/жv�l��)��*�ҍ�{���?p-$���x���34�[Y^�M�����:����.�����X�e�a�##Z���.*˦f��׊�����:�%k�{��so�{1�dϢ�m�9�/UR ��b[N9@no�ȍ�DC ֠ѧ�Jg�K�-O�*�m>�\v��qO��a��V���6 l0/�~�\/��#��}@kk���8�����r?�y�u��Վ2��e�CTG(}�`�ã���s(_I�&�K"��� U�&��.c��?�Sߜ��C�7'��v���S3:�K���$�q�ۆ�����"������1�nB�L���V��)�j���s�3|�����q4C���m7D	�H�?p�nC��r�x�R*pξ����D�/,�+�BJ˫k�>���<5��jH�~H�m3`�g?k��5�}�#���~�M#�}'w<7P�1�y�@��Q�b�ZZ�P��T���|�qU��{�=����'W�^s�U%�	L��8��7��|�2�%819N�ȣ%-
��8,Ԅ.�g�'���U�G̣1w;���Ӡ��O�����>*��R=�Ǌ�ဠ��������.i�	��>�'���g<��3g�ʵ�/P�ج�n�655�,�Qz�2��u�8d����1�g�)�m�J��B��K� ��!+*!GG� �.SB��C!�׶��z�x�)�Q9w�I����|� �=�l6�?����]9w�ܿ{W>��C��ӐԿ�˿�_w>�� �XM`,��M���MJ产���ףv�x�z�~�"�^j��

�������>瀬���\tH vccӭ�m|4�z�)����A�o�/����g!Ij�E-6�{�L�ݨ�}v���I���o��`����sV�^v��Ԫ�6��,�T@^>'�iy���Р���drrʭ�ivfp�n�.�1� J��F�jT��_��<"���p��8��l�M�t�'p�20�O3����}�Z��i2M"H5<�^��7��ҁO���;�X8�*�^�4'��~q>��A֠v[Θ�G� ��^a��$yom�{̢�����xb6"J&�I ���0��ka*��1��Sw@�ɾN�0��iU��Av� A}%��R��t�2�u��!�������j� �'~/z�ދ՚��pa΍�7 "�t����x��{78��r��A��v��Z[��;=N��>�
���M?)w|����j�p�*IH��:�ߪS��u�p���ޚ8�����b�����0����$eQOv�Nr�W�uĊ��܏�ꩱ�a�ۈb@&n���AFC�t���#)*���{���N\���6�RL(H¬��Bq�>֞,-�x>J�
���WFL������u�����0nw�V~� �9kָ��P  k����b{C@����O-2�e�b4/a��@�rZ$G���a)��ȵ++,/4�DJ�������^;��\�r��,�n�r�����/��+����$[gN���y�qA{d�դ�)��'��W[��iTaR-�4����'��{s_�>��g�X�g���T�P����wv	\�Mf.ș�ڑ���x>%.�?$�hʍÿ��i�! ''Py� �;2?��15
<C__��+w����S��L��*+�zQ��_�ǩ��]ǛÙ]Ʈ�#ZI�-[ۛ���N8�� �k��+�_~Y��+��������]�|������d�P�	Q4� �
_P9�P|�v�d�T@9 t�y��ζ�S� &u'"ř�h�D��J��.!��A9%��~�d�*���T�� r�^
��P�T\���Zy��>�Y�^��ѵ��Ƀ�Tࡪ�\�� �BM���Z�ڴ���G��ѿ?�J\���g濌=�I��TbS"�tr��V:@<� 6�D���G�.���m6k���\�|q��Kr���!�*��vfOu�9M��9��̊�e�e����u�&\IHDN��#�<�s�1E���ܣT!�``<ʅ�y�� `�19=�����\�~���y��d�yq�������Okl��n�!O���[0d�HyS��mĄ�O?"��m|^\����zS�k[nM�Y�q{|���@���w�NN���
-M�C���H��B�� �
p�9���0l�f��y1>�y���+y<�
�a�jϧ���=&�B���x���8nAZI<J�`@Q���T�BO��];�-��p�_g9�_�~.N�_�vMΜ٭�M��ܺs�ų���o��d��G�XQ��1g �߻�P�W�,=~$��[듉�	.��ki�T���H_^E�	ZY��p�ԅ��"Kyي�_}�V"2?�0i(-g�p^�M^U/G�� ��4����{�ꫯ��/��������S����ؕ�}%΂|7��(����j@]�Ã��e5��{*5d�X�5�.�V��6�>7�4��y��a3���S? ��҅BM�i�^�O�CoU]׻�^~P'�95}��u��R¸�޽s�Yhi�|�����`�����;ri�-��7oʆ�����?�ɳ�3�[�"�B��#i��Z��e���qI��I�}����Tm�d,��->�%c-=����Å��dq������)�;�g��� ��U����
��١7��� d�ȪkK���z�n������/C#�$���<�����j����=l�]�!t�!o*�����<?w���yDj|xaP Ď�i�W��mc�9B*��o���R�[ ��Kc�!��|LL��ZS	�\s�)�f��)H�ߘ�@�DۤQ׹3V���U�-d�IA����Q���X���k�s��h=�*#���[o���8=�<b_tc�կ�"�����hC&�(y�5Z��9lΟ;K �j7�����f��p��ݣ��9YH J���3/�4Ԕtdq�����Η31� �m<(��
���O����{λ�h�^��#�|���h�aO�����Y�:Ez7����b��^,������k��b?��A>�u[l�w��t?bC�{���$�?qW^��}7�K�N��y��t���ގ��1"L��=3>�̹�4k�D�	���:��ֹ3x�6��{5�TG11�� Mf�� ��jik���,�������E ~�s�(l����^M�Ă���m(Y&wu1�LL��$ ޾y[�Nqomnȵ����PA����"���?�+3���\�*�Ct���l9��G���*3%�ٓJCf$ϱJE��z��Z;t��Y8�Ҟ�ݦ��4��BKm����ܙ��3�)�$���y0r�*VS�ꠘ�� Y�}�؂G�K�_��_z��}���!��Ȕ�s
dbl��Yd!�[���ȑU"(�2��Gzu�3^|34�7+��K���TJ�<<-���^���hF�D��h�TA��:`��1�3 ��N�XY��T�/���|�7�+ׯ^�N�}��M�}�������3$��W��:�7���N�`N����]����B�rP���/�^��(0��� hlxl-p�*���S}1N��f圳�A�\Xx@��@���~owK޻���}������D����u��� �@ݏ�������LTsM�ڢ%M�k�E�ھ˷�
�����Gڹ���s��R
³L!�u�(�c�s����s$/�S�>T����~�xQ>��C�_��O3�y��cxy�QKR�^X����!��{k����GU�0��x�6�4z1��!Dan�x祙:��������ӕ�NN,�)�5���R�������}�!�_�={��9�4�j�\�|I��]�1��)�	�{˻��$� 1��$Z+_�J������Z|MCs5�wO��ɽ<樶�P�e�<�݅a�B����5������pt��W�: 2�F��w�*Wdfv��sn�����%zsPEr���̭vb�7.�Y���-��,�g� -���l��%|O��=�c��lNY�`eiխ�L�'�ddt\F���~�e �<���:�x������	X���!D��޻�&�;��c�VB�����c�YS�-Ĭ���S֐��^�v���0��½r�jN�Nkȸ�K��
��>�;�,��z���o�����_��$^�ȳ:�+�-�ѡ~933�6�v��y;?����N�Cn8ko�}=|��-&4��[���`nX+�p���Z���y+i+2Z�n���г �/���oܩK
}�[�+����^-�Uk�ق�z���ʛ��q�'�ff�ɓey���
.^� _~�+�X2����`6�8  L990��n�Uo-�i=؊�<0cᴬ�*���Y5 qM�E=�T���Vm!b�i?��9C5
Jn�����5��XH�Wb�6I�'-<zDF?keu]^z�e���S�<|(���[2�?x�@p����5����"�BZ+�j����q�$=�{�{Vg��E��X�Z�R��g=:x��S�^�%�͛94<"�Ο�W�r�D�~�ۚ��5b֦{HTdEC�'��ܚ8�}3<:�_����r��}�PL�69����؏��r��������CV�V�*=�v;g�ԟ_��m����>_��M9}�<	��g!o
���wޑ��|o$m����VO����.̱��!)bxd� ��	j�h1gEex)ю�y*�� ��(ѷ�K�b�ʇפZx����i�y8Mg9��K9v�$����R���������k�b�8兽�>������0�X�g6�t�����(�VIh$�}�B6k�Y��ECx�����S�C�K��ƽߓR6�\�Y@2|O�j��ez[��>99�Tv|!b�:�w>�)wnܖ��5YFy�{e}{�{^R�U��)���AO�N��X�)m�� ���eq�E$��ߕ
8?�ޗȶ�%d� ^��.Q.��nSF�el�@&�����;~���{os� ��Y^�A���cV�)��$8��<���s�#����	�2.^�c(�FujF���jN�M�(:)� ���j	#t��"8�b�D�G����y�����>�
@�3S�\�z�ĨOn}"�n� �5i�Do9�v}��D�Vj�΀�@%���ϝ9@���Z�@3z(�-�/���\�0ܤ���N�]�ʧ�bW�.��O��5 #��&�QbY�!"w��UV�De`�p{�Yf~g������A���OX� ���`�a6n�P|��Ad�ԝ�a9�1"�N�~*�
!�&�ШZl6#�b�R$�,�6*0���U0���4�Nۮ7��7_����.� w;~��Y#��̏���!5���?�7>qϹA���v��M2!lA���H�XK�;3�l��V�/֝_p�$�G�Y�虅�_8��"A�HX~]`]afL 4}�=�)�q
�(?�����%	�Tw>@$�zr"���� o��>��XVS�<���\�0a��p���:79�N���-bj%0����	��C7��[��������*�}�����YH����<0࿬���6��9����ե5�0#|fY86�:���Rz�vv�l����Pqk}���:�v�8��~���Et6�z���?����d�g�b���3M�1)� �H!G�>�c��/����2��6���=�_��1�k ,�Xc�<|8�kt퐇46>ʄ���p.9{i%��Pl4�p2�c�K5�^Ӌ��X9
k��\*��ڧ�}���P�4��<Y���4�T̐K�_{_�$�q��YK/�a@+	��(Q�)�J�#�`�a;��_�,_J�|%R�j� �:��,�Uu���9Y�=3 @��>c�Y�k��<��� �u�ʫ~�ˉ�]`��{靿�d����s�������ח,:	HwcZ/p�s���S��	�t!��$��  ;KIDAT����A��t�������muO���˒��b�����;��8%�w��ð}g'��+���\���'�7���i��P,�F+�z-��\��X��Q�5ߠ�}Sy��UA�T��ׇVc69<tD<o�KRd-K��,�d�m݁A"�gZkY�,�Su�53 `$x��;�у�D��p��k�o�8���?����;��ޣ��Q��݇� g�Z"q4��&�c��9��Rʹ��%�[R7���}x)�4͝G��D��D�4����(��^����=y#C��s�G�I�ٖ��;qiA��Yf�c�P���:g�=l s0�㝬ol������E��7X�����V͹/q61��4�"���}!�t;|�sټ$�O4�$L�`M�������e�u3���i�]��6�)\w��^)e!_�xI����ް
���m&mᗿ�U��ʕ���������;����3��e��ƙ�0I������~Ź��������t?h�XD���i��8��}�E,i���~^e��Y7%�s$���0�� )� !i��$:L� �G3�@��(ȇ뭧��p�.]yx�Ǉ�£��a����˂�r�J
��L�B������i$�:�M*Э����j����h.ZX���V
��HX�4��牸|��k�fP� 5J�I슂qx&f��`i��҆�=k��E�b~���Lc�qv+����m�J�H7y-JU��a}��0�s���mEB�`�>U|����,I�r�Y�!�r�]Ey�i��;w�Q~�"���π��k׮%�Mk����ة iE6X4�������V�:��Zbgq@Q\�/��v5��q���@�L��D��
�@^v!�������' �k��kӥK�Y
�?��nx��	$b�>E҇��d��%�2c�/���VKEf-�,����@Ad���x��D���lu�i���u���*B��Ҝ����;�$� ��_����z#(gR��J�n�m�0�6��[~��]A��P�XK�"'Fwj����⹓�F�X��_8�@NQ�bv���vꆁ1���k��eS��B~���[�i��'�������K��
R}>�Lr`%�3�5DL�!3*�m��C ���puI �bU�k)�eAuL,{�A�Q�P{���Bk�療�UT-�A`��
5MC3�Ԗ΅WJ��V����E�US����]��<��{��@p��5�w���a ��������/���U����Z��/�6sBr�7��Z\��޷Ƕ�!Qsj3X��C`*�Γ���^ǫ����*"�?�Ldb2���]�p�ni|��<�#H����4̆��M���%��!�	&b��K#��W���V4(:�\x�}�\��G�~%K��d��#�Ht_�*jJ�זu��Kq4����M4�B�"ag�0���6ѐ�
U��5c]�^LB�4�����4�=[M����x� ΐ�Yΰ�+>(*E%���St��B|?��5�
Ǜ#q�H}�/��;��1QB-2)�E[����ߦ��=G���p�Z_�~��=���6�'�a�~eeK	z,�r�î`������=������೯�X�y^��R*l`�r��
YI5f����{K�z�WqLz���Bf�A�6$����˩n��	�?N���a�X���9�OЅ���Ŗ�B���P��x[B��f����D��D�hf=�r)<���"^F��QR9"-���_��<��`�r�U&C��_��9iZ�Ozz�O�8����ܞ��%���f��k�b �=��+���]���������������N���ã\����i�{����P�##�S��6��6�=��y�����6�XS�k͖M�C0��6[���@d�xS��2e�l�;��M�{b{B
[����j98��wss�3%5�� d�m�t�۰�QbO����8�)@�O?Z|�;vegу���jS(@tT��֬��������0�$yv�W���$��UQ2��c�({9��>�g�?3�;�jp�^G����|m	WX�eFk����P�~��e��XҎL&ېl�� �W�E·�n_�.�|��&����w��wѝ#����!zI��2E@�=5���\�*�K"F���7�o�8t|<p�(#�����s�Ig��a=��,�%)��ϵ�ƈ�2G�eL\��x2q�X�YHd�߃�v>�,��r	J��tFd���E�����O�ӈҺX�� v69߉�A�j�������d���`�|{�~���c�-l ���l6	�����R�m֊ь�͑�{o�,RۀCw�'\t.un�ڹq�.�0B';�9)�(��(��;��F^�Cw�\g/�ƴKy������9�v���m��\�\��v�W��5�.T
�K*V\��o	���d8=uI�dp��"Rand�$$�-�?!z�z�scB?0��ko�VXq�����0ǂ���W�i��,EZ�)�������4Μb����1�:��>��Nt8k\h����)����'4��7`������{p�P��Ik~;K:�m��I�C?�H��ĝo�#��,���]�k����W�ww1|�72��͢Ö���be�"�KP_�U�P-��I��Vb�h�:3/�ˉv��{��_���x��	7���`���85�����T8�i�L���-x�]*�o�H��]&�%��{L��;
���]j���Y���R9�L�:`"9:BAW>��.��P~�([��;L��a).P��/�c�;�`&�K�n��dk� s]\�>gP,<�����I�Q0��Y��FbLOZpF��Ap�Wj܎g8j�(�����\��*�������z�~!j�.LY?�������0:�yք�j�L�v���:B/��"7![��ig���*�))X}�<^[��ɿ�>�*\<�$�QK�cX���ݟ��4�
;K�� ��
T��==�Rix�k6�t�뒕Ы���l]�Y���ٞ<�Ō�b=�mF=X�A�8M����@&`�%�e͐�u��I��9��OK����VZ��5��Q$Φ��A�^e�d�p��AV-<���N��M0v���x��#w���d-���udz��N�W�2�=���Q gl�6���m���A�aA=zznVA,�\\z�: �tg�ɖ�5�vh�R]�'�v奻��&�M���<��2�NȌ;�/��F�BLz�TZߨkc���&B�������,��
a���y���S��Y*�6)��~0��}��3Hc'q֕���U����K憛I��bw�*�w񷽟c�j3Z�@���y�_���m�KT�%yvWjm�0e�XA���.�OB��CX�������W.e"	M�3:&j=7��:8�3q������&���B�q����`�������^r�>���0$��P�G�ģɅ���~V0Lv�̜�h|��x�@E��|X?_���0�,6a��[�Ն�뺙���}ʒ|hO��&�M8oF�������@�~o�矐E�E><�M# ԕ�����D��TRy��=g�{����x� .9����gnh�	|��L��:�).g�=C��HSUr$ �a	N����P���L��!��qT~��n�P�`M�;xP�
�K2g+lV"m'L�>�@���Q��2�NE�j[m.q��X�uU�VS�߶A�X���U��?a,�fc�Nق�A��$�
R��|Ӿg԰%�oiZH#�����,J�������	?�P��eYo[dCX@��62�7�y�� ͺ)�t�-+y/�)z��+c�W=τ@�sP�	�1����$ț�h�����S7 �p烀� �'�=��^�����F�}���<V~H��HU�)����bAm�P�&w�яO.�NL��g��L�ݲ$/�Y�8F�Q�+$^�W�BAo
QY7�I�܈XR�}��[J񆀏u�F�_a�N�Q���d$	��3u���>o��qR��8[���x�[�urG|����9Ƙ�j�GrV�G�x�i��K0�>��@�u�J{���%N�Js�aV�vL�M��o� ��)�¿���xr/�^����Q}�2��� ��V����Z�$�lOwZ|S,+U� u�SF*<�
C)�Z�����Ή���T�f�n`�N��b,� *?؜�.I��w:P��_@�٠��Ui�?��[`����#�/���<�h�<�#(k��.�]�uJX9�(���� ��"_m��xx��O����B��.q{�r�߯]�-q�K�4�oN>]aZ!�҅����BTOL��d��酎1k��ef��|�$�������ZP���cA�>[���}��X�&�̋�\��/Tҡ\�=�H�d#P��T�e��d-r>��N�L�"�c}5	�5u�RO-�{�U�;d�\$F�>��Q讇�S��Qa������}E�;	'�8;JJ���)o�ֿ�&�E�D;�x)����qE����ʄ|��Z4�^-s�-�	��d�&����j�XD'�S}F����Di�!�bL&�#4�U$�u�Q���ʳ�Sj��S�E"������C�c��L=E�������¥ak�h~���V@_%���>S��PI(����!���u���J�c�IE�Xu`^Գ!%%���4�Ӧ�Ѵ�Tk���y���Ac҉k,b���ʓ v�����h����;-�R,�&�`x�+n�UI�"�A����tx�/�Ƕ�m7��(6޾�����.-�d&�`R�:�B�~x�آ�|�#��:]˙6`��2V�����W_��A�|Sl�S�G7o�c�z��s��NE��|=�3T{�DM!�I�a�>���N��c��$��p�9��cjͼ�8KˢB ~�����ԐA�&�J��}d<���n����Ks�r�q��iD<}�],�� �pb��0 "��v�%Sy�l,�����0��QH��?�VԘ���ae����]{"\/2�%��(?`O�1�~��%�C���SQ�;I�5�y���ӝ�lے��⢛���ByH7������b�G��1���M��<5a�(k�3��j��M�Þ�.��v�����sC]��}��+/���i���9$V�Cm�����xlD#�B�D�y@�C"�#W�-l�D]�Hz5�r���SjzU�=J��"wnO#R�"���	���ZЧ
n�y�B�M�40n�ejxʥ���%چ�(��'�<an��=m����5b��G��X<G���K���܃���׭���*�Ti=n���$#�AJË�5�J��l+��uo��dll���A/>o��sL$F$y=G1�v�9<=|UK�)�VK�C��o^c8g�O���ԟ�"�ٶ������h$�}a�E�jw0g��$l�9��CHH�Y?�����s�5��
³a[=��z����ȥu�O'��g]N=L5� ���y-�U�R��i�L���ˤǆV������SN�85��T�n�t)����$����Yܴ�-����������I���u��1����n�6�6�G�y�Gd�]��O?�u}j����?�Uz^U0!W!�9&���9��,OIxw�fB#&ri�9�9٨+� ��i�X͢��G>i~߁�0��"�Y&�K'�7�͂�vscw|h�����u�_<�	��z�WU��+��?q��\�ƚHy����+N��V�,�=g�{���+������V/�"���%���O�J�y�P�|P�f$Ѓ�V�O�9Ɍ8r%���̐P}�5@1��{�N��L��{�d\ ;p�Q�+�������~��9��*�[�`��U_tǮ{E���r%T5(^�v�(-uv�G��� �����بbYDc#�LX�PQ�"���u��j�s��b��m�Ie\$%[&�@����3��lA�&�*�qT.А�J���W��b� ��aJDY5�)�R� �h�Z4� +�ti�ul���ځP=x�;��� ���WG����0�g��+R*iF�H������+��ೄ�I(�p�Ɋ���aqFY� 0��
8w���H��\��m�/+2�-��p��^�C���r��_������YU��ߧ�L5���=�l�l�L8Ip�����Ͽ�:��Yt4�˦���QG��C�,����xgV�˦qrw^a�,|V�r�4�l������x�qi���hJ>���O�@c�^\ˬ��_Z�q��K��!��s3۔�O�g��+�o�g4���}H�6eH[=�p<�b5D%�>I��G-�Fd{��6�ӧbx�� F�%$�f��<o����B�H�T�)���` �3,�	�eR�l|E��Z��dG�\�l���?r����R�]oQԖ��(I�%�7C-m�#����	u�pjiP��mV5קLQ
�K��c��:n�n����f�eCq�a*���+�����J1�*�w�j��6��|ZX�o&��+ Y�y*��p=�P/�f]��ߒ�Z�" G��A���n}�����'[ß�V'AƳ��
�?����aߘ��?�OR"`R0�������:ʦ7'z�X�d�(��e8��h m��j?E�2��s�v�[FB�}m�yeB��gb�ǘ������"��|�	wD��-oqJdͯ��(��]CI�jH��F@c�S:r��>�:�r4�mH`�(Ȩ���K�.u�E�2��>4&~�ZG^%}X��@0"��]<���|(k߯��>�ݺIn� �7(\̡`�,?�����2����`U�x��yr�$+\�w͓��r�w�JZm!'�a�)�` ��y���?��E)'����k|`*��Z�_���Ϩ�؇pgP����_}�#����\�{O����%_J��@m��`�����:�=MS���]�>M�p�yS��z��.�X��6!T�J��
���Dx¨@���=_<[iN+[��` #��r��'�}�|�NYD#_���+��Z�6˃m���i�m[�/�D1GL8�e�>�^��j&X�fB.�GP��'קb�Cd�n�Y$8��rK���ɮ:�?f�&�tg���l��0Vy��V`R��pS��J�nQ.S��i*N _rbҴ��~�!���ɼ��)�b����Q���δ�zMb�T?��&������ꩠ����.1��i�?����q��y�~u?[����
���Y��'#� V1������!��]2R(��SM�7�Mw����5��,hxKq�	,2���t�~&�43��%���J�����qT�a��(��p\��7�9P������t`������dZ4���FA{?�o���m�E�E �R��L�(o�C#SK�����h�9�
GEw�?�kKD��kXd65�	-vL��6���ڿY$��d$�J��3}��K����p��\��wqMxB��^e[��*�"+�慅�h�`����7��Bu�H��=��w˞�"��cz��l��ѝY�q!7>�?�Q!�X��6a�9��L�t�W�l��U��q��^�?��m��S4�� F��#W�%�k�(QS��Ҫ�hM���A��)���[�GƬX�ˈ+��l��$E'Hb�/�ɚ�H�^X���:yȌ�N����MN�ﳿ�*M�ʹt,��s��F,������Qz~6Z�V�����k#b4a2���:���6�q&�8#�S!ْ�h�6f�b(R��Z��[h��M
��:�q.��>QS�!��n'k�E�(����b�/
5l!��
�!�'����ѧ��e���.�I@]��jz"�b0A���s�}��>&pY'	�7́*�w�'��(�<�a.D����hYI�FS��tZU�D6��`x`c#@>F�E���a!QH�餳I��l�	^��:&�*P(�t��{���8>{S�#��+|gE�_���e=�W G&%N{tQJ����j��Ћ���I΀N=D>�#i�X�8۹ؤm3�=����W�#)g��ƜL�������;kP�᪺��FƐ���[�_�t��،����[������pG��ĥش}�'��p�:��6ՙ�)4M��T
�?�Gf�cbJ
�4z������:�΄X�e��-�Z����zi޺��rG=E��c�i"���˵~^F�c$��_�ɥ`N����|�WFCB;�R�ce��]�+��$X�%cZ�(���zs��G�&�
�%w���P�+e�qGۿk&A��.F9���(�:X����#�9��$9��R�Crg�(y��q�M]Y�kA���������<)=^���ub#�a����jV�O�d+���ח�Y�VeW�K�{���h�����z�2�=N��P%�)��*�(�V����>�e�7�/��.y@o!���fM���(��XƲ��i��=i�8]e�u(��ڬ��V��D�2�X��>�5vD�����)zU�6(������nB7���s�ީ� 23������(֊�� FXԷt'�Ⱥ��T��Ό>)hN�ER���&��+��⎉'1%�F�Úe� +W��&6c�_�<�����תflX�ٲP�1E>���w�f��~)/�89>�"� �]��%�:F{+ŊҌbn�GV�Vk�X��I�ܼtzB��@����Z.�	ko{e#���GHnWbM~��|9mf1.O7�YT��	s��L<��4��;u1�Je�2ۡʺz^��R���K��"�3�܄yN^��x�O �b��zeԜ��S#n�4�U#GH��`��P�o��80�k&ݴP�QYr9��wZ���KM��xNB�e��S��Oɳ�<4�i��i�������UW䄴�<��ȕ�蠢O�G ɠ����l�a_2�\xU3ġ^����1&�"�4�����[8��(k�M�[�K����=�xGjK��~�1��.�� ik�P�@JQ�W"���t:�,�q"AA	|P��x�ey킓�H|�R��J8Q W���g��-y������L]�B���_Q�4����X?���N0[��^��n`�Bn��-{�.|lhPXZJmj[�#�wwAv�����R	��a�b8r�-	�P�t:�J���T��j|�om?�s,D��5�Pb��h*�O��pd5��=��&��4��}���n�z�4MH$��<jr�d�ܹ�\ԋ����E7���Q�����[j�����J(K�$����*�rL���enٶ�鿱��~NH��=	����}����|�pk��#�S�^Ƌ�}�?!���O��9�	�0V��X*<�|�R��־ߦ�l���p��J2%�2�]���� m�j�-ַUaXkb�-��=K{Z�aa Z��f����]f݉Z1r�����vV-ԉk��ZF�f�+��6���:r��7^=����,�(��i�!�7z��k��%=�$����iU,@,6���R�VjQ H��IUV�]��h�zӰ��(�C�l1T��&�'b-c�^�s�<b�̪��0FZ�o!8��bS+�B���HO��g^�qY��ڙ%~�H(�L��a�:����R:P�>�+ĭX<��cv��ZƀR����5\H��;7O���ϑ�"���󺬽EYJ����:5��H����n���s���K�����4��d�s'�|;��$MW�T�J����0d
wv(�RK�&�cb��~�hPc@����P�V"輟 !-�e��>�-P���֦���*�;n�I����R[�V:5�ň����q����.;&�Q�jܿi�`� Vr��|�R������L��(�W#%�Q���3��)���̖]�&7̅�|1 ���d2h��z��M-��A�~fhVtvNE�=���z:W�e���ʜ4�=�M�YP�<����:�Ysϰ���hV�Ufu��j^4��!�h��	B8�[��wː��"f���-`4��r�Ncp[TN5)ZVJ�4.��A��d�D#�7�͍�{�8b3�	�0��2fê/#p�U�/�b�u��T�Y���A�������m�"�e��6 @��7�0���[�k��ʁ�A��&^O{�D����rF� ����l��.k��(�`��#/��J�d��pP����3iX�K��qB,��S�U�����\*��@<�پ) V������cA�B��r
�*��� ���/@�+�b��O?���t��[a����E�3�k��H�D��y��$���ijf]��$+~w
�����x-9�����@�oh�`�	j�����w�Y����kZJ?�$ջ勐3���i��^e\>��z��U|���r�$J��n'�4XPc� �:���h�`M����{�e��I��0�d��9�X	���n����.���hi�2-P�YiW�W۸��n���Jʫx��;)q8��c�7������z�o'�0��3G����{������:�t��J$]�1�����Z*���S�a��7RԽ$�w���[���σ���:h5�&Hr�	_�*r5�-���$�S� R�k��҂�������{�0��8͆\=��EHQ2�D�kL*��Xw���6I��l�)�M)��㙜��J�h@`���6p'/�Cli�sW��m7ҟOH�M���T���eͤ�*��D�F+�"j">�~��i�N�9��l"oǖH�٥a�n���-!���j��{!cA�m
��'\�(/�ڍx�iK�ϣ���?�)�1���w7(&�}�"[<M�EuǑ�VW�4+��t��}���L�$����k�����|����Nt�t����$�:Ş&j4:!/�D�����l <e�	 �<�ӏiHv��ͬM4�E ��7�N��>�9��5(��{��v��-Ouq8yi���y����?�g���B+�@� S]�X�͘5']�e��P��H+|Ͻ�����R�@
��)�0��dtE���d�o��%�÷�f�r0���~I�+1�������Zi����j��,>�(1��tkQY��ߗA.kS�6�}��*����#�_�+Re��D:ǂ��<	�H�,?��it$���x�f��4����%�ĸ����/լv�%-j������eƯ%�go��\�c1������9!�\���h���4����q���PY��q��e�l�Xo-K`A������EJ-�c�&���
�/�`�szV�CAq}`�=	��Z�#$�WIK����ˁ���XydVK�ZB�(��ާT�%�P��M�䓆�B<�~�a%NTu���ZD�/�]�����o�u�r��
*\ֆ}0	�����?�$�04�D�cJQEV����6�g0.�T��TWۅY)H�L�H�f���F c3&i䕩F�آ �-�5�����~��(O�G���n�=��]vX?gZa��+o�Tcxv�tN����TK�b��2`���zw'�#lka����(�����7��2g��g���K�6��-:J{�'S�0�P�|�EGj��["�1����`�h8�r	�<�\��X8+g�Q���u��5�;��P�¡�%��1�����o,s+'D Y7�d���1;�|�vY�9�wMg�+|��n�3�P��k[��G&�����E�Ld�γ"V�й����C{�8& �� dhpyu�Ҳ���`�]��B ���l��Ƅ�OX�m���V�5��:�:�"�q΄����yN=�4���O|Ί�mf�v��Cq�m��
K��MC^H�\8�C��~�O��TS�3$j9��N4���u��9���P�#4�ЦǯJ1xl��H��6���ӈ=���bP)��ǹ�b"Ǧd�.i�*o�ÎY��Ps�(
t�	f��zn�D���݂Q�݀�f�!�}��&˺�FT��jn��;�+���!�\�Y���P rw@��1�|�e-�)t�`Z�)4�N�Y�!�i�����h�v ���Y!m���ʊLr��54�ߔ{t�^k����㻐%U-Nno�9l}�������@Wa��T��b&~�8��PF���G�Z�O��497�|�S�Zf�LG���]��Mw=7���Ӣ�8�gm�\V�6���~��P��.B��~/�Β/��9�Ʈ�ʌ%q�d�J�M�S_����ge-��m�պ*ۖMub4m{������J�N�f�=i$�{�r�4p���_�hA���}�{c^U?��w0!�L�+��?Iقf��K����B��|�+�l\E]�%T��ӝA����tG~qt��1쏥0��w�2U\A#��Q��*�
G��r���$gŬ<.3��.�Q�pY��?"3�ȭJc�����N�kW�P3L�u6�NZ���r�_+)<1טem�R�I���g/��0�F��1+��vrH������%*J�+�U���s��9��{N���?+��i��#O�+�K�b)i�pտ	�u+_:��
[9<L���\>tsz�~�}��XT���mԨe���V��`��w/w���	��c3��%��ŭ�QfQ��::c��Qpc��X�:4jT�F�D���T6���U�<��� �=�(��!;�����&��]!�_�q����|�9�U�Y/� H<��ٶF�wT(2�����{ǽbE� ck;���y���$�O5�UU���$Cf4���M��4h8x��|ʳ�B�h��u0W��9Ƀ�Y��rחz��)�����Q�&��߁��Y�Zv1�f��#�N��_ɸ���ƅNm�d�/�?�Xt\}���[v���%&O�J�r��`�6J�j"�Yۿ::��+_ז��W"�cΪ ��a�=����|Qh���v����k�m��-�V�C�����X�z�c8���б��Hۡ~Z�/�-��\�x2��/�?�4^�;���H�<z�t�v{�&{���C�j<T�,��W�:qs����J+�c��d衆�J�� ']"O��y}I;k��^X��}�k:j��ׇy@� )�d�2�)�@�X��ȁS7��x� d �y�����`��T�[Bq��9F�Mg|+e<|Z������OS'j�N�N�ڿ(��@�T��A�X��E�Gq�`��ץ� �8��D���]��s��-�^U�{��?D���ո�y�$(�>�{��z���9��X�I���G=�K�&gV��,Ԇ�y�>uJ�
|(�0�|���W��%FtA����]\�2��G�xXk�U��<���y�\o�$��d]t7���|��8��H[�
2�\?}����du�C�,��|���5�&fۛ�P����d�Cm�����i��7�Q	��a/H:�C($����cDT��%� r��U�t�!����2�������j���#e�o��_2?��߉�BQ�Bgoh�RN��[�?���ύ=Ӟ1�8S��릉E}O?����[7��	��c��3cNن��G�vYX�%�h�����Y�0�����̉�<�4�E��V�b?:��|�ޟ�|�C��{�U�<��ѻό������E�|p}�$��2�|��T?������"��%
�=�Cu�y2��ޝ�0�!�����j�8�{=:�]<�X��� �}���O��lY}\f�|�[�OE�&�ͦ�v�Vݜ!s�;t�@.�p�Og���`Ӌ���)eL�RrΖ��JS��jt�xt�>g߲]��@c�͹���y�Kuq�w�Ew�y'Wm���Jc'}�;�A=0����k���{YڿI�������:�.�RQ|@���s����B�}���s#]i�>I���%��ڕd��A��s�������o=���:�mp�� �R4y����H%�z&/l�Z+ �
'����	�"�\�A��j�߻�O��%$]LG�7+(QRҕ
�t?��~��;�?����X�$&�ÃSW�e>xoy=d�
{�ڞ�ߘ��>}:K�ܻ�<�"o)�;�u����,[�����ج��1�2|�L�'H�;��o��gS^�����J߂�ϙ�.��ŭ<U�3M�Y�OF���%���̢'@F~�I�}��wյ͓�>�C�.#7�[���q4a~C�����	A��ġ����D����`�[��8�Q��H�����c������g��6��k�.�-e�f�*ɉ�#��7w����q	ʟ�=E�[dK.ʔX?;
�Oٟ�IM�I0�f5gHS"���W�1�c�=:�x�{�8�G����'O����9'VqM���\�)əZ5ڷ��vm�\���}��$��-��0��iپ*�B��X�rI��r�ֈ-��Iqf__Ԫ�fA���n��	Ta��;�D$L��d��%���V��=���^<�F�ϡ9������cQMsY���T�f+�r�㘠⒁��"�l��g��t q�<�4v#�!��1K��#[���G��.��_!�l��Q�����w�Xﶉ��A��,k��U�ME�|]J^E~_6��'dUro�����^U���t?�sz��	I��Y���q=>e�m��������[y�DMݾ��������u�T1y
�ɦ�vz%1�3�Ԗ0�|;�|���2_�Ek����#>�ݜ�e��\6�-}D=fmH1����:��������8h�8�W��nn�W)t���w�469 ����0�<�Ǭ��9�p�����D�������SӲp�����S��*R� �� PK   ��xX��MY��  �  /   images/6959c78f-01fd-4792-b095-b0ffc5233e8e.pngtzUT]�n �`	�ww�����mp��n	Npww��apܹ���xzu��^{�쒯���P ��O�>��H�+���qm"�}��Q	���!:Hk:��#����$&���GF\�0�4ޛ`��P�~/�������B4�I`�&������n��]�9"� 6�E�|ڑ
���
Ǹl��:�$�5e�m4���>7^?�9vJ�_��a?[�BCCv�!Dٲ�"s���#�6�Ķ� �5��Q��ߙ�0�o/lF߶�&�V�PP�<lxk�ylO,����i� =�0�#�!��yU���T��gBy�zΐ�
�X�N��]�#h3�5�\�񶼷�b�l��`��� ��
���v��r�Yՠ�#���O�S�L���!�i�%f�6sB���y} >�Xǔ��C^�e̜�۹e�R[��8��bT3����4(�V���������WId�RPɒ����%�* Yr:k���H��`�A2�N_�8i��/�9��J���#dI���%.�~�bA�t��B%�/!7f���q�!(�/���Y�ǥ�"��p8=5=�*5u�ʠ�2��q�$g� �� E�Y%��2�L��8G`�$�:[Q���NP��E@(d'߂�wr��#��WDhP_ͰMܸ�B�>`b
3�WnB�_�?�3��&�����E6�N�7af�,^B�"��f�W��&w���$�F�L�[z�����YJ�;]�k� �9,A,Ta`�F�ot�i�m{_ȟј���(�?�ͅ�^˷mYa�t����b�9<:-"���G4�%h]�($D	�hoB&�������/'����3�?��ޚbI��6��;���1 D�$�r@,���r���c$~�30\���$���C��8�X�p�i��u3hK
9�;�e4�Y��)�<�����_ ���;�w4}�����2�q#�4�$j��7�՗���}�bK�}�p��}ZX���/F�fJD����Yg�g;�r)8>MȜ�B9=?48�����v�
�)��V�9��߽_����C�׫� ��e���Nû]���K�S�i�D.��9�߹w.D��3�1�u�,�GS6I�6�ڪ�1��z���2+?d.X)�+�'S�	N��M�"��ú�_)+?��w���IEP�5`���-zM�BQ��jl�#�Hf�\!�|}ڲ�:�藀%]�D¯@M�(��i!Ĺ��U���:�:���U���L����Q����XI���ղ�����s��!���Z�9��wܷ�[\tTu
&>\�W0���,��QP��s��L���^�;"y�3����O8�3��������j;o&7��jw�R8M��%�d2���F
]�Oe&n� ګ��C��]&ڐ���&�NrCg�`}Xy�X�&��#��9�/��j�Rc�v1�����!�?/���ک�����͖��^g���~ѣ���~hm��^/��t'Z<i�ef�y�ˊ%�����)�dlK��)F���d:��q)�?�'ݿ\�\�Gon�dba0�$wyݢzW�{(��G4��d(���=d�'��ɜBcebB���Yju���LY��s�4ڮ���N
3O�2�ے��w�Fܟg����J�¸�I�4o��H�+��u���9_5M��`�L+�j���7�"`�������w��蓻�lT��iJ��h��Q�vaP/,9Α�Dq�:���YI�v��ƨۭ��;/X�+�}^|�c�9��L\c}�;c6�hh�^O�Y=�Lh�G��Hx���a)�����{p���:6Kݏ�/���5���e�Vc7��|;ܸ{��k�ϞN���7iA�!+�[I�؍�o0�Ũ�ϖ����4^�\45 �cS	�@�F��uf��>Ve��j��D�Z�>h���r��:����&����/ʍ����8���g��۞���3\5��u'<�aG��r��5�IV���(�Q{�+\<M���ׯ_-ll���^!�Xr�/�רk��9�O�_�S�#R�˿:������n���EY����4)|��K���i��bs����6�|�y��5�m�x6���÷ۏu�J5O���_?�J`5dƨ/��1�D�ғ��|�#R4<��E�~�F�LJ�P�����B�}ك}��.�K,Q��	P.�|9v|>k�M
���NrEڶ?mq�1o��m�=/��s�i}q�Ѕ�?����!\�(�Ps
�@�iQ:4IP�������Z�-
���XkAX�k�|�K��Y��o�je��ݿ�g��
gꈾ�}o�����23�����zf�IqJ��/��ֿ��B���z8o0M���oV^i�G�6�"!I�S���g����P��#����hr�����Ϻ���ꂏ�yD���p|cf�˹�s�P(w���!�c]&o!yB���.�}�w��E���F�|^e+�-g2½���c����
Q9�rx�ta4r^�}��� �m�Ԕ������P<y����P|�-''�)���z�K���|��'��6��,9��p�X�wS�UgkZ}����^A��RW�����Ѯ���*�ܞ;�:�0�A6�P���6_/w"�N���ҍ�2}��W��yyw�x����8-���鯚1�È6+sPY%���/x�ץZ��Oz��q#�!0N!�F5�F��_�Q��Q��(�8J��q-4mH�	Sl�;9��X�D�j�5�c-d�䵷g�� !������98���G���bOSш��01��9�=@�[Go��\���@���1eKQ�����i����{ �'��7ѽ��_tb����+��y��iI��Y8����ţ�uژ	h�@�[�aD�	0Zc�r�f�m��a)�x&Ӱ��gt��P[( ���˙��É��D=�A:�h�����K��u�,���Ӻ���u_yzz��mB����lQ���|�+`���5{����TLP[' -[w���ޭ8t$&_sɕ��Π�_�]�gQ����͹܀��C<��F����J�B��c�*����c�?����b3BC�zRنʦ9�{u�\���Z�V�+x��a��+dDf��ᕨn6|;�J{,8=f8,r�4Et֕��;ܽ���Rę�C:8�-b,�8Wf�Ջ��$#�&s��v-�9�R��	 Kw����j�>̔�S,�,5�6{(�P�(�\�Xz��GL��@�?��Zk�7�<4<l�:��������������T����h��1&�|�EWwx<�*���1}w�N}�������m����
y
�����ު�ΰڪ�Ӹ�PU��h
SRv�(�}�N83A�]"���J�誛����i���b�����zzz:����^�~h�#�>�6�P�G���)*��J7f�O�����Q���>8V�|�:�h#���m#�ئ�����Q�l���Jcc;�)g��G\��E���͏�Z�z҈�潶�b{�p�0��W� �<�'������dE6�oq>����/�TH���FN]��R�X$�����&8�	k�[���;[�8���K��~hcͦ�0cy7GhN}�,Z���j��8�ٷ�����㐴�.h/�B��L�]��%(:���_r��1�񀗗*��0��S=���z�]�7�0��İ5翤Z\Z/lI&��{0��#LFZ;�#J֦�V�Y-�Jv�55Gb�3����n�>�϶v�g65��
�J( �ê��	��XO�Ozj�^�klLA|���:�^�� �b��ϑO������>��v� j��q�?�n�"��e���X�8��0�/��V˱��� �Hg�����^q/��ڃ!��� ������[�Ewb{A_�aGd�p�J̑�2?T!�w� I�+�nB-))��>39�g������a��ni�2]�k!���$א�P�8�F�Q/u��N[K��X�=�hd�ܤ=��������e���D�o�.�.\	�{�L7$fjT�%��Bُ�M-��JrT����j�/(��4W��M�U�sD|�o��8�n\i2�F&����3�ug5b��̲�;#1�~��=W�a�;;���T���cu��3��S�d�܀�6Å}�I�x���м.Kh��:�6.
�N��>�#!<�u\Hbd�ٙ٢�𣅄����`M�'}غnޟkd:ct[8l�Fc��q�^tc��Ew.����ģ������k��t�Ce5F�d��y|T~~����B����CN{Y�h�1�P�2�+z,��	L1~�>zR�����;��3u:��7��/�eU�5�s�c��FK�e����ǒ"�ݍ�[��f��H�}��jC��[-�^�T�d��j�}���*�b��2�k-�����-zs��R,1w>�Y_U�ͤ��d�4��ܔ�f-J4�B]KW�����Ա6f��>���ze�<��������aK�d��l�㊶Ɍa�{s6Y͹�]&�$���2O��P��}5L--��I����>�-��n޻�IR��=�h��][�����d�����b�h5�԰���|4mgm%G�Vh��C%�MЃ�x�J�	P�#f�Xy����4�B��Ҏ��RU�P�����~���YK����k�e0�M��A��yq`ۯ����3\��]�v��ҦqX�����Y,���D�OdB�9��9V~
��DC�J�~͠��Nf�Hň�E:��[��b<�[�L�I��B+��S�%I�S�]ed(��c��+V`D䖏N��$퍦�w���$2�͊��5~ŪϮ-@����i�T��@��`<�X�s$dGX�KY2hh���&X��~`�m�NV��Ez;`��T����D(B��|��� Wf,V��}Ã���m�8�JĠ��O_c��ʄ�^�8	=g�%���jw�xB���o�J>(���(��O��ϝu��Y���a�w���7M�L����}�c���B�q�E�VM5x��BCq<�5s8L}�
M�_$�t�MW����Ĳ#��s�$�-̴U�����H���?��Qh�lU!Ę�t)x/+;.~�6N��������<��D��CyEAI`L %t��Y���	}>��zh�zPep�{�ab��U��������0���D�����y7K�<��/&s�f�6�"S]뒅9�h-{�sޞ���,a?!��c������M�6��@��˻ �m�x2�N��c寽�n!Y�t)A�d�rUb���29p�'LZ�o�b�$�.�gn�1Sq:����U���vi�Cҫ�WlB��8J��%�o_ $~T�v�VV:ꪈ�E�AU��^����P�C"4���k���R4��7�(�lk+0-�� OT���Bo"�! ��bt��v�����'���^����R�ܨ8�f�V��w�>�_�WоN#�����8�ڗ>�!ak�b��Gjė��1��	�B~�}��mc���҈;�bG�3/��tT�؇�mps8Mu���{�hһ��}���m���~~�	��I����h�tT����MP�d��n��E��!t˟ޚW� �o��^�Dۨ�6sLtH|>��'���]�=�-,�����`�"���^�F.(��HR�<�#�ԉ^�=E�A� !�q�Z��WML�X��I]r�$C���d:�l�c	��g�|[�:�`$�Y4Һ!H��/2155���7b�PfV=r�t�FI��_���0Mú�O�Z��T�*D���S,S�n%f��ߕ�N�!S,Q�fԖaV	1���i�~��,�2}:O�^��<J�J_� ͒��#t`W�g6�t��X���a]��+2O�$yN���5П��$R�#
qLe�R��;��X�|����R3R�qJ���z��ʐ߿O���d:8�/�������������n�>3�U��l���/V�����>�����;]s�dA�d\�;��^MY���?7O�b�������o�B}NLSS,��>-�p�/������_<��
������+V�#�R.��-D�p���E�C q�ŧV�������b=���Äew`艚�M�����8�^\�����J=�>��%	HP|3��`��u��#82n���}�1�f�;ň� _�S��/�p�;�m�NM[�AZ7���Q�S��޷C��f�Jô�!�x.�����U?�v ����+	���\^E;�_���gӎ7<�"{� R�b�u���E���P>VEY3��kb��o*U��)������ԣ��=z�L�F��8��z��8��}K�G__Q�rշ�~.�	�*fegP�w���*�	�G���F�?������ �U���
8�?�i����Ã��2���')᳸�����nK2w��5��MŃ�+��e���Q�����4�j��*�����t~�B��ة��OE��ӥ���a��bG��Ee�I��v2������эG.|��k���q1#��%l�	�z]�^/��x�q�D_�p�'��C���'�t[�=_��OH1T��{�f���6���_ 	�W�t/�+lj�E�b�)�O�M�U��R�'q��b�ը_{��>��dY,P�!�o�I�4�U��{!��N�
��!�o�bt��n�p�D}���zf�Cj�����28`�e�ZW��j�Ӧ"z�ޱɶp!��%��ސ��R[U��RU޵���#�7\�p���_�u������M��a)cp�ɶ�	={���I������;1�T�#:�}CY�3�8���DL6���ѵ���8��۟ZʢЋ�զ����1~Z�\��#�X�ٽ�!��=2�������S|������͓��V�-���o!��Vi�YW�h"&.��A��'8�%r�.Z(�'�����;��I�:F5�gJC�l?��Y�:���~�V8�U)*�d�a�m6���lO(�����:.ݐ��aք*����Q�	v�e����J}�sm�3�\�L(&�D�+��kR���W�Vd��6���P��N�IR��nr-j�e
��6L�W��zU�����x��,ި���f��r:�-n[q�׮Y����|q-�
��Bl�2${]�X�I����+����i�3�9�W�����L�7-��6	�ǡ���A�0/����y���5�����u��ɓhFH��S�I$���S�j����2�"��K|��z!��������	����o~���9-d_#�k��*�?��$J�S�.:<����q��{Ӻ)��E��������J�݋?�-�|K�UpY�����>S�r:��Zd�}%A��	/�g.�O�O3w��(T������e����:�:��w-�4����W�tÇi ��Bc2dJ����K��I-;j<^�.�f�qr���1���|�.�:V+�����+a������B������ �Sñ��~;YSDa��_pÝ:1Eoث1&|��o$�p�%�_l�&Jv�庠�X_��!]O�܎?# G��mԜ��&F���R@Q
ho%�*qCMys��s�$�Š��f�_�l���6spk	�`���Г{�zt�0ѩ�[���,:�W'lAuw���<ҝ�1<_I��(��z�
�)�2�����9B|�,s����ߏ|��6��x�r=5�h�N��;�!��d=1�fuZ��Хj�\G2��:��ܼT����(?b˳�5�KT�J�\.��)j0s�LY�+)�;���z�,O���Y�[")5�f�ˁˉM
���"tGY�˩t�	n����|�Ҷ��*Uh�D\�rwmq��fc��/s���2���x�T1l���Lh��& $d���ȥ0[�'��:~5J"�����������QaB�����Lc�{�QN���S�͝�G��4�cؖܚ��:M��4A���_:0ѯ�������xlq���0��7��K�_�S0��/��G�a�����Q]6�bEd<������s�~ZM���.���}2�j<�拵���LP]��\���7�!rt�tWy;,#9'ᗗ�����)Df��,�@�7J�d����IVwy��׎����~م��ɛ:���%�ŝ����Zoo�޲\���*C,S���-�R+��S�Mx8B���4VlYp�]R	e����6y���	�㛘v���h�$���Q��Yd|Tx_� 4tCv�\����3(S�c���>z��ٰ�+����`��h鱦�#�o��'��ͪ����6b�Yv��7��'��>Nd�Zy�7�w��a�쮃Vp/���.��i��uə~ �u���ۧ?�V����Ǹ�Qhw'�t�ǆ��f�(G�'����h��ʏ�I�=(ēcq�؈��w%ae�0T�J@�]O��V���ڒl~����S���(�Fv�lf>���_F�l���n-l��f"1��|~2Xs�}�B���B�n�xHٿ�H8
�{�rs�j�����o0=�8�{y�����$��k��hUO=b�M����H�C���#�[N0�&�y��+K'������I��Y���5Ob��
�jb�oQ�`A}�-�9������
i�|R,Gg���PK%�:��oLqж���_��a��~$[� �?5��I��GR-	^�oٖ�\Q����{�|�t��jv�ONHt�m]��T�u-��(^�l~�����U0G�5OK/lE��o�KD�$�����
�w�������]�8��
�Ķ����ҝ���&V�$,[@��E�=�Vi|��m9�T�����9�U	�8����s~�G$�d6�Ͱ�[���֬��c��������P�k��v"����j�>�f�$���ĝ7�1�7��y��N4�_��T 6�ϑ�V������q$Rb�?&g�Nr�ˍ�����2�l�aA^�;�C%8�WH�S�,� ���f{�h���ׇ�-�|�@�e�U�5Cjn6����0'cwd�lp&��|,���8����mS!������L��x]�boHi&�mp ^�v�M��/�t�nc��!��4�1bS�u���P�ٲ��"�1z	���Mz�z|De�نv���sb�<y���Zw2���j��-�+hՕ�la%�5����/N:�sL�I�\.�2����ދ�^�������;8��,�y��h�e3����S �WC#�V�`n[nV�_���Q#��> ��1jݥ1�^����q���pD2���	o&�1U����-N����������u0�nɂ���U�0{T�Ki����u6Z;���j�n������<��/$���j�q���W+���}��'��K����x8��ӈ��\ʊ}y5�]<�cȤ1��.D=
�0u!|J3�E�x0�)o8��dؤ6`�h3Y�4\��'Xg�9����Ei��ݺ�:�4����!Snc�n�ܯ��ȋ'�4C±��8���o m7�%�_��$��&�݈�*�ѵg�)����k~��J��^9�<�~͈$�m�+����/�Fؾ�}tYWr��؈���d�Ս�fb�\Cg��Aתp��*W�~'*��d��
�D!^��=���;!Ɋp�ޮ��������7�gv�K;br�>��j���P"�,�.-��*�#fq �N�ĪK�O%+9­��h|��6��r�iߘ2�lZ����$���va�|���8�~a��c�)54[d�s����GJ�̫\�!H(8R٦N��8	�"�v�L�=;�h�D��j~:�دT1�H�#F��~�:d�S�bS��_�����}�^�=q�p�~��y���맼߉�B�����W�Vx��������{XoD�']Ha�����Lk�ԭ!���gj�4����4��P�P������2���f���t�|e�] ������e�P���X���g��Uh#k�@��)���v<@Α#'E)QW�n����<+s�F[h�S!+���lί�û�=��^#_���z�!yS�,A�����?{��Ȉr��lv�;�$�D� L`��ߝ)�As�Ț�Xr��@��T+FW����Y>?�쁆���A�!5b �����'=D���왣s+U��QgE��������$�4&�e-�r������c��Ի\��^��\O��c�o� [��*�yD͝�oe�6�p�N���n5���ʟ���s��q���*#����n�&�ژ�'�p)�=��,ss<�p�<<K�����=��4tak����Cr���������eӲ5G��E$��P��)r��Sņ����ZV�>�[?�ݜ�1�W�2P� ���G����O��w�27�K(�Ǳ��2*jכo<�1W,��9��g�ѩ�c�/��?�2ㇳ���+D��o:�KG�3q#�����ژ���EEl�E"	^KQ��^h�AB!��1���̗�������<�rA�U�G�q���W�6s������:�KL����<���u�io\z3�o�l��i��InM1o��\��alX��MNF��8Qщ��e:����3oDp��#���M(2���e.�L^=���0�b^�Z�H�w�� ����WyɎ�ty���q��uy���l���O>"��{��F˙��S�]��D���\�����R�����m�L(��ct�>< �6CϹ^!%n؅i�X���X�J���wC�,���VV6��x&=z�(�Y�(b�!W�B��"�͙��qmF��0)p�����������yS��.S|�j�5�2M��^Y���ew:b��Mо܌�8��" �\��Н�؃���O5Z��7�oa�ۨ ��S�X�_00�^���3���O��<�74jZ!?�r>^�i�[|U��	'����=}��K/r���-q� qp!��xJ�q�QMi����V?�r��~E�s��m��%�<F}�q�4�!��2�u��4��-�\Y�ndw� �٩)�hn|����7�F�������g4�o�w|6��(�����B���`g�"�@s�J�:�_��A�z��F�	�Q�M4��9�a�O�2�q<@h����X'Ż�|w3����1�Q�!��{7GiP,Il�/n�ٸ��zJ:����LA�!4�C�E��p�H-:1u��h�֝�oL��hMgϺ��;�	-Wu��%��/����V���e����	�կ��<A����t9��#u�kl�'0e.oY8J[�m|oooc�W;��l֭��w�]oX]ﾣ��ff*�l?&<2��^��f)Q *�'�)'�|ct��`3���U-�����ɓ.�9�����5�|VQ�sУ^��w�R����v���9�%q��!É��=�#QQ��uԅ�����}h�^w6\����D�j�U���q}�������D�o=!��cD僻(��@���B���
���xz�0?�~P$�$y:%�y]t�5�9�J��g�����^`顮�o�PZYZ��#Y��Xp�M8�#ލHG���s�c��_4��Cs�q� /��b��ř��Lb"���lAw���SY�5E°���[���P�Ũ�C%i����-/G.̑��MAj>�@����4�{�Ѐ��!�
���]�:W����Y-j͉�))"^���/�yfC�.�PF�O� ��3?�1>���x^���q/5]x��l[�!��[~ѱٟ[LX�D˗w5����-e�cd��1�(
e��\�4ݙ6�#R����u5L�<���L���O]u��9�:��.³^��#;0�(F__?���
�l'����Ob�1�ЕOM6�ǥ��y� ����U����ҁ+�Y��G7��O�)m����sQRHeE��_�^D��z�n���ck�&Z�P��db��Dp�KRf�.�;@��K#��S}���{�w���tT�����!�.=jTƽo�c��+��5�x�7(��/߫���b�\L�>���"�a���A'\]9�k<�RC�|�a�o�X3�ybj�ѷQ9R���;�z&�'�߳����9=��4��Tk7L��P��G�v��o�C��E7N���a���C������ל�қ�g	�!���jZ��gIY\b�/o��<���WO��p��N=F.f�H:,�-y�2+�&}��J0>�'E@v�>!~����I~f�x|�k�E�@�R9�Ӣ%�|g� OX,b#�	P�9������m���̺p�t�R��"-V1�Xy@NE�kNv%��?����=�ͽ"����xv;	St���Z{�Џ��"u�GZ����LeS�YG�֠@wꇪ�d6x��=7�hb�Fgc"�����D$;���l=�G�_��_��;�'�o����v*��TQ��B:T�g����|�����?c�yT�żo���d�.wb3�Y����_r�%�3�X�d���ψC�xQ��?�AE$�3.A����Q˖�J"2~Fڮ�V�
��CJZ�����y��,>�\�>��Ul���*Zl�2I��[N��m�͆�Z,?�����Rhb�����|��g�#{}��eR��{�HA�����d����*�-с>�|#�#艿�E
'
��ɔ�^Y�R��o�?�Z������ ⡄����	}����M����5?���[��*��ąK
@��N�Ekj놎]K9����-��}_>�m����7��ן���mԜd���>f����f�K��q������0��I�oVg��1(B�f���B�|I+���^�_?���6����G�6��}���o��")C�e_Ry ^�~A���޷��N�BK`XN��T$1-į?M�N5,Vd0rC�M��X�To�����p[2@��8v"�ڣٛ�m�C%�s�M��T# $ە�z��j���@��EmM]6��\�h��� �oG!	L��4_m����8��ɳ;�}�я�ő�O's"��}� ���e�'��&@�t�	k%�FĀ	yj�R�8sǢ�׵�gF��8n�;X�̢�o��8:k��bY���-'�4ǝ���[�_�x���tar���*T!EE��k�V9��
��̬�1��qC�K�؈��wae�%9����H	�_��ﰤҥa�a��;���KX?.r�Jj�T�:6n�"$t���5�����w�GP��dha �PfSq�t
��U$�����r�"�4��kq��HG����Y�;�Z`�4�N����
T/�E1Qk�2�#��]8M��C�:1H��]ԟ�*����E�H,��On�f��M|6����]4g��^gɚoQ+���#�<�Q��=�E�׾g�n>���_[�)�
%Ao��Ur�&^�_��_/"4�Sp`�a��huQ�`���`�S)܌��l������w}��
�V��p�|�Q���$"�<�O��]���s�`�ۂ�8��jP�'����k� ���.|)]]_Wc��	�/��.!Vǉ�q�{Xޣe�7�W�Ǯ�K���ž����?>Y|��ph�Y�p`G��B��C�^w���׏x关x��z'�P{yQQ�^F/SR���n!�e\�vʡ��⽂w7-��`&\�G��)��Z[?�Ƭ��<=Y��_��6���>�kJ�X�Ǽ]��t��7;�u��EZ���鞇�y�˞����|�-;�'�f���4�	ޜg��K��v	i�k���^�W4uЊ�)	f�y���="BTwz��?
��N+�q\ڦ���m�!I��A���:��ڝ�T�.^�a�t��XBn��\u���u߫���rv�ߦP�5�_�6Q0X\��7*�_~z��[sy�.�ZiC����-�>� _������%���ӎ����� p�"����-+��p=[������e�}[0//�|U}7`eE��$@��=�a��wR�[������As�{��{7ɔݕ4��yT��<�#�j����������5�u�t�O��J^���C�
f��$F��0�V�M�L�l�O���lӶTS�
��������ǛS��{��qꚻ�6�0�3ڢ��N����F�@:���ZH��ԷG8~�n��A�!3V�M�J�%06rm����ƚ��D��B�v��I�=dPp1s%$�d���ޮG�%wֱ��x>�6�?A��A���[�z]O�T�ǼN�1U]ތK��cR;ߒ�؅��D���\;��_,���r�,���x�٭�hj�)��K���^������n��ү��G��`g��i��z�&6��b�0�9���_(D˴�i띡�{l��5�6�r��kl)+�u9Xؾ��Zj���v֟�8,�R?p˒5l�2v�F����Q�߻�N�˰E��O��DR���ĠU�@�^�G*���d��҉�>6�(g%�!ApP4����xzVQ(�ᗄ�4(8�F<8�3�S��(|Qȼ��"��%�z����V[���B#Yډ }Z����Y�u�^D�ڈHU���P�RA��ǯvK��>�.��@�?�}/�5\m����A�Sgkv1�m���>P�R7�K�� ݄���;:^�Ŗa'vQ%�6^��=��R0�|�V�P&_U��������%�D"Gb����b�%��Y��}�.o���k�U�����Od�ȦAv�)��×�4���2�v|�̵�t�uI��gq�+D�:`�� Q�z)-��j���-�GiP��WNY�
��1�.Y�:n&=̎�]?ߩ��������`�j���V�<_tŞ�65�d�3mx�W8�G%d�
�՗������o�2�b��i���K��Z���m��^�������E�{�6b���E�Ƕ��{�����5�X�u�����i��T�jkkY<�L���d�����a�A v(jѫ>4�����a���;`ei�;_M��V}i��Î/�Q�.���2Q^l�H�Ã�����u���AO<����ݍ`�1�~6H��{���l����3�K�9|��̤M-��q�1�CB.c��������N�S��
A�.}�|�s�(��k&L��J� m	�Lg��]��ep��>��OQ
�=0��٨�d� �No��A
u$%��߸0ՠq�PB��x;*vv�[�F��^�?���4��?�@)�F)�b����G�����'���p (����,`�c�����1�Ր����כ�*���A���nn{ㄺ�A��[=�>K�7���D}�tx8B�csI�;���%s�8d�J� 1	��F��~�x�,�����Е��C��������kA��0'V��ts�.Q��
9�z�eźJkfK���.�hyby�}�m>;��y>�g1T���+ag[�K�'�����Z��g/�����qwoW.��0�-���(8'g��n7Q�v r���=���FK�q�i]BbM�r ��p�\�V���).�k��-�Z҄ZKҦ�/l-j��Ŋ���~��Β��o�`!$���8�j�W#����\�1��A[Ԭ���""* �l�ǩ���in֜�Z����|�F�p�ƋI�u4l{1K��p�(P)���kS��{���f����Rw�dJ`�Ύ껵?�Dq\�
�T;#V�s� �8m~�"�p��@��y�&�+d*�}EI��i�J�v�����sRZ�3ϳ�*����+A�2�tX�<��% 5I�c��]��J\F����q���jd�/)W������I�։J(Zpշ��}o��V��d+F6��ep��K� Q�qς}'��ϾN��	5��,[7����#�q)s5K;;��&\�5=�n�7^_w��
�s�W��b�Ji�%�u�����vLQk{���+_�k?�q�= �&#�4&��+����C����.ˏ�@Y��U��#��z���(��|�6#Bݗ�����Z��rS�JHȬr�~��������6�T�z�&�zi��;ޖQ�d�g�O�[Pn�|x�����'�0����xx�3�auK\��rQUhd���ճÞ0�`]�hС+�d-��L��ǆ���`�F�v�V�I6��N{�+|�֮���U���U����z�2#�)��魊$��d]UygfQ��FYLwZq"�����ׁl�D�K�H��d�-+��ѝ��|�:���5VŇ��PS���y����`_�r�y�k��BT�F�gk�}���ԆF4�(NM8Gi��}X����Ub�9��H�?9B�n�������rb�/p�d�� t�ϲ���,��GJ�#Ӌ4�m+&nL.ˤ�*R�ë��_ya�_p7r���n8)|E|�p�,��5���(��z�)���uXvL}{����/�����[����暛r�*�5_���_�"���n�KS�;��K�}o0����Q�����vO�1e����n蕋�+���8�hK)�	������uU�	uh�`jތ�m�R�r�a+1������Wb�>�ٚ$��Wj�3�PFGZQ��.���d�2yy��M�c����d�DZ��{ˠ8��[4��www�w� ��!�w�����@plpww���έs�Nչ?�jj����ٽ{�^=5��:�\�3w޷�ܓu��!���<�[�x ��]g�@��=W�A��3h���đE3bY��`���_���ßŅ�ʕ��=��puO_��H���K�G�=IB|g%�L�A{>[[ ��'{��^���v���)�~�b���:y�]�b�'�BGh�f����~�ȫ�Af� �=�����a�����>j��)�{���sk�1y1�dh��G�Y^%
q���2�<-J�[�,���7�Y���
�D���+C���)����� }�"2믄Ml����Iis=�Q��݃�6P�]��2��!��S�@���u���qa\w�0K�B� j��P�C���[=B���6��R����fˁ��ܤ�_Uc��C�!�tJ�}T�a���T3B�����@�~�*l���@��ȃ��?� �rl�Efa�;��@h�06���oD���I�~���h�y����xZb�o��br=���wP�8aNA��
���ƧkY���
B��t�JV�����Va�+:ɘ<��
��5�x���~�C�h�z�X	A��n�cT:�C�8�<�b��l�mj�~[7Y`?܆JɤG�:�"�4Z镻����N_`e�K)�k�j:�p��,�.���~���(�71�3C�K���oa��}���K��Z�J�W�)ṝ��1׾��)2�ChSLE���'�������F��K3j�7`�C��/f�"
�~�������������c�nL�Hʴ��~�><���J-w�I*F^䰹��k�2�Ij(Y�K8���X��s�U����$�W��6�!-������=-?ɘA�Q��8)�����_�����$%��qv?��p�S�~�F���xl��0�~T�jY4��D���rx�X���E�	����	�-�/�	�����9(�R!@��V-�y��NgkMÜK��Y��Q
���k���	(��\:KVj?���}�,V���,UZ[�(����!ZY2�s��O���i�~�&х|1�y+���
t���suI�s��ެ>�F��.@�+���{�S2!�7�� d�;/ւ�*� vy��g1B�}5 Չ2�e`ט6���K-����6g��
Yt��9��Vh��b��Dyݿ<���2�/���Jz;Ylpl�C�;�����}B0m��)�[��Q[�ܶ1�k&����Φ�f`�pBȴ�I�Y��c�(;��J�6��g&��Xo�Z!��$A�c�d��x�h�my��6��W�[���,�>e��t?���_~���J��Cp�%���[�����2R6:��y�S��\u�o����������~4���*v���UM���G�V�v8�����k�u�oc'w��_u�_��xH����Uڼ���4�#�v{3���U�r��V��T�r�ž���B�	�T�nA�]�|w���d���M��+z�XP6µ�JP�7�Y����]p��Bx���-'w0�6�=��w/pcP��Bf;u���gZL�u�-�[[[,�0N`�_�Łd[ΰ��$�0W3}q2:��!zXS�}m��<�Ň�d
��!��qi�q�NPdd;��p�=$#�96\��y�����C4L#"bbѣ�0��:\J�$�I+Z<��� aoM����s�Nm2}����׸�܅�C�� :���E���0a�'��,=�H�-���� J�A��?}�D_�-�RR$�O�q��2���t�:�;�Nb|i#�hVw�lݧ�^3�xYjH��x���ᯮ����Ö'������Ó+����-~I2���m��'�a�*�ha�
=<��O2*)���1H���6�ځʖ[��)D��Vva+��π8�3ǿIv��D����w�c�f,�~⢻�N���v�P�ys�b�=��(��nd�	��/����y�'�b<͋:0�`�P�W2&;�s_j�C��v3H�z;��j3���B�����&$�r����p�t#�V�\���,���U�ɤ�Z��@T1ߘԣ��_��r�#U �� |4�y@��ޢ�v���Z��w���0�{�d��v��x1Fx|�ӷ.�d"}���'�4v#T/"��L�9j<�ҁ@L��3�P��ѹ�ڊ΂<V�|;2<�0��]Ќ3�U�6U_��⫱����1|8@YS&ZBS���K��	���bhce 6��W[�������%�?=�e;W�\9J��x����h�G𑸞,�B�1ݬ�q�����96�����֙-~��IG�r8�����|����s�؛y�ޘ���k�JT�q���3	�t�2����g1�OD尠왦Ƨ���fƂ�=�����*vB��k�a�n�S�=g��N8ב|='0���vW]x�xY��ãP'�4U�g��8i�³���qA��tH��{�8�D��u�Ʉ�^2�q�����D����1�4�r�Ւ���J���mեΔe8N�S`�=����M�"�<��E��S���B������Nw����G)�AB�*߇�'/4�ᠼHd�N7}m��d�R��t�W�St�8tn�A�A�n��<�d�5D�8�޿&���6���ORe���͓�c�jzJ���F.-�;��|��k�_�Wi�i8E�������S�3��sR�I��:�Z�P�oQn���Zw��#d�;����e����7},�2��\����e��G���Ŝ���;d`ϝ���Tӿ!/Z�z������汛�I�VE�s��'VYc?ԧ��B��M�ڸ�|X��8{�)�����<P�Ѧ r<���p|\�?v��u��/>�rL�\�g&�?r�bį�/�ۄoU�������y�ⷞe��ӗ��^����"��7�-p������-vP���=�K�\e�g�|;��K�D*�I�C]�K)cߦ8jR!��v����fĸʔ������*kv	��K�N�p��*� %�ל1/�rC�4��y�t�oc;�5 �u[R��M�ZQ��R-~�}�_3���<�^�>Y_1Ru�[�����f��Үh���}��h@��'�o�>���:���ŁC�8�)�>1��38 [���wph-S���;~@�C2ʥ����Ć�V�$�% 
J���"^��o�ϣX6<��!��R[�L�_�`��{Ha��.�g#e��㙬�y���_������ ����Ň@g+ct����x��Op��+D��+�imm-?>�R�6N�pw�G6y�e�e�:�s2��D�r� +	No�2u
�>TPru}on�`J�ĸ�-J�6�H�)Rf�F�'�����ޱU���q��9T�s�h*�H�!�����P8F���o����:cԇV%�8ح��X�]�c�v�:���h2�K9rݜ�+V�U�2j2�k�� �4 �������y9���ȴc����p�,vu\������!�}��Z��G�-���`�*�{<�ݐ�|��!U�����R�Ks�Г�n��䈹(��nw�'�����>�E73J4��������b/O	�-�Ǽ�i���A����]x��D�E	-�[��j�G4�z��U��P=1�����(ci�y"��V;EB�v7!T��&Z Ճt��aa1,q�}O^���~�����͚:��J54�.S��s&g-�.ܑ^�f��sk�d�!Ϙā�~�Cu��qr+�3�Ӵ�I@w��1n�1��aj���ۡ���.��X����]�M�d��������Y[�P�87[���X�z��t�p����{M��YH)�� K���R�-Y�q��ծ�'eZT���)��@��� 3(���ib�'{z��}(���*c ��`�;d����;s�~MW��G�F�������
���`q�+C:g��[���Q��ﷅ7ї�~]F4��[���#�����T1�zi�:��O���=.{Y䈸�C.�8W�TBp�qC���MMܒ�����X�`Q��*tT������d����� U��N��#��;5�)�Ӷ���?5�[5>�+RS{p���LK��_,�z�d0��9����T��u�˝��a��?���ml�)��*�6���uyJ3��!�Qwq��afW�����Y? 4Qw4�2�&^�G�#k�c�ʟYd�����9C�h:Hu�I�uc���bq�u��襬DO4H��rE�'�d�l����#�,Օ�V�l�9CjU~��ulů3�d5ND��0(�2�-����V�l�w<𸸳�B17]Hr�:4[4�W�ǈ"��rx�{ /ö��:ڬ$�a���?6)�0;��gY��x�����A�o�$�gd���{���Qnq{C���Z�on�Ƴ-^�;D�FE�^GG+���E}L�C&�y��=�`�E��$���#��G�xr~����QG�ۋ���AC�����dy���}�X���+���<���%�����
Sǯz��f��'�7@!d��7D\��ܚ����Ħ["���|��5[JA^R��-��2���]:/�Ҏ~!� �2��p���I����D=uc.?��pR�W�y�1���|�O�*M��|�u�v	f`%dG���\t���	B��,������|di�5jzM�~|��cí�I���n����
H�s[������g�xwk�W�ki��~���+83&�����e��
������[(?�_-Q�(�p|˓����$^�<��Q��~}{���͗�xd�Ȕ�΁=�z��'�����\{r�i0�Ra� 0�����q�p؅!��~�L��n�Ϳ�1aWw�852yzz����A�S.L,���O��,�hy�`�t^����!���m��®Y�W���Wfx<1Q�#�xOh��I��+��p��鶌�Z���n��/j��('k�����У_=kSK���[��nO6�1�TD3X����B\��c����.P%]5�.+ёt+ѴTW+%5(���K������x�i�d�ZWt4vKP@��q���׆�e�wg��Ch���)�|
�������5g�5s�wS�c~i��Պ%2`gd���LD��`����Z��LM�����}v�.C�\����]���iIr7��s�'���j������^��b�j�ٯ�w��ٙi��sU�H��d�p><8�TǴ����|S�EE�xx{��h��J��w���y��g�M��}�'��p�����<�#G�<G����v�o�>Y.z*S�bJ�S���-�7�W�UcDP�(.8��L������"����R����fMR#]��JQ�p�!�]�։忪���.��x@��}�-��1�o��Ʈ���%ZK��Nj�+ᩛ	���8��@�*f�����as�p�%����Z���U��o*#l��������FH�q2�֩i����?6��Iqfj;�M��^��к����DJ��F�͛rs���*S�ۦ����h�4���_H��L/�����Ӣ�_��	;-�E|� cw�̤��������%C���Ɵ�w��M��R��J.����oK.�[�X��FS�P�z|%=I������Y���\�_;���L�%!�q_�����8Х�U��`�����l8f\N:r` L�V�o|���V�>B�S�X�UF٘���#A�l�嘞���:��ȋ>/\|��̙_a�JQ��SW
��D��)�Yr���m P��@���P��|��T�y��t)QCsB
��<?�CC p���A���-�W9��r2���+Y�=�SAXl:���R�����ab|�(�x�2�HVǓ��[�b�;F�r��NV��Ί��`�8�8��_���i�`|1\�I��F��K�׌�ٸe�EnK�����m�a@�v3������W�c<�Q�l��vH�R�@yx�AWwn�{EV�\�y�(:�?#HAK1��|3�+6*���Í��b� �Ǩ������&n��u����b�`��;�w97�|m���4O8�~���f��9m��\��?�*����[��m�\���[�T��m��x!���g�&13,��Cg�v�����⸌�KAZs�0���9 (Ef�[b��]��Ӎ�ș�5Z�]��|	ݰ|	�2j���ny��9�/p�ἦ��0Z�)Mt�d�+x����s�W[M� �B���%Zk�s
��CpZh��)o�,�KE��:�ki)�[��n"�0�U���UT��3��m�hşH����3$��q�]�:��.��4��ڷ&y����q{�-E�)�(��S
ډǢ:�-��需_�b����!T�2�,�D��&������G��\h��(lI����	~讥'��E��YVM�ݠ�	񬁭Fő���f�4��ԍN��/�>#xfE�FP�~���d��e��3�z����Q��wK�
�6����L�.��ቹ�ng~1�e�"�өARm�z�À&Lg���:�؊j����/�
��3�Y�I#k'NߩF���f�L�=��i��L.��z���?��tyq�d�6��ʌa�A���>���Q�/�j���T�Z<RB3î��N7-��������ݠ��H�ۤJ)Ա�'�95���u���shʶ����ՠs�*'`~P��<W�1m�QDf2�D�Q=��V�-�Z��g��G2�tR��./b=�~jr�ɫ�2��I��k'F�Sg�[�Id�to��|	��iB[�a&St���S$>7)
+�*o��Xs�`�|wqϚ�����^�q��å+�p\�5i�����$�ܢ���:\t=l�\�|73��b���6Ę6���ԙ|�s���m��j�#$�U.ر����>Mp���e�G}e�n�7����m����;�8nC��a>�3jZ����<����@�ݶ7���t�#$ R��fmq G�㎲�M�����uZ˖��������!m��@�^���։�O����4H/bվ����
���li'��;�;�є�����`�R�%��Q���e/���pppk ���aK~~�6��E���A�_����Nˆ�@�j��թ�9���E�3����ڥ�¢�����^d�I�9оY,���U�h�drݩ�/�e�9{�.����	�#[a��Ŭ�N���U��HDd��L�t�rY	m��d�S	��FGER��Y���l�jEz|n�'<�͗�5����WJ�ͺTO8������/���Jǅ��S�0��œ��r�|RӰ�:��c}�zfj��HA���曇�2�C��J'n-RbjYu4MR�UD˓_,��ki�Q�>9z�֌�-k�qA[anlP �Ti�	�@�*�T���n�2��t�0x���'#�s���`��DI��3�����}���o� t���v�	�P����g3#�XiB �6>�ݹ��/���sV�9�XAI��h�CX:ܰ�����:[�8�Rw��,�������Oh~��y{jÇ��t�ĸ�vd�a�w1D��t~�p:B���2\T"�K3��E}7�6���t0��mq���}S
�/i w�uy+#�&����������dF[)��./�������h���9���o���s�&1�	�JT�Ќ�%��K`�� ގ���&��?�l�H$J�tC���u�vy�#�*?~�u�E��5�'���;�b:^_�w�����a���7b4}���_9�����>H�{z�BDl2Gp�@��M���3xf;;�܇�����&�-�2����u �6��DL�
`�3H��^�,�/�W�LЈBkn��L����鯲x��l�\:�~m}�	��e�H��D'C�`�Ί�xM�3�-a{%E=r�D�	]��:pK���	���j��Kj4A��G�/�S�?��L��X���rA�5�LҔ��I��5w���&�E�B)�� �+lO��m�"�]ۇ�9Z��Ձ�ܒ��>�9�2����7�aJ�-ƽW��j�˞���qp3���>y��.[���c�\i}f�wd�'���Y��^䔙��qkb�L�@5�#>X��'����['N�,T��8���oI�'�H��߸j��	�֛�)/���ys`ܗ?R~k�X�
�z6��X�~Z)t�jza@��8��D��Ù�e
Ң�9qR�Dii��\�wo�n���b@؟ 6�ʙ�)���@�!����~���f=�"������ #"t�E����E����|�(���
�L��3Ol2�@����\�ɟ��"^��
^�@9�_�����o,�d�o�K�"�/���d�ԑ���KN]�d�؄�H��X�'-�z|	$���S1��~��&%%�P� :���Z^�+fp���7?	� 	����\����uL+.!Q�L��,��h��Eq�hoeE�a+�?�m��'sny7?CA�pE�םSS�):�"	R�/)����܌�[B�ڎ���bg%^�(�X#e�;E<�2ީR�]�~��Z�}���T
�(�O�V�Y)y�P�
_�m���f[i6L�;%�g����Z@ҙTH|!���%�
7�!� �o��
|H V���ԏml�a��%��;M�����$�cDt�=�3��<o^Ð������sVa�!��+@�޽Z:�9=J-%����;#��>8B�ר�|�gٖ���1�&"��`{'���z��MJU(,�п����4Z2��W�����7w'��~�7���{��� �)�nW����#�}{y X�tWZG��1�F�(HK�����w��g��}毱�ܸ̰�)��d�u)b�Z�Ԯ:݉�\/\}J�9e�ꈹ<eQ������5(�_��a�ǆ���4������d�FV���PLVG����TI��� T�����כ)��`��?X�]|4�f띞�5�� ���w��u���S������:��D�>��,���N����<�����GFy9���	 �s��r�c5r�ƿa�8�µ��=Y<4��HL�"܀y���r,\_d$U�_��Q$�A�?����xq�43G|Zf��Q��{zQ���R���W���Y��t����b��q���@m��ݩ����Q	����@�3�d肂���*���	DN��v��p�6ԛ�H(� �V�O�6(����>��A�R���A�c��-�L����u�j�]��E��_�8�S.��f��������5k����*)X�D��Z;����x�(F�Ҩ�J���mkm-���{�p���Osb%�e��s�hd3!���$�u�
������p�kms��V<�ySNdb!��	�x,��cT�3�����aߞŐ�Z�eTPL��8P}����E�2�N��N�Y���9#&�ř�1�������s)���T�@c]Dk�Vh��R|( @�5>�b�T2�n�l���U &�f�iV&Z��*�>d�v���ad��G�W:4Y��f���j6�|�Be�<����ϊx8~W����?wD!i�R؀'H��=m�n)ɊrYi��%�6*��v<��W0k���r^�<����4�v�	�?yq�+�r*V��K0����0�M�˺���n����j�g?�=C��F�������5Y���V�n#���?ǋ�{�
e�۩�>r8/c˭J}w��n�"U��|کg� �&��*�dK(<5�����o��סT�ѹ���h�/^;�u]����Q�X*���2�V�v�l�A��������D������.��X�ڱ��4���x=���:F�Vf�-9�],�y���$�ʬڦ~XoAVk92��(�%B6�h���o�]'�nD�!:&=v\��0�j;�`�]���*e�����,<������Ҭ���zAݔ�qR���T>��:�nfa)�<��\�i�:l��� �9B���|O��ö�T�$�V��� ���T9��G|��f�nH���Q�Sl'�8W��#�r�pL}���%q�(s2;������o�
�:\��x\"��]�9;O�NKqN�F�VP4��()VX�V6�T-�X����ْ�S�Q=���G�^������u@Ӧ���f9yQ�����AZ�ޓA��2����Fe�4P�o���Va����		��]�FD�ʲ5�ro�W}X!�;�i$|�ؘ&ֶ�ܥy�4��'��S�v�+3#�郎��W�����~2���8��FW�acl�V2z��h�w�E�`�+|'��M�����/�a�܈��^7������I�'���a;1��wn	d^7��~W��ie�ѣu�V�s,[x�\�x#�?��.�m��*��WE()��>Y<
.T_�gb�F��q�\�0��J�ό۲���|�rS�(>5b�R^1�SW���5F�ps ��i�3��30T/�pa��dPlμ7�?���M���?�-����:��=<_�����$]Uɋ��:�v�}	�3 фW'�l��.�����sJ��YO��Wm��'^;e�-�9��r\�ܶ�}�W����[W������#��HL���5`��DŲЇ�\�O�2�PO��Z�E���9�"T���\`���}�����tE$tŏ@�!?Y
u��4Bb�
[���<G�4�]=|�>MSF^<LW�z���?�=����
��&
�!��W�O�*N��-{|P`&i���"���Lפj��9x)�b�n��U&�Ĺ�	��#���|Ć0���k�\D�4�*/Qlb�
��-]��S����;	YD8|�F��a�����tS7Ҍ � a����4�u{��v5mE�#�}x Qb�6�N�og�
'f��^�P�wml�6��.`<|ܤR5ɷ[��ʹ��R#�.���@6Rz<���Ǣ�c�����cNk�7��U������y�֎�S��h��p��--��H��A�=G-m�uk�K�X9n]�5�m��ʪ>�~��D>^�3�J޷ �˫��~e��~�}�b.���Ζ�1_I��)��B���c�.��K�	{�L�싘�U�������"<�#|n9VbL����M�ejo���x,x�s��n,�FH`�L��u��B���A���.����
%:��%'H��@���M���d�ٗ=��tj�*{�y`1�	>�t:<P<�l�JЎ�"}���{�8^�xt�a����M��7�
3C:�U���*�D=�Ƭ��*���Գ��(��B��q�����%�VRr���*k�R3 �oth���H������֭�����C�q�9�l���)�;���C�9B��Ȑh5�SG�{8���tњ� �CK+ewS����;b�E�\���A�Gb��Gb��zǭc����\��t[�/Mx�H_WǠ����ޮ7x}��a'�w���zWU'AtS Nhf����l[��ד�l-�U��#����������Jm��0[x>�!UJ�Tx�=�t!�]��HֆP	r���z/��S�,�b]�:D+�Y{��4r9
��֊��	�[3����k��|t��~x��ڟ�<�-_�ۍK��5u�V�8�^;��H�Ŗ��u��
�^�t���>�	3oىd��^(be��54�Ps���tE�@�y��m���T��9)��k�+E��7�\��
�B�:�L�����t�	���+��{M��q�Fw�����B�"�K*	���~ӻg�n{|�Q���Eq�^{ϟ������u]QQ&��������K\���Q=dsws;���L��:U��(0ob*�U�����,\^��z�Y���lt�0qL�?4���+/�-�7����^�4~-�XK~#����F�--����^��H��qga'c{)��D!�$�?�kc]J�])2���S�,Ҝ�aaP�_�n�Y�5�Yߗ�r�ϝ/�|�'h�������˹X ����9���O,F�F	i׉�_ϧw��	����
U�$��F�� �\[l���~vtT�^�3��I�r%mk��R
ʼ�:^i�.%�!�f��!�b;w�Njq@˧˶UT�+�D@=��Ͻ���=��_�!6if��}��hʚs�źKJ�#�j6��B��|&/[|<A㝳�`�oG3����#<N��pm*@�쁄'���
x���:$��Z���8����!�4���{�)c����^!"�;8�Ɲ
������}(��;�_��Ws_,�1����6!O�Muzq��u�J�ip'1�pG(��K@kS�! �؊�=�X����i��EJL���{�De��;-��҅��uY��Y����)a%q=փ�1�J�.���j��w�K��N�]��|�|���y��m	�M�n>��N}����B��U���E����|L
.O�Y%W��,����k����[�(��������QdKq��U^\�M}���)�:�z��	^]ʩ!���Mb-3pE�˴�^A��b��>���v7�w/@�qu�с#��o�6�;{��N�K0�Vb��}c�Q��u��W���f���VdLu�b?M���v������1���^K�-aǍ]��f���Y�y�1݉e���i�L�U���>qd	K���eu�{0?���a�s��M�,C<@y���V�o���Y���f��"N*P2d��$&P�֊�h��q�A�j��KlԿF���"�=��g(�ˏ=;��ߍ�&�<!$bKi"����'.�������h�튍X�<�ԜHi��4� =	L���)����SH°2}���=��ʴ2�6����G�5ѰZ�����M�S�uCxt92O[��\�)7yB�bz����k
��h&�o�lL���4C	0g�d�X���/;m��Z[%���Y����*�T�ƅ{�'�R��.���&��u��R���s��a��h��s0��s?fx� �>�{Ԏ8db����C�Z�(��z"�=[��8��B���*��֪�WOʬN��s��B�3�	���J�8�8����4ژ�˘�R	ܗE�U��(SHԌ���gd�crt��`$�C{�m��T=�tѰ�Q���"�Z,d6�E�Cý�f(e�U�2T$M@�v�w�����M�n�1X�����U����NǠ�vf�<�G�Z�n$>b����ԡ��l�DSa�pCC�P�3cw:���Rc����e�Ϙ<����f-�)�܁?�SmM�ڰ����_�CDYjLS�II��~�Ha��aӉ�@�Y��\�J�tS�i�9����0L���8��y��@-���w�E�1�h��TOX�IS��z3�@�qO����vˠF\;���x�m2F�1����U�qC���k��d�#q��}�`$�=H���<׳�^�䠪�uY�BQA��P��� :�`�S�u*4�.�������x댒�����zߝ_�\VT��}�p������y"���	��������>�`����D5����o���������:Þ��4�ѷ�H	:��a��z�GQRK}k`ݝ��-']���s�)��^�x1nH��w��ùۂa67���+��ŷ6�#jj;��p��o��7��	Φ����t�%̓���nj�ӳP�Z-��@��]y�9N�?}��J�M5�(��	aTH�A�"6#��!�xẌ́�F��$�PYs@�v���w���*R�e����.��W�����Os~@�)E����,�~_�1�L<>��8�,�������J��X���ꪅ���&�Շ���>e���Ea�:bj�È���E������?�N ;���<�t4EP��s����FN=�&x �U(;��.�^Z�D�ѯ���[Z�	B!�*w�Z���7��mMg�%��6%@�yl{�-������S~�^���"�2����3�ٸO�O���N{��27�*���,~ �@F��K����pٔ~��/���B�EK���K�ꙛ�Jt�Ej;�]{
D��bG=��?�"
g��G��Ҭ��}O�P����J�i�����#�����Xr�)vB��s��X6�oI����7j�n�d�O5���f��N��B'�}>^	~�h1j�)7jc���u�މ8ӏ2Y��R�  
b�a�:�.�%V��!�y��xB�E��a��� a��mBllh�X`G�]�㳕I����*[�;,�0z�T�`�dV�:�œ�9�S�|�����}0d>������|��G/jƼ��7ߕ���.�t�nm���O�]��C�Oh�ȡE%/ ������������ͧ�޹ϫ�(��dt��)%9w%�#qu�ؾ���F�??t�����}���/��Lt�
�u�"3m�Pϑ�%��T����q?��[h9�hGS!����2�xl�:r�^c�TUf���}����6��3�	��̫l�=�-b��q�]-n�&X�t� �)�������j�Յ�0�y�sZ�Y0ՏW�糅@S{�ĒW�ko����	�nx\��&�Td^��W���Ρ�g�.6�ˏ�D�H�s����`{��P\ ?k_t�g��J/��J~��˝�m������0�r���X�@�Y�1�j�֜ϺG!��ְo�u�(��3R=C>{>�`�o�|���Z���Uz2%�����^�X�� ���'���+Z=Z`�����tq�0���B���/8BX��qq|��O�~���Bm/�0���Fr�n�3�N�t��"��}�/FRG�AKD����s�3�|@�fzHh�7�W[�]r��w�������}u��}?��֬hЙ������&ȧ3����j5~�Mᵋ0�R� ]��˝��c����(kjR�:C랆�ӡ�9�@k9JRy�o�?�M�6/,u8Z�R�v�����ܞZ>wE@:��H'��S���b*a�'s��:�;Ĵy>pi�$���d�e��Z*�S�:e.�ȷ� �/�0f>(SN�EV8��a��;L���$7��+����P�3�Ƿ;|A�^\���(�<�e�=	�1U�;�G�!�V��]/a�%��N=��/КR�R��}ρ�@3��,�O?����oUm�'�:vkv�[���J��-��^'���%�x_���w�Ƨ)D��#l��r���N�yr��8>\oKc��$~H^սdđ6�����b���3H��ƽ>�:TIC�&:��{5��O��Q8��$���`��������%%$oA~�d<�B,�t�ܶ���=�?�<iK)xC��A��9�S���z�J��j�2��O���G1p�}]�-öʜ�e��j�ֺf[�Z^/��_���
d�(�4�r�PJ7tu9#K������*jmկ�'e�i~�*W�ɠ؉-;�r,:,�,l��$N�Ծ~�^��e?��F�'�`��i*�6����r�'�,���Lif������s���2u(u����1�i Mm�S�θQ墣 m���~f�]�g�뿃 �(ֆ�7�ڕ\~!�g)F��I�T?Z����S�xJ&2jB�h8�Z㬽�d�i���O���D��yS�$�:�]�X��'w���!�e���#��˴�*�'`��7A��53����k[���F��ڰ
��������h���ˢۜ'opv l�B=�c���8z�E����K�Sf/�_b�&��J���߯I��
 ���>7{cs�gIK�h�^Ղ0XFA�Չ�A�q�3/p7y��<j�^p��U%���R�2��RH��K��1&����>��m�	��-*����D�w�y����OZF�I�'�/�|RI��n��33!��f`�c�s�`A{D6�U��p2��Ji��+:s_�oc+����6�� @���h�xIY|ˡ_�41�Ě���8t��׳k�o�,����,4���W�4Vp})���b����P���.Qnr��	CI�r�v{�� ��ބ��f�Q�uB�s�T�[��]�/s0.��D���)����p3��=F�$n���_��K��y7(�]��B��>5���u��gx�Zu_~���H���O�Ɓ�,w��cl;��f�����.��qg�j��(�c���6� ��[ ̧Cc��t���)�%Ά����t�[��[����5�Vah��ݣ�b��޿��_)�����w����xg��9�b�8��R'}z������� y��={�� �M�}�W`&V�B�d3 U�_���$j�����4�~�v���'<'�T-��A��xd҆=$rY���Ch;��4�m˖϶wi ���Ѫ���Bܵ�b�� ��>X��P�Hk�"�1���q�ʍL���X�ϭ�|d
�*@\��[�k��h����VR�4^
�����y_�"����X]J&����8�f�q+w�]��l��%E���e/�%7�����n���͎0��8;&��K����G��թ@���[u������ ���)'*���&��f�fVun=�Њ
�����܏����;�k�]�|��y����3�
�W�$��������+h�Lpw	n�.Np�݂������sqww����0���5��Z�0�������ڻjױ��{ֹ�t�������x���B��ƫ�����}�_�%n�Ų����ۀ����Ҍ���G`Buk�43ݹ&��+�ڷ��ڽB���Α��}�bY���8�$�9_n��$xܭW��i.�����m��,���qH���U����d!.#�ï��]�s�9���Z���5S�H'�!#U��l]wZ����]�$V:IQ�M���z�n)�dG��ȀS�6��Y`j>e8�&�;�Ѿ>^��|(�Z�ݎ,���R��N��i�{�;ᕈ�V�U�l� e�N�i&Ad��\�u����C�?�㰃��k�Vm�Ϋ�9�
����O�~�E����~PYE��F#� {�1����u�����������l�Y�.����i>�Z
��yg����(���4�f|\�3کk]�lJzVH	�z�s���<o��{c�c���;$�a�u�j\Ҩ*U�L���k�md`=��j{�¶���	c`	�A�������{ډz��s9o��Ͱ�yc04EU:��S�*��A�A�z�����~!غ�)����1�䮇fB�"�x�ѽ�}�'1>�-�����v��8=1���Gco�gF��AZ>�EH����='+���q��"���\{}&�c;�",�w�L9����QXe�6v���2E?��b-���_t�$��"s�?�vÞ̹:,ȅR6��C{t����9q����l_��f7ȉ�7U4���=��fۘ����\��»Q0�1�8��Ю���0�J ��������%^ýkʯ� �r�Iu��uW��Ic���wk�s�h[	�4	g�w�^�������8���.��8)��?g�(�<�_@�~�����M3�����)^�z8����AP��s����
��	����Z�pl,���|Bp�2��wWn��+z�݅ug-�A���5Ԭ��%�[�sB_�6��R�8T���jA��OuH�eƀl�8���FD6�	����z1������R/�^����;s�{y�K��4H�c�9����F�6͛q�!�IQ�^�(ڙ+��C��0�����M{�K\@��,uԶ#�. ,0�`���C�4g�y%K��H�=wC��0�Ú����*w׬!ܟ�����AnJg����I}S�����i�o|I_�{gu��QC�0\�����Np�ϛV`Χj��E�ҏ�a�|y3S��u��Y��"s�e'=�;n}&����9�2��[�8NW�ڤ���0SO��݆O��.=|�D���6 5���c%&Ժ'=}إ�U���ҕ�O���V�����C���t/K�:�W�S�N�hVF�!�K�QĥŮ������̾�_3r7��wٝ�q�����u�3S����i�u�)F�)����>�-D���B�,ME���S�sZg4G׃Sv���l��l�x��P������t f�;~ ��bH�6��J*V����0�e�4�f^`�ڠ���}+�y���f���n?�xp�u���1��χ��ǖ�@�kT�َx��ni��%���>1r����s�c��<b>��m�61�Kܠbq+�n�����O�VF���Җ_�Xh,U�2����r[G�Rk:||���.�-gՂ;S�`�ǆ��k��;.a���k�a�t\<�#����ם�*W̻��%V��" /Sk���i�snU�԰ż����2����ёҷ��*����,F-&l�� e xwy�01TD؇�_m�K������،~q-Ҭz�l�p���a����5�Y?T��(�s�Z� ����{��y�&��.�g$XI'1p;ּ�JE��IB��D���Z�|�u���(t�w/G��J*����vGD�^��T��0���p����ji�k�,�09?��5�g��;�)�.=���*��� ]`S�S��]%)~J;��}^�~�(�S	%���G�摤c��Jmw�t��t����G,{>����K�5��;��!R��_�ȶi;+4� �+�Z�NB qg��ּJ�ui+ |ek,GQ�ޝw�����h��n�0g�v�T.w���rs�>
�V'�۹�E�l�� '��Q�
V,N���U��`�EԽe<����L����Ի�!t�Ƽ/Ѳz�0)w���}�CAL�V9F_W1Z+
F)�*��0n���}��yht�&�y��ƪH�������N�#��*փ�C]l��pT���*�hǔ��/?J?��u�������6��E��8��~}���3r;�nu=8���iA���ob��ԑc����q,����C�L�Q��<�"�N���������H����gւ@,��L'Ʋ� �<���)V	M�R�%�/�)A�2�a��ȝ�Pݙ�����y�S�؉>>	]?X����\�l.��=�u�>�0Mw�p���-����dr
�BE_M����s�]�o�Y�[-;�ܥt����ܳ�Э�U���H9�qiY�ڄ]R^V�f۝�%�7!��	0a��%_m�5j<Q�4��+:R{��,]�S}.�U�n�O��Q@?\�@+��F&���6|.�Ƴ����?̝���Z�&�Tյ�#�pO�.�9��e��rQR{�A��'y}פKq16��
DB%D��t��d�XJ�I�ul���J����)�ص�� m������v«��D���<���R��r�/�鶀���*�3v�V����H0��6�՗���ޓ��Y�����oA���f�f���6^��G����kj�}�~�O���!�G�8$r���$�x�^v���^�T�7�XY�E��4Օ�����)�PtAگ�2.�n���y�W�K�%�uy���v{�(�̇R''#*1��[+<��Niu���%K&ZP9~�=�;��s��4B�!�.C��R���.'��-)HSBz�u�e�I���A����g((�K}�Lų�g����E��V��osՁ)͂��!�i��%G�W3\����n��Kع�u�6��k��蛡H.Q�Q�>��\�l���� 8�/�K�/�L�,�)f��,sB��YyZ����@(��R�x�R}}��LM������HH�
���UnΫN�ap�ӿPb�tK�O�&_?��S0�n*��8�?X�FR=��ٳ��ھ��!ޠ���}�&/Y��T�y���������=�?(3/�G�=/.4w�? ����/��6�~ù?|��V���p��[m[��Ȣ��j��EqX�c7��Y	6�W���J<J�SZ�Q�(��1��!��r�k�c�w���S�䞉 '��;�Z��3D[�Kъj�n�JS�����#�3k
Bs�|t�)�r��s]=��S��1��$��#�d7������i��3V��n��pj2BWmP�s� 5$T�nXV����;�r�������iE����o*g�	���1�2��&���x�?B#z蒭)�^`e/�5d1�*�FGsJr�w�]�m�'�����&��8A9ˀ��]ES����Y5�tU���=:	�c��(�ؿ�F�ڪ�"��i�����J��d�H斔v����Tg�Zc��[��� Ϥ�VIFrz������"�]���R�ѥ"D��>��H���E�9 ��d����k7ڕ���t�^����'����PB�@������ؔ�;`g�,�8�ƓC\���|t��UQf�E�ː�f��֘{Y*q�*t�<����M���ѭrJ��i�R6��Ps䃉��r�t����w,\����oӰU��a�����oA�)�{�%�?�>P;>{,�O��3,�6���,/br�f�GNd�Ќ�+�$����RGp�D*�;�Q��O�1�E�j���a�Ʀk��'6ս��w)�������=a����êW|�n�;B~�`�,B"|ҭ�K��m�)V��O�p��
��r4~}M͐�7�Y@���E��zjQ/^����;T����9�oo?N�U���&ew`�HG���1A.Q��I��cc�
J�t�ɪ lP-�YvE=�J��k賐�"ҵL�^�,WMUHQJ�����}��!��q
7t�����0����V�����o�?��:<�f�"�+���#}b���H1г�� ��W7�f}��$CcW���>N����< �p��}(��9���ɚ�S�K�/'�!���8�rVV�ྒྷ#�+#d��O��<�-����K&����j�wm�ۆ|��F�=�>�]�����C��O�'}}}5��4���b0D`��۵�:$(Z�6c� �j�p�L���������3�����������2��q��3j�X�Q�����&jkC�����Y�� ���C
i��U;��v��1���֤�H�<n٘�T�����a��1($$?7���J�6''g�+:��p9D��H����ϟ����w8L������YeA��:.�I"Z�&Ώ���`n՞�������a���-�Й0p�V{
�K|S�=�k�CC���5!�fN�bn�S�GC��pxoow����7������&H_�?��e������Ē����ԛ����o~<�.Vi���ة��C:��,�|NKK�ҥ�������}Ɵ�"\"� �֌����2�[�<�ި�րC����2V�����$��j9O#�Ń��C�]\������E�Ύm�q�O^X�ӊ�t45X�ZQ�qg��v;�~X�9H�g�ebd��z� j��)T�% �u9��E�^m�����=���������
W �q�{�E����� �ѱ0������-P��뮋(=h��y��tk�s�����3{TX��rI>0��z���(�8�eL)�	8Q�ׯ�{�_NJV��b�WW�Ηk!-,,R���t=�w��t�L�?���l4X$����^4�t���˶y�:��Sn�uѩ+ңT_e��6�����K��P|�J�QgK�����$qt�N��3��8�ڔj��Z���4[�ɼ�	쬭���FEC~����8 �����Qы.�twvv�q5��'��~Q��)���.�\��i7�	ä6��K�h�z�of:ǹN�����?[��&�An�6@ϲ��p��K{X|�{�$FHDV���6`�3Ĩ9h�H�l��`n�*,��̾�<��@+Ms�;�e0����\��Z����i�3g��?���� ���(���*wo,ZM8��c\��P����Po3n�r��A�3ێu�xa�7}���{�ީ�B���ۆ�S�Э�aX�W�پ�
�a���p{�s�>��^i�	�Bں��~O�?��&%w2�g��N۸q��̂��vx-�ج���L_��o3���~��Mu�����c�V��&@+��Zct�i�3<�{{rX�8�z����TSv���\�9���i ���{���^�ކ��Q�#��j�[�8���yj����~q��&�#�qV��W���F��L�s쵘cGj[����?��'�߼Ħe/ʌG-��d�O������|ן2����Ki-���桼�-��a�^���G���553�7��Q�yB��H�����L�l֚X⨶�X|^�P�1n�����H7�/K�eU�[5��(Uc���xs���wB}yM<�em���Et�}�AAy���-�`=�쎻)��Ά,�-NL�{�zӨ�/՝�wZ�����g�!��c"@���gv[�e�m�="F������B<T���eI�z���̐�n��Pe�31T{`~~F��p���y�t��
����`��
*Pawӂ[�{�J�ɻ9vj2�SΜ\-y48�[�zF�ӱ{��_����Xv�/�v�E�����,JmX�&w���e���xBv��受�+�~����,$'����нJ��B��A����l�����erώ���T�e�3_L� eߙ��._h4�'=��MP�4)$���]��S~2����֍7O�k����J�xIX��P�D]����������>�!���yF^�����@����Ǜ����';VB� /�@��Piv�GN��>�ݮ8䘛_7&?O0�cO�H�o�א�N��:I5�%{�sVEy�����H`���ZxS@�R��R[���p�֨aT���&��5Ƶ��@�:M���5�9�Jj�]IBn��:OC��h��71@��-8��)u�Z��G,S�M�Z��W���G]��[��x���S����[�]�O����Z��l�3��5��7띖Z*@�Z��Z_p���As+:h�쯗�yTX�?m�=�4E�,�����ѿJR �\����*�UM��I6g~ږ5��A�/��^Mm���2VA�R�!��q�z��}�kzF>��G2V�[��5�t��=���~�E��I:;V� �%+-ߺ��u����cp�s��۽\�c4��$��9wф��O���F�gY�oxz�7�[DZI�B\�P �.�;�}�
�����*�k�nwvX�1�,G��ɤy˙n�w���Ȉ�V�	�>�� ҽ�}��w��J�"TU���:�8\B8�j�rX�?�\|��p��w;""��X�T9�5>`j3�m.=���C�˻����VT�XH�+)O�.iG?]v�K����Yi6 �n�EfW��~�lC!�ɢ_+�S��R�lq |����[Cԯ�=�u{n�gN��s^�7�d��f�Z!a����R�^��^�������������Zҵ������k*�ŌIAGx^���P`'���p�+?Tv~uU7pWWf���:S�Bغ������tX�2�=���t��&<�������,��|[��4��%ԙ8�k�����׸;��p��-�uݝT#�﬍DIJU "@9xs�cRf� ��B��9Џ���(�ꆿ
a�w�VV{��i�1��i�<�ibg��f�go}F9���1*2������x�c����r5	�y�y�x3e���3'�t��X��v��~h�@<�����!�|W�IZ)s��@i�KOޚD��������f?�*Tp�z����<�8�=��\k<��.,��L�Ǆ��p����R3�;ι¼�'�!>./��,[���u�a���tȚߺ�oS��s��M��8Pc���g ���|���ZYCfS����(��"E5e�mCȈ�}%��E�}��� JU(�䔱�&��P���d�� �*e�h����Gu�u�t�+kl�E�L�y��!���9!���`�/e�̡��y�U��X��l��_�M�4�v?QmDt���2c�Ldsӧ	�W�j����"��b F�#4�_|n'%R�Z��	�M�Oh`٣���\��=2��t�"���n:o���iF��1�����$/�=���;��@\n)pu7�PT�$�y� �������^>(1�ĔCP{��z��HI�u��{�G�Ę�����]��������1�X;���MU)�ZZ�B)���%YJk�Gb�N��	y�����<��]�(E-ɒ�R^� ����x��)N_\�J�Ɓ^�ݴbi�Y��k��n2���l6�[�R�_x|_C�=�ŉ3k�eKSYE=�m��G� �������E�ƚ٣��?�'d
L0����m"���Æ�/�E�9)�:B�z�����b���P���9���^������)P�	� �G��r8�[Я9уy��U��6c��QM��� Ր��p˻.G��{-�x�>-6TG��O���Fo�đܺX��[<[�S��$�#��z�ܚ5=�\Ҁt����&Zd=آm��rK���G*��}�c���\��:�Wf�p�/}��p˼ص|��>�@��ts6��Ix	o0��i�Z���'��^���z~ �͡������0{��s:i����~w_�-�a8���@�yJr�}�H���{�H�a)�Hw:#J��/�K��Q�b�~8��_�.�5�i�c&*H7wn��?��%�kS������ל�2��e:Q�.q��� ��U{��p�[��߳�}��G��?��~U�(��+p�̲�<r���IK����4R���\�[
�I��)n�p�Ѹ�S<��Ԍ���W���8���0�iz�@�����%X�
�xޣ���-jЙA7�ɼC������h��D����tЭ+�6�Ϭ*42�ݒX�F�~��>gˎO����P&�]w{�`�.?��,���Kk�b�_^:VZq����z�&�«=:,6��?�X�7ɂ�(�3y�Ģ�gl]���pFۈ�<��1'��N�?{x!t��Ҩ�Ъ�V��:��2�MWq���-��gs�<a$%��"�����(�6��*���=��,��1>6����XsB�ޖ7>��N*�������M�z`�p���Ǒ<Gm�OA��Va�&6ӻ<�'�~{.³���f�[����el�&t.�I��F��5��<�r�,�n�c�|K��>X�/�����/�	ł����kh Xn���]Cг��C*L���Pl���a5���T!� 7j#ǟ��J���ϾX�g�%��<J���*c��o�����B��[U�!~ޭ�-�,���P��!P������`~�^�w���/��	Y�q�Y)�ҚR�����9�Zz[9�T�#��_��I��3N���@ʧisE�F�ñ� ����5o��X���8c�\�\`����~�D���Sx�����חxn7��ڧ��t�֜l��SG�_��ԛ�j{\^:�����9�{�t}l�[/j*���~h;�I�0�{o�6r9A��뀭�g��5u�=�Pt�gШ�ڙ|���R�OV�~\	oV�]7t;a[FK�qz��
�	>%�5EE7���3O�;r�>Z�X�N�Z,��V��߄�Em��S�R6���*���N����f�f��u��n��� a��m�ʋr{���-�ݯ�7�A�EA�����������!-��Y݃�a��[V\�B��&����mE������:�&t����u~,���A3�" ��j��Or��{�3�-�JB��w�u�<&��:b��ýo�߉*\s�ER}�پlq	�7�B�[͔xau}�&�}�y�y2����~�a%ê#��a���y5�����&6K�"�S��a��fW�J_D�ϡ�ӗ�`�e���0��uø���L0��l����g7Y�R<�hAwy�[�{����7�	Wm{\���m��[;��k�^��$���"�u���Q)�<Ϝ�����P�aO������y���T9�YB��o�'�	e�l~OW�.�G����5Y_��`���P�u���շ7o=�ʰ؃����?D�/{E�T�WҜ�9�Z�锫���z�'#t^y����r���� �Vg*��Ap58F֓�]��Q׻i���P5�;SmhJҾ�\�<��g	�Ӧid�7����dK�\��Pr�ԗ	_4����髋��ݽ�?��9�ʱ&�o�󗝊G�+�%Ǜ&�[]��w�Ni��7E����F��A~�ْK���P x4���}���x��W2c�.���3���������˛^�U
��BF&�,b���2�|�rf.���/�)�@�UiX��nʔ�.��?������7��Z���GKk׋�iֺf&[}�����;��?gX���D�N�[:X6� I�xF�������eK����ۀP/#5;JqW��D�5
�����E��}� [1.��ߪ�G���_Gؙ�t����b&g��n~84K�m�89.��5/2�1͇��L��3�G��G�jqV�\��]�tvcA��0��^h�F��qF;�}������a2(��$�%�������%o��|�p�R�O��țoFq��|�f�({���E���Ƒ��a��*n�L���;�yہ ��]��R(��3.����s��"�2����YB@�8j"�?%�y��h��l��t?�Y��>b�N���7�s ~�Ei@��`��R��U��V�)��j4���x�R,�#[6f��)E!k�(�0���.��W����kF�Z��1���9������>�IZ���^߰ )�&���Aݙ]�--�2`��>kM�BMf��$.���N�>��a?�8�	c���~Q|��h�8PS��0N�#~�f����Dm.j����h�+�7����i��[�ܭB`�F�|P�c�7�x��Ln�Ӂy��@��
Y��_�N��k���%~� �My��j��%�j �^?aO�������~���|����iZ.��白���V� ���Z���{2n���Q�{|�xMz��~E��'�c�̀D�ѯ��ޛ�r�A�k��74v������h.=a�g�`��������7��~�{�`��I����(��E�>�+b`�%��4�do��������޶漱�am9����ꇸ�d���ms��Ru���m���[��8�r_d|%\��!��%�HY�)��5ӈ�������@�:��']�O%�����N���u�yi~%�؉>Ƞ��5�u�yj��p�bI���U�8ש%����������'G�8��N�2�[���y}t�K������q�w�OE�>.�h�F��*��i�)O�L���n9I����xi�i��F~먵�R��^7d-��u������jtf�3.�!��&���M���⅙Y�s������W-W�ӨX���(������O1*��l��1�V��`��fG�fNcNO��#я��}�{������K��4y��r�����~�6�i������0�v���f��\|�� -gQ�2;b:��,�JY�V����
a�In�mȒ:*EJ:YD5β�|�\T*��d�V�-��o��x����ǲP�ܡs�U�9V��h<��xЯ6^D:aP�p��U�����0�{�X����+���7pu�*c�6���2���٬m�u����	��LyM��Φ��&d$���փi��R��o�g��j%�,S��P寶y���պ��]�
53]&�N��: iLx�ڔ�Ζ�o�;�$G��F��e�ǰc�Û�V��S�0Τ;��Z�a&Anj�KYV��|X����i;�_w����>�b\�+Vki�ב�K�=�q��>>v�mȬߐ�Q�MM���f�s�ID�^�~�H�/�l7ڷ[�k@=�Ǭ�?���ɪWܿ�U�����K����"��k��N��b5H"��/W��v�}�[�9K,� �INA�y�d���k���ʊFL��#�тg�G�O�Pbm��Z�\][�_!�_���fZ��P�=R���Nm���/�D����(ɡT���.�_����ŗ�y�v�jI/
?���1ٕ�p����n���z,}���3�&�-��f^8���l�#������(� ���G��S��kZA0�z��"��}�$�:ܹ�'*��R��=��E=6�5H�˝`�����u K*�1n��U��#rI����s��sO�3�?Y2[��=�K�#6ĴNQ�<���#��1:r��k@Ç�Z��N�Q�����w��Ύ�a�[�E�nҳ"����u����?�]����,�i�偑:+-GNG�AF�ߍ�/�� ��ѷ�xTf qn��m wb�e�MC�}X�R ��,3/'rQgqm��")\�CPiyfw����e>:�bo���.�m�q�0�i4P��Q�D˱���(�}��0
��S�Ǚ��>VV�ƪ{T�'v̶�m/��_3��>�IEIG�����x��4Z���(�@�4�59�Y��)��r#��n퇜��M�����8m�|;">�B�tI�*h�'��N$9��#3=2�
Uv=�s�y����0Qf<�1��p!V2}�#�F��8�p!���Ud��r��^�vG�8����H������V��r�Yeb�� rw��Qs�1���F�����%����5��k.��o��|��b��K5�ꏒ��ӟ�g�V�Ȝ�{ŦL>��_<����7��7�F��H?��'�z�F�ok���PFvy�)�����,%�ۮX� ���y3ЛH,�ܘi���6��n}P�[�L�2b�����L��B����*n��?�?=X�\��n*q^q���e'o'�PԷ ��@7*�Y C`e�8Y,M�b1y�Tg�|bS�H�oŋig�B<^8Y�Q�^�J���j�g�����ݜ�j�R�Y��Q�a�K�f;+�z�y���jg�����,G�U��W������@��N��Zz�/��Z�TK�(&�k��-���cO��^�e�>S^�o��A�ɹh�f��<07�}?��r������䇚�0	9K�Mv�!���%�Z�`e�����EDE�-��x��$��$���)�7W�nD����#���&�Db�nz�}/z���\��\����ƍ��r��erd�=�kˈb-�Ž����^����3%���AE�f`����6	��Љ����A�mRY��I� ���e=J%Q����~�wv�P�5\� �Ap��tJ;���I!{trI@��Ek��Qu��;��_�Mv���v��T$��͊�B@q0��l�@���5٠��Nro�ͷq�z��q�غ��X�>��QK��Wf�i�JDb���1�K?�U �<[SϹi[׈�fǋvrR����/?��������#5j�fr�r�בD)Q���,d��`���'�����+a���?��ӟ�{�:	�VP.:z-W�g'��U
M�$G64����vٹ�bMj���B�u���%Ύ��vH�vP*��ԁI��rP�iл�p<J����b�,C#�s�"�م�9r��Q��B*|�:�h�a�կ�j�1U��iqV¸��[0��4�/��*@/�'�+���C���~�J���Q}�v��b��W&i�F�ݰ{� �l9#���@V]S[+r�"RcuGhl��#��\���ʯ�&Cv:3�� ����k?��0=>_o(5�����@�CV�E6��a�l7��S�������?!G��i��J�]J�����դ8.�/���-$_�g!���i#!r@���N�$�FM�Kr����������fZ���[߱7�G	�V�5��F�Iޔ�N!}�)'�n��ǝk� ��V�0��*D�Ux=X6�:m\���[�CGl��vo�}vb1�|�E�.Gϩ���+e�{E.1�a�
����|*�y\h�����FQ���T����Q!�9#�?VS }c��F�z ��NԆ���|t�����7P����87Q�W����i�zO�I4���|�n1D9�y�e��|�,��;$%����cn�:N�@Ԩ���q:ǧ>�Ν�ͩj|��:BT_+��
��57�i�,g:>�f�Cv�x�{F��k=_�y(G�O���� ��ҥ``�Lc��g���aF��C�;v��N�<�Yl�b��\]���Z�;�֑�R�j��=U�C	[e�U�ٗr�߿���	�Sw~(�r�Ng��)W|�$zf��]R��S;�s$������F���w�Lm5�P�rp�]��g��(�R���,��$'���|D�!y�g�	��(����j�Ϗ�(���Mv�!���#�\���m�P���q��-��'޻Ӛ=�N+����V��@Y�M���;��ʴY}[�XrS)t����Z�5���ݫp�l�<��Iկ�<�&G�㼼����
�fK��	$�-�
|��o������2�xFط4C�J_��&{�����M�N�T���V'/�J�`���k�B��	F�ҸEslSѯV,-�c@�D��Pl��|V5��Q7�94h��#K�	Zo��Fw�g�G�� \�<�Exp��mI����0#��A�<����	7����i22���owՙ_�7+��_^#W�L�(M���u�c��r=���5D�"���ٝ@�F@��������|���k�A��'�[Z�'�I�Nr�P�{.4D�j �K�2�C�����'��(�T�\%&��J�g9]�~��jv;u��8сv��F��V[MW�;�f�R�M1T3�6R���r9��8[���=�#�4���!��O:�A9Cd��W�1��A~��Ģ�>nϑE��瀍�K~�P�
���ު����=!���/�Y�?6B����efaWC���]`�wK>�E���ռ*9�]�\(��|��Ւ%,��S�}H���Iw��-���%O7+�K�[A�2��vAT���sS�AqL]e���KΣ &�nm�K��)*D9����	3��v୓���:�������zO=C�e{̿��/#�6��h���)ُ�=�9�n��Њ?F)~�,�I)�=*|��f�v�����M��BE=J��4�����̵I���6A�����R�0���uH�4�~V�z�c�6
�_U"[~D��~
���O�-�2�:���&i.kS�|�B�
�0J&(��@)KxD�T/-6|*$��,~�+��MC����³'��Z�[���Š/�Ք -�F�5�r���g�Y�����J�,��-ݶB�G��DV ������֨�4�Yf��I-����Jl�F�a%�WQA�R��3�S�:�[�.ob�N����eSހ˜��=v��3��V��˳��lY� S��4 �0������x:�r~&vF�/[�������t#֍�
��j�]x��9O*#�
Uπ\o&W��������2�<�3Æ�9����i˶�
�	����j�v�dn��K�F�W���:�V��D��e��#G����X����;sy�n�#��E{~�T-����K��FmdIi�Ə�Qш���>+��8���6��UL�AiHV�q(�2�j�<���J1��ó.�D��׃q�t��k����7�<�l�&��n�̎"9l�Vq\�lRHWZ�}�M�"t�/�$����C��V!�r>LG]i�	�Tǰ��=rF�r���l�={�u1��g����3N�'��,��#��N��%����u�E�(�%��*���-�ôL+�[x=�������np��.�6������=�U��r����z���id/�8��s�lY� ��8k/^�%�#6����f3��$��LdL�k M�06K��s�]
�1�|[.KQ�9����s�IG8��7�s��$���$�AX�9�K�Y���@�=#����ν� ����m'������<�w�f�3�>d���a��E��>��U
zc{�o��̱����v��%n9X�٧piGG~��G(�:���L���п0��ċ�3�hX��(ҳGh��D5xj�'��<�C%��V]���A�������둰!<|�n� '�
���"��&���W5����!�i��_�Bт�M��� �hw�o�J������.�E˂
�HQ�'��ȫ^_���Ul��F�?>5"ok�.�E=n_B?-YU�E2U��iwE�ph_�Ȇ�M%4�Tg	���1�0M>@�Z�D}v�F�O���#�J�v6��E�'t?�
|Z6W�[ME�5�(�va%�÷��%��{�:"�#��o7b�V����#$���[�����A:��Z�ɉ�cT�� 
c���aG���K4RJf�8L�e����r���+eI�eʽ ���N���A�����f�����m��t۩t�γ�R��!���L%\yD�V ��*������/xN4��NØ�R��nm��@��2��!m��>R���EC��`R�㻩!��+�����j��k�_o?���-���4�J,�t�o�l�`��H�p�/	j��CD�y��ίԔ���l�ߘZ]�P�}S��F ������J���ܴ�`RP��v�J\����|-��?Q
�A�él�>��6��T�[�z|�-������j�k�>I��/K�o��IA@7�|��p�m�r9P��f㆟�:M㞺p�PU�l��*���e<�����V���D���Ff��.'�MM�}�����i�q�<���4��,>Cz1����YE�\�_U:���'U�q9"f�G	�1r`H�V~7-�N��2�g�"��;k�/����V��uX}�Lk��Rw��Mr�obЋ<���jZA�s<���_E�g�2�=d��8���D�Rs;���/)�0���%����A2�v0�N��� N|�%rs]\���Fs�v��A�.&o�N��ŦR.����qΕ��T�V��u�(�ш�Rl�Y�f\�v�Sq!M�3v8l̈<ig���Tg!�_�$���������
�-]�L(�GP���F��KC���I&-��ɭ�@O�m]�,�P޾!��=I�T�޺��v�����
 ����[��̮u����H��{ڟ�`�PǇ�˝��Ҳ�\y�:����*��v�z����������l�ֹ�zW�wƘ�I
��p;8���I�OP�Ty��XB|4�nǳ��^#t!�t�	O�LW��1�¾��L�Fz���V�ÆHPl��@D9J�.M�aκ�/�GZfÑXN_C�`p�l�gn���	������yU���Ǒ	�X~�	#'�EabOl�3�۾���k�j��e}�hH��阗Op��i�>�*�R��B�2��vdU1��	yPO���4�M��O���W�(�Xh!v+�D��M�B�l�^w��+��Ο���-c��K��T�d�i�7Ҁiu謂B����3�5LFq7e��xr��.�1��Re|��YnnEX�8�zjj2�%�!>�%�^��p�!Ŋ$�Xa�%'���Ȼ C���9{.��+�!�6�ۺD�ˇVh�w��j���ޟ���.����x0���N7z���o��(��k�������w	xp�";�!$ƖE�o��7�Z��e�J��U�wC۰�2��6���Y����.Y-jU`���K��WQ�3<�l1$"ׄ���P�ߢ�����;Ap6_sĵ;����]k
�(��;�>r$��������YC�bM)���B�)k����`�4*�f^/S�U�J+Ą��Չuޒ��E�x�����2�ք���m0�jy���O*J�O���$0���Xޛ�Q�إ��k�9�:�Vp����
G���d�H�������D�i�)��Rn�t�Y($�7�����8��a�4�Y^jg@��_K����J9��[GvS��]J�g��[&�Zq��~;��Y���o������h���-�B�t������x�z_k+����?�/Ii���#}����F@�]�N~�Ss,}���Z��E�p,.��!M�^.���p�Ő��gdf"�]�� E�4<���?ԝ��9�.���vh�?������99K�8�b�H;>1'��k�,ʗ
z    IEND�B`�PK   t~�Xq����� W /   images/6b3c47ca-37ce-4ada-891d-054e310e4230.pngL{XT����r�����ݝ&20#��ҨD��A@���!�[��Az` i��;g���<��8μg�{�����9|PQzFz��*  �0�'� @R �N_�fǁ� .:?������6	�}�A^� 蚠?�-���7�<�tQ�7sq{�d
����X�Y;�r0�w2Oڐ��{ ��C��qS�.�{�����:�R.�X.�xE�B������*-�l,/Hu��Z�Z���sֳޏ=BQ�vCI����JA�V(K���D�0yǿ/$92Qv׌n?��\>L�5��wن�j[g`�ά�[�o�n�y�e�����{f�~���țGѬ�7܉����Q�ϲ�!P���%o��Q����0��Λy|�G�qN켖mk���v'�$]���{]g-f:2�1'|�yH��J�feJƑ_:��yY�w�L���x5���P*٭��:4T�c[�&Q��K ����rj v���8��F=���i߸y�L�y�J��0��p{�޸�a��ԭ����E��.xj����qB���O~���?�3ؗױ��z�;T�n}�S���)�cv������!{;�I�Y����N-ͼa�w�cV�*\�hݛe5�������������jjj�*#-Kl��(Q��B�ucrQ�S�A.����\��cR3Նj���I�Dˆ��ΓO�d�%D��cn�c.vگBnL�֦⳰���c��� ��_��bJ�����s��w�I��� ��:��.�tOY�&���;���9�>z&~r���A:q�n��r���՘!n�8�WSi���4w�T3�6�ε�`��{Lմ�		�"��a���q�z]��Q��VAS*mR3��h�/t�Ż4.zN=��8�0�zmϰY��w}bp��D)�_�:_�O�ɻ�
jc�)�n�Q*X*'��])'�j�`֥Ή�'���ea`W��O�ιj���
xk��nd����C���1��\S���c��j��Z*����4Ge�@o��=O2��v�R����=-��jdg�೙�n]���z�D�q)����Ȥ�Ҽs�5��0�q.�-hR����V�-���ڃ��ŅM.�)�-1*U#;�ď~#;��"]�1�o�'JG#�EMi���JS{֫�AH93�,E�K�	� ��|"�|��!l
%񼞳��eB��yD�I�Ts�nf�L����y@�&���k4EE�k?Z�a*���U�iRj6�������ꔨ�AO�(i����_.Q��0"p���D��Z++<�PIH^{H��Z!���>h�2��0I�	�d�5Sޮ�R��$��ےnޞ��Ƚ�A�*��/�3�J���ʀ��G�=�]����0VX^�ǫ4��<��jܚ�S�;����qP���;�-���v�x��j�����KR�ğ�{��.H������>$���ڥv����N��RJ^?�u��)L�����:)!51A�Ϊ(˺+56��F�L&�G�Q�n�x�
V�ZI	~Ձ��
̇�B.�����we�Q֑�-��I��a����,;4��q��(�&����е,�8�;L[���U��Z3ā�;����ϐ��H��O�@�O�9."�<���7�};����3�Ӧ�j=��C*�CM��7j�{���a����%�S����{�_�Dv����]��{W%Z�>��(	Z��z3��$R�ꎘZR��Y�3��o͞/ko�I��Q]ހ�N�c�_�c'������mgI>vW�q�A2���g�]�Ӄ��>��A�����OѢK�D��i�]~%Cb�p%7[�����Xd�����ӡ�=�
L���o���m���2f*�w/W yǯ2���&mk�߱� {CaL0ys���������B
�L��8��ɿ�s�\���8����ˇ�a:�O�0%��pk_�&\� �-,u���F{y�LQj���$�UԱkZ	)�ػξm�^��/�[K�1n?o�ٽa���z�g��IFy�5���!F$���2*%�侳���X�IϙuI�g��>�����䗆uT��nfn�J�''Wf���+�o����������gE�?���S��{��Uw��8��8 *���$�3��!�d�Z�b]q�qJJ���6e��T��<����2��n�_�G�'�~L�@[�D�kXMԈ����d|�ޣ�;�۷�ɛ�$N��)���vǞH1=��e<R~|a������i�߿�Fa.��ށ�Ư�˫��(��L��]�-TІѯ���B'ْ����N�;��������U@T��RE�䝚��x#�D��~%"L��(_ި��	�n��wP`��+��R��k�2��4g� l�����Y�e��2���v�Ab�vd#�)���ֺ�g�(��<�N�O�+��҃�f��$�9�,'<���Ӈ�^#�}��ôJ�3�ޞ�mz�C��)'���)#���Y|�ttݜg;ɴ��Ԓ���P@�����
͒�N��v����iѤ@�Æ��fG���g�����чP�j	2[��e/�4��q���Y�L�:�
�&��a�2��U�yA�-s����s��RK�Hk�;𧳉�fJ�fo�#�㏀+μ��X{�#x��j���r��Dq�r����f0!o ��wN҅��{Np����,���m�_eT��'�'Y��J>'��&�ԩ�>�	���6tK�K��RB�}�JB��E�L|h#*/b�EuX�[;��Z��v��)�+��bz}Ti�ۇa��u���>���2�������0p�<��sZCo��uq4��l�~#1a/���C��.�<{��h��&���<��qpDe� ݿ�
q��F��x����nWO0�q��#� ��zG:�X�'f��	���R6?��2�B)�_��{|T��X �ĺ�VY�&�##�����($����H	��w��4������6F�Թ�=������kj�F�P/z��f܋)�����i�J��F�b��g&�����Ϛ�3�kX�7	�SR���lU��%U�Szpi������`*(�q:%8��]��["��]7��0���W
�1"Ɂ�!��j�Ό��A[Z�gF���'���M<L�i]�^(y���f�z�˙��~La�]8-R��fȂ|��e3��BV�k�`�=`b.=��J���s�q��܆,�����A��$�G� �	�9�tn���!Ǩц[���7s������#%A]�Fq嬗vdc�2�� @I>]�%��Q����_4%v�<�~%��-;k���*�K���6��H*`�[�ޠ�l��R�Q;�1_͒�@�0�`�����eBD���e�>C�V�����<+|a/�ឌh����Q��c� |J���5	�A�g�H�Rc���0Ȣ�c�f�%N�=*�����ؔrNxn(���E@}��f�тWV����q�@2'ٵ~��,4�"�:��E�I�8!'Q�����wtt�a0D�'��B%ڇc�g��T�y�;��K�}w�]��k�}����1o�n�U�j�ʜ/����bZf9�go�g���350;zM�c(�e���{Nl��w��268
{R�iW�{FZ\
�ߵQ����J^���ϣ␡P�֗W�X�{���t��с6-N��[}��S?���H��ȳz��4��!�8���`P��. Y�JQ#L��L���P_��7Q���H~�J2?cʈiO����eZ
�߇'v�S[�xn�ي�c�����x����:M;��\��\���a��H��'΅�N���P��0Wh�A�lX�⸉V��A[����BJ������o��&�("?(�	\.� �(b<��o�r���jr���'ߡS8��Ʊ�b�u_�O�H3p��8۷��&oH9�^Y��˞���(�� r7�����荺E�bc�cY�t� �x ���Ɔ���E����p]��1"���hzO����+��\N�0q��LP��.�� hҟo��i9E��������W�)�a�9���(*��8�E��1��|c|�����MB0�W�PkC�Z?q�=��<�o�cs#����J�,��֯��J����Wx�Tyn�qk?ӟt~��{�^;`J�*��c	�����0�@Z�cT
	���k�ޔ�:�7�n��+x�t����)��pJ��E_z�v�L��\gpu3�x��;o?��z�y�D�a
Z��|��#k#�Y�Gջ�0�e��e=O��13%BQ�rs�K�����V���� C�[���M�a�(7��ŷ�)-~��%��XE$l�>L����3�ǃ��zۭ�O	;���c'���u���dJ�m��m,.fAf��� ꂻ���|m��j��ۙh��t�aL��B$ge�ƭ��7��.[�������^��N��^��A��а��5C/y�^#��V	Wh�6�Kuw�1`jXtۧ\|#fz��q�m���R�@<��g���>֟�f��}P|�FUa�1��M�I�a߯gp�FJ���2����#�8� ���ꡌԵ���9|G���e)��QA
K��1�b�P86{�6g��oٞ"�'u���E�5vv��Y\�խPM:1��9&�(���J(�ݚ����uY�Gz4�_O���E��Z��%�G��L�ov�C��K�O�2��3��en��zF��5���V����lx:�5�o?M}A߆�6���i���;X����	�0��zت}�e�ѵ,l�u1Á���/��gSY����F�M�� _
Ul��x'��B7A  ��J	g�S�ۮ�R�7i4i�4f����bj2BY��nT	��.4|��nR�.�m�4=�0]*=Q���Z�!�fF�d>�T�Qg���d,h��~��%H���Ka}����G�*�ʬںq�9�V���W�O��)�.:pR܏��Z�F��k��-p��@�$U�+�w�	 ��D�U���H�d�/,k���*N|fd�t�g*e�y	*��-��s�Thhy��o��p�պ^s~�]��ܼ�w&���;;��=QSSkz���Ԋ}VQ#�Z�X���%rG#���m!�b�9�1�p��da��q= ���%o���;QH ?��j�[F['�X��.@*k5��l�*c�|��Dzy��^h�x g�-��np�KBF�ƌ�]����n�;AS(!�YZ�M�Ŗx�]�=Y��`��_�u�������86�fQWrZ|�C��+t �*��n���P=h�?��vǮ��V���@G ����xlQǱ)G��5�������p�^%�.`�֍���\+�Zh���t�b�x��"}�v��&U��i��~�T�����M-z�.N�'?YaR~���V���8�
N�<>�Ͻ�fn�29�(MkY��C~��`BG����V:Si�q������V@�d�M)t ��Zez+\�/�ω`�����}�E�I�D�$��O��C�v��sg�`�=�R8󾛻��3�޽s��Ux�����[�M߈xA+k#l�^2r���BY��3z�l9X�uk�����1'�bX��X+�o���=�sB碍[E	�BL�qq9��0���ea� ��_f��p��v��׃��d�	A�AoЫ�����%�T�f�M�F�ڻQgX�ņ�����!�6�b	�.x��l�B��;
U�q%}o��2�~�������'�2���b�.�n��c�d������unj��5C�ڮB��"�ĥ��`)ĉ$��kMȲ�DB�}<��jf��d0�$�B~��f:�9x�ҟS'3�4B�웄������n�pB�îMswW�_�U����޸x���:��>o^���'E/�U�(#[!� F!��UFp"�������Ì!��l���%@�	R�4!.o��f�m�j��ـ8!�s��c�s�.�:�<B�������<���tA�e��Ǌ[a+�2	�B~�����@�1���C&� s��DݧeA+�~�<��BnڰK|= �IL|S�bu��ܧ��2q�}C���0e�6�zL-�W/Ŷ=M	PdB×��B�A��==1n"����PW��`1T%�L��y�պv�nZ����"��ί��g���{׬�b�[���j�U�p<P$8��ߘ��Hٵz^ qbD����p+�*�`��r�nD�-��ःi��>�5c���Oԭ>�:4u����چ,4����c�Z��*j5	!
v:�QI7��5��Jn�1����CC���0v4A�������rMM^���x��pnq����E�M�)C[?$L�/��_A­���_�Ы" UHC{SzDt:dG	^	r(��V��K��Jr�~t�4g�}p�?_965�!�r#��_(���m�ؙ3gb����rP���56�7�t��m�׿�Y,��ng�!���@���:'�"�����n�~Y�Ա��|9q'T=���,�K���6fP_ġx����0rE����|Z*��st0N�� %���#�RE��V3�pp�����C;�� ���D�h�&(T���@��s�08"�&1U���u�Q���@RRF��O��_~�oW�Df�D�&_���&������v����k��B��'z�8�S��Õ�S���o�gs�>4E�g�{�����Ξ�|$sTJ�e�i�p����iΟ#*�a�	I��6�3
��X	C�[vط�	C�GbJ��VĤGW��3v�(ڻ˨{����g)q�c+7�͞���H�?P]��L(�At��Ԧ�p�%��e�Ft���\�����L��8�^	~={��m���Q���* ��'��y�ֈ-��Y�*\]�c��Ƙ��E�̽�.l�f�<�a*<�u�������(��nOI�=ǈ]��W�+��=��޵8:W�K������slXoF�-d��<�y�^4�&,�3b�E�ġ&���O]^�����9�'����N��A)"վ��u���L&�7�2ݥ�e}X�l��K����^F��FQ�{&LX.�
v��=�V�fY�Tc�0���3�0�p�fe�����U�$����Sx�^ݳ©,t$�C8~g�|��F)s�@E>5�;���Q���G�3w��e�M���5�+�S��岴`�.{��LݲA�~�+�St�r|ގ� �?��)�	�:3�=ϊ��¸����8�B�+aԞg�߷�!�D��;���\o_��Q�vOt7-�֟��&.=)���^Iw�w�νLE�n�P���'C�v-"�{�ƭ��*?�Ov�,AK�n>����}�PA�+z|[�	�����n��&%�x����A@����;�Xmw�� Q��������K �R��oJ##�0��i=vAu٘�q��m����Ր伾��]Y$�E���2�%��s3|���Z;_��ҙo1�����t�����`L
k鎞��eEP2.��f�2q4�u�a��Hx}��I\�q9��E�XtN�C�<��u�^N�g�I�ə�A��3v�X��	\xE��*�+j釺=�ha@�!�J�A����p7[ݭZ)i3,=�s�s&.Y@R#�/��s�#��8��^���?2j@WH/�A:�O�}(Ҭ�D�NO���E���TQ�w�����`[�0��M�[oǜ��#�N��a-Em�0�f6`?���J8�\ďSɞk#���}�+Ty)��s�� ��m�.憻�w�:4x��Es�a���8&(/�/��*�1��MG��1�+�Mp�p�R\�a�L�;��S�Tŉ���	����st}��=$5xy�~����+Q���K���.���]����/���{�1��D��G�m�La�G�C�杝���N8�D��-JL�r$O���(;ty1��ݐ��A5;|�=iq�b���d	vͼ5t�; ��2��iP�YQ݇r	���⸋j�Ss���H�X�{	H�/��r+
b�7�N��|�T�ф\9{���;��'+~2T���9�,㙩-�=����\2h�������rƎJ�r[�e׆O�H�ljP�3��w�~����M��{eYE�����/��	�Eb����{�6�Ho������+5}8�l"����n���铔�R�B�;���;R!�!
+�e�6M����~[�mu|��%��_�t��m�������Oܽ��q��
$0��H��?Ѽ���p$��y-4cuL�S=�~u{a�VW�>�z_tgl���5M�����$#��b��_>{o��	��
��U�^,�u�U�����|����Fvt~�eL�J�L{��3��c��D{� �1�_���u��WZ�n�#��Ou�lW��~�ѹ���<>`o)E�<�+��|�H^���9!�7R*~�з
R�=;�A��*��0o�8�$4���Yp]>FjS�勓�3�ߖ�j�֦s"/�+aI1]4�/R�V��uƷ�ܹb���=I�m�)��H�����:�͛�Q��7�i�E���n.�RE�C۵y$x�{dQGL�bN�R~y��8��rb  �?��)i���z6$��N�P�mc����."�)�⥡+Zv>�!5;�nh����"F�I^^R������뢸^-���Q�X���M�2q�|���g�8��a��OO���lK��|s���Ƅ��`o��J����皔�1�T�������E@�	~�KI��Ч�d@� 5�9��~����F��/�²�g������Êf��wJ�y�wF���󯟅��!��dB�Ǘ���3����:�uT���>x�bm��{TY��iA2j�L 0��`���X'Ƣ>��fb����bJ)R�щx��]�l�8��T��Ưcݴ ���(yV1S���׷K�ꞝ=��pB���K��+U�e�prW�ho�W?z7���P���wXW�6�M� �����#�\�%�,5=�1���ӛ���;�y�SW ʘ�x$�!z��z�M ��[�w��~��X�;��=���f�gr?�ӏ(�'UI@ǪU�������^��'
�&�3\����1��q����q�&2{$��k�XyW[G��y��uD�'�۵����S��\�������!+/�]���K	�G<l�ǽ^�MNBI��H���y-�V�[��/�;���~���]�������#��$~̗w�Q�`��\W�Ӈ���#�k��eξ�]�f��]t��#����OI��?��O.ո���P�d#ϝ%�Te���슾�]I��������z��M�7�V�V�O�X��J�H��wB9L5ۿ#��M������>���Qږ�����Қ!�:����53O�
���Z���z̻����i/��Rn�����a7�����3R�+��f�tT=����6�TL��6��Hˊ9����ǧfz?;/����Rd7E�R6'��[��%����k?9��W�ɋ2�F�mi��Q�{րz]%̫��[�;6
=���؇�ƔiJ̀k��-y>ΒN�^���|<Y0�x�/B���@� _�y�ڥ�������Id&b�;�m�D���":���פ�� Ӆr��ՠ�;�w}'��@��2Qy|Q�x_���ݻ���A[7��px���v8 '@�8qLa�S�|c��%PeX?y�z��]���Sן)�Yiz�3W}�+�]�Yu�8qpiږV1|3� P���U���x�TZơQv$���7ln�RT߳���\@ؽ�LX�U�W�TD�V�%ԋOR����eu���)��@�ϑ���j"�����e���v��ΞM\�ۢ�|�e��o�}� 4�[�cu]R=�����F,�
H2i���û��0�=�����*G�cz�È���0ll���D.�`��}������216b�ُ[#�Ջ�%LO�	���K|�ۯ>-�;�]͕�5�q%�d�椕�D|�U��H�ʬ��Q_���c�h�BJ��8p-j�ѩή��1�,
λ: �T�9��wl}�h���D��RNpf�]�c�2���U���)~�Gmw����ۢ�!��/��;����QW	�$:����ώI���wu�_��[��N"r?奟e���H)u�U�H.� ^�b��ۓ_Q�)a�b!j�-�fl�R#�h�~�.����_�����]��t�f! M�%�I����n<�LR�q����'`��+�TGtt��Fۤ���0��R��5�BO��x?2M�2@D��6H9�˔ ?�6=�1��~P�,����O�W��)Ko���$ ���,}��l��.~I���(5��zG��^Ӑ�`��Y43!O��[Ժ��2�Ǭ��a�����h�#�apJ�G�
����gZ�T��F�bW�9��{��t�#D��
\a�Sb��a�zx�@8�� �E�Xa&�f��'|	=9]�#!
r� �[Ǥ�+�%�dfg��`���&���O�@҂;(���f��)V�n%џ��Rs2���S'?U�'g��ǄL\0DY���.��,5����N��T�!��3Z�lc���Ih��y��9�֥����p�0�e����v�3 1�]A����C*;�n�M�]QS��U���<9��:CE�A[��LKl���6o��ǟE�j�[��BC+�Y����l��@<��D|]��)�Vծg��}�؃EY��a�[����D�+�7Y�})���ƥ�{D���\���͚�W�|����}N���%� 2@�G�'Y��
.�$j�@>%���«��bOO�������q�Pￇ��"�ʡ���L�naY�1"�n0��X}��̏����/�ư*�\��d:.������d�oN<;�:�P�r
=���t���
8�fag��$����I�|g����<����vp��	/�x��Km8��C7��I��� �,��8���;�?���z����-(uY��Y�D[���j�QH~�iʷ�R������б��tu����](�0�w��s[k��c�b�?��T.G\Jv��M��N���рԞ[�Ѣ�&;���8>� ����?a�Āu�-X���g����X
�3:.,ݖ��j��5^ZJH��>�!O��Z�m���!.d{.�VH��*���k����IS�㉆��+Ul�n�}], Y���j-K,E�r������[C*�W���b��x7��C�_�HqsP�
�~��t�}n��SC������ڞ����o�Zڵq���iR]cao��T�׎���YyW�G���~k��+(|�;��0OCQ���Կ�4`⮞�BB�J�ջ��*�Bbɼ�~�j�a�9C��؎3\���]�U\8(����s:�W\�h�Y-���.��Aq�{����r�B�yyo�`��}�	�-*6��ox�R�{k���}=E'��΁�G�-#�s���bI���TC/�4�au��]U�X�ڧ�)�!k�c��~���p���:[n�� ��C���p�كk��Āa��i�V�o��!�1����}r�Z�� ��I,��Ҳf)��7�W�������j\CA^h|2��T�-��Ѡ��p4q.y�Y�GT��uV���`���.o�4�����8bb>�U��$��
O51��у׾��j!y��#��5���]j#U-7�>C	��xv��=z�S"M%G¸�:'[��)��:� �5�*"@e�
o1\kxD��m�a|'�
B�z��5Q�1I�T�W�0�7����x����5�:d�n�~��7�ҽ�t �[����I�s5l�H.ەo*�
JK�hTuM�ø^�2�`%��T�t���p�s�G�B��_(��iB_�=�ݲ��+��#	(&���Y�C��	ٷ�;]>]�-���!�Q��1|��Jl������#\W=}���"{]��:���%dc$.�Q�;��i�'�|Zy66a�@�(w�IтS4��Hi����,���q�3���f�+���M�?�~��D�t*'��8Ik��N��[�*�n}��w�����x������H�C�*PyV��s���EU0t�����ӗ1�c��J��ӐC!<Nj�>0O��:�\&D1��q���<�8k��׃н�OW�݊6�8�;d2����z`��j��y_f� ,d���%����A������+����j���B'ǐ���ҁq��d��4*�'�+<d�s��Q���Zi������#���E����Bx��J��^�l���hv�)�u�5�V��AA�ؤ����U����߳�Fp���~�җO���/�����n�A�,p8��8�F����S�tq�t��Ә֙	�9l�\�\�~��_�R��r�l���_��]v\��/kk �o߇���h7U�s�t���:%�˳fb^��d	b@�*�&��y���d/��V���꼶i��P��=�@O=\)�~f1KG���s���s,�!���
���R���P�TwJ>C��9�4�;K��l{��p�� %�����Ť�\�6�\���k�i�EO!iw�������3�U`v�
�ν`;� ������4�i_���h:#)B��A��Al����]g�'G�C�@�8��%����q��w=o�ڤ����J���躻@��v�)�m�Ր���6���e���N�D�R�]UIj����K>u6Х-+)zb��{�0f��tB_��h��!�M_C��=����Ļ��8s9�5F�pڼ�m�ӯ���!n��l *��xrЕd����N��d����hi�v~?*V��j}��L>Gn���7��BT�#��VH��y��Vfj(��mE!�)�S�^e^�� Ɍ<R%�{s��l�n>E\�19����5���
���̞�Ρ���\K�7a�_S��v�ԕD!5���Ύz�0Q9]lȢ'-��d��#m�������Ò��I:����m�tԫI�7�m6��P(��V��[�����%Ri?�������'|��W�7��}�4 .=lv�W��=yU���R�}�=,��W#%g7�~M���H	ӹ�h[y�����8B7��W��"zP���>|�1-��⹠p��T���B����5�G{M5�
��Z�!n/���E�L��4�&�\Ĥ@�ɉ�S>�0���#�'͈ا�����hb235���v�w��K�Ob��\�r6�ݰ� �W��!��<yN�b|Fά�|�>w-~�h�;�$��� ��{u�W<��>^�S����>��5������P���V�-�x0�׾<�����}�]@p�w�	�����w=��8�+19�K�ļt�:\E0��T`�CM ��|�_����G?s�r�ߊ��
6Ky��_��%oH�  ���*7���E�X4*j����X�Z"n��UӨE;Qj��Μ�7���-�1�� jE���C҇&�[�m��� '�觘�۵��)@�'�J��ʕ%��Q��%�Z��X��X,��h=���*iHM����Gy������7���A=y$Hy��:�1W�(��f4�M*(�������E�Z1�tQ�ح�|��:�o���\i�hT�\�b/�.�T]�
�����L	��ݴ=�\;�2i[���y�Q�`v�@Vm���Òv�e:[jQ�h`dW��r��5pj�޾g����q�hHݻ�4�u]7�g��qFWȎxVSwF<0s@�+7����ʓ�uC̛�4rc�v"%�g��H�A�c�9���{���G��_Q_"��%������Jc��[;���kg��/F�����y��S���	�1��^�!H9��u�i�i!�/�BJ����'o�l�i�[�]2�?ٙ�bw%~��Ik>6�2��VN��d���-���d�͵ב�R�x��opI�%ƹ��)��ѵ�}ފ��/��8�k��i���c��uĶ�	�O������ŭ\���wM��8�����HEB�6�8^�+|���͙�g�E�*��;���ؖ�ɂ�b�f�
�Z��u��c�m�t��B��+���6��̚��}_Ͷ��Ӫz��Ѿx6O�=75��"/3���8�뾐P����4���R�aެ?G�)˶�98(��ۺ�%=�����m1ISU%��`���� u���E��2 ���wn{�grR��3JA��֍�@ʭ���T������|�x����Hf&B>�*˞�>Q?c�*`�a�P\�w+g��B�lׁQP�t��fv���m�S���>6\=tU��ר�ˮ����-�NE҄����%L�ס�%D��!K���ȉx7DK�Z܃�r��Q����	�)I
ɂ�x�g�E7[�0�,!�:�	��(�\�i�ָ�%�*v��F�&˦���W^�"~o��&ow:?ڇ?i�����o�}�e ���]��Rv�n��<������ZQ���]��R踲v�p�N�����}�ˎ[G��H[L�ti~��� ;���Yߛk�x�C�:���J���d�8�6�y��,Zr8�!�Lĕ�E�� hd;�3צ^f��<Įr���Mn=�Dn==+/���XV����G�3�*"���*{��`	�4���g����A���,�K�.5���������[I���L߽�8�kUB~���T�:�ne�+������C�rjҸt�����V�"J=m}>�Ekn�����SC%�6W�`�3D�� *��YI2~�E�֏�9]C��A%��Ϲ񽁿����F�� ���p���qN}�6%�@�.[cy.��:>�*��'�����HWQ���<�>p0s����f. �I~�=�l7�zZml"4�!Ib^�$!Ƈq<\�(.���+	0���!\�gOL'�6-o��/m�M�-F��c����m��$[��ɯ��%�������p��/7�3�㺇���b_�����������A`�����M�-�0[wTA�����Θ�H��-�'\vo^��(��g�������I�@�*2�^�I9�d�Xe�?��)��o�V��6���g�]��*�	����\�������a�,��lڢ_%>9����!-�*�Ƅf�X��U�`-��<}_��j��	�EV�^C �ث�4R��P���x�{�4zxŠUJt�ϳ cY>%}6��7L�Y��
�[٠n�pn�����JDŅ.3q��d�=WzXen+j�+ٕ�[��awfF��v��q�?�o�|A̺jF�����>�F��纨���&�t�⩬k��5E�޾Ԫm��i*hWQ��|XD�ۿw���e�g�d��Nj����"öT0tpz���}}:n'Fm���,[��9\����k�۶��"f�U-}+��/�k����?,�N�G.��υ�8S�W����j�c>Z-9�y�ߘ�x%��ʼ���ti��zB�pS���N��rg����\�l�A�#�%_�غ�N��iK<��]_��وsɘS�CV�g�1��C�(��Yb@;�RڃIY)�J;T
��3u�:M�	\?ʘ=��U����Ax̚RGm=�Q��e��Mޮm���a�����^��B�8�C���� �铆�%٢<��5�/}L���h��']RI:2RQ*(�@TW���uq�	��_~kSV	�ElY�����#!j�U�<����֢sIHUoH�'f��ԇ��r�AN^�kg���ӝ���%�k���q3T_u����M��z1<�	�4�n5� o��b����냶3>Nn�Uç�׳���5
[�J�^/�BRF�s�zc'��n�Zq�M�`�3��^Q�{u�1�I���E����Y���c*M�5��:�+��u �~J���' �<��z����~B��v��-͛A���b�(	"Po@
y8�/34��A:���ׯ�/pn�����-��G����%�F"��ǋ��	��k ��G� g�\5Jc���f���.]���|�B&_E�=���vm�1�p��T�h�k �����{%R%�.ꧠ{����#��\*��A.��u�D9��d�䧇�1[7C�-W4?G���RC �N����3ׇ�GH��2���"wT�Aߦ9IUL�kO:v�������ˏi�'KO��m�n��{O���}6fW�#\Q�%^��d�hB�];�N��ݳ��S��������������؜S�ě����wM�։�����o��ٿM�M
r�����R��[$�^˿�Zl�՗M�m��O����b
Q*8=2I���r��ֻp�b曠��X�H	O�!?0tR.0���h��PXLĚ���ņ��dG�zwH�{���5T!�s )NI�<�	�Gߨf�Zq_Ah*]�z��.]FQ�;���9�kL�����kl�$#?j[�.!�����摫F��[7;��5l�����~px�絝���eK��ޠ�m�~�-�4��z�6;	]���W���'�s�)��6Ϛ�K8E,@v���Y�WׄXN��>ِ"1�};7�a�����~|'��. �&|j'�/�V���&�>9��q���\��F�=��}�_u]�s��/��� Gɡ>�-�3�-M���?5	E>I���l��kR�A_a�6h��/B����Z���p��!����׿qN�7�l�V�"�pL�:4Y��n<�N�z��@Ԯ3xV�����)��������m�X[-�c��f���%��5^���T3���m�^W��F��.��3V��1o]�w���Q��K��iy����|WI::��1F8�a��8<ىm���l4� �=��*H�����z1��5D-�}𚝴����u�J�1�~��ۑϋ4�j:a��1sD�r�6�qK��7�D���r5�qw�F!�j��^�S��#�K�!����m�CJ��sD�/燺l�����a�]xJЌ/��,�߄�,eO��;<�ܼ=�1v��nT����R"����� ���~�<��]7���]��0c���*ڸ�h%:�H���׫4��c8�MϞ��=u�N�6��<�D���xo�/�7fL#���V7��ģ�^��?�����R��}�'j��K��3�� MP����0�d�`3F���Aúu�o����X7�7�>(u�[W�{u�Ӟl�< ti��j�B����7?вf�JnM�����7�����Ö߀�͸,zg�giw��lX����-z�Z�8��l跕 1�9�I2�p�ޜ�}�iO	r�*��G�v�����-t������o���v@�r��9^ԄO���=�1�u���ے��*��$'f�<��)���)��-���Cw���8�&��ݓ��A����W�wM�Ӕ�uz80�������V�X{�������� 1�P�t"�Q2����e�(J�
��#�@
�+�lP#H/�d?��d�i׽���WJ�~�^���`1�#�:W�,suӼw�g�q�(dn���i޳����L��~"/qi�{ΆUf{֣,I�鵙�P�}[�=h�눽$O�J���Z{tlw0��{���;Y�<�Z�dC,�tZ�^9o�P���.4R@�ִDo�׽n���ؒE�Ň{{Ҝ�g�D�M
��[@HWp�u�`B�Q��u��w2>�9δalG���/ORk��8�}}5��˦Z�rf�=K��9|������c�ش�<��#W	��Ĉ��̽gTUɶ6���"�D�� F�*Aɒ�h $� q۶�i�`�HR��$Qh�H� I�H� o��v����{}�;�m�Ԫ��Ϝ�j���WGl������=n�KY��
�w��N-9�n���z�������rZ&�ގT����GVd�	W��w����v����'8N.z��L�	OGA7
x|z�`�,�F���8��Ʃ/%�W���6��:o]�����ȧ�,p�j�Q7~ey52�7����.v���6GP�{��3��OT�\(����ƿ���`y��)��`i�m�K=���<,�Y�k|�;�`�W�n�7�׿�R�W�/_�������E	��M��e̠Q���o�(>4�{J���-9���{K��;0����m�;�7l�-�=�|��|�}m�&<�F*\��Y����)�"�Vt���W����G
�6�Q�c����#�7s��y��"gc���5������v�Nrv�;��������(����J]�}������hHǧ�I$�*�3W����(���>�U���FeTp��x��Y���뜲�Pl'	p����ƿ��&��	`a!�q�D�Gy5݉�/v]�������<a�ߏ��'B��,�~}\}V?�)q2�-��5�����Oݻ��ڕ��ө�h�@P-�4qb"B�G��;���BV3N�F��\��Y��ݯR���:��;x�<��@E�_֓ D�+�6㳗�:BS�~#�U<#�]�ݲ7�ެރ�ΰ㸩v�������j��u��P���#���s�[���[��j������@�z��:��ڂ�֠���yyXj�`v�L��x�Ŗ��y�g�cɒ\����²igիǿ.D;Jr������\l���������̘Z���*D���MJ!̎�����ߴ�_g[�{�T�.*��ظ۠��wȕ��WAH=����o��ܡU+v�K6)%|�}�,5��{�� ���ї�ʹ�#��$ i3諔������(�KOaJ��,��ϗg2��?Q۷�e
�Q`��iӕ!�MlF�NV׎�s���qr[�G7Ѽ9��-_����|F����A544��f��W�A�yT� �{4qk|Y��a;�X���W�+�����_��pN��n\���i��W�{�bӇ�0���c�r*4͙,!VSQx�N�V��ـ%����j����*悍`a�o)ט�|MO^P�6�Q� �c?�a���3���m�Mǋ���k�s��ć}���_9��	k���뼙�[����S9�VM�b$��������Ö��z���;m�����ưV�|ħ�K%�4[ǧ��h�W����j�A�-����&*]��	�c�X�K�tF�8}E�b��e���3X�~��G�֭q�#�Y���]0:9d�.��� I�Kb�)&~O�式�҄�u����JP/��~�'K�E�e�垺���t}�]@�*ӫmt�s5�n+I��'\\i��H��?����o.�����b�-�M�{}�?X6�	�(�h�0�
��a�~���KZ¦�V��n[�7�)�أtX?��zJ�7�Փ�lΧ1Vm��q��?v���2���{�y��gh��f,\�^��ǔ��v���C=#�vb��g��rg�=�0��g��q�1�x��O\ҋ{H�z��~v�i'�>��,l�񎮐}U&��&�<��*s��E�Ĭ��V,�d�j�%���������rE����޿��ā͔#8$�
n�����.�{Ϟ��
O0z��a<��S/
g[���hG��wc��̑\���[��u�~ob#�z����.�/�T���L�ħB�0Q�vP���_y_�������W�u#����|i���i�� ܝ�#n'�&�pt.B<���`�c m�d��`?{FOp��<�t��o/4�0�=�5��k�K�TL56Z	��N��ɵ
�R
�M�9��z(���z�O���w��]��s�CAl��$=�X��oXn��#-��d�|��ќ�� �/�X�J�y��kt���ۤ}!�G��
f��m\��-Q>V?�-<�K�U��|�U,�����-&z�jO&Lw�Yja��<�ە�0�wR
�����_Z�o�[��g��?Hc�wsG�8d�Z�:����Ĳ���6����ۿ�w�rd�c����$�ǹ���[�������]�Jl����|��k����h�� �n�����Y����.@-E~']i�J9�sWs�-����e@��jR� �P�;Te���'Rn��(��X�{2��^P���OO�C�ӏ1V�1F�8(gf�w�v��o��Xyj�k2ny��p����,��w~I�i�ܛ����A��G�ރ�G�q3᲋��н��"l�W��8���� �C���T��Z��u+�:��I}���HF���Q�� �9�>� =1�*�l*ႥRG�6�{���4����>���#�e���|8r�a�H�$�}h�I�Nc���&��U��8=r(��+�/s}�����E̿���Lȭf�n1�<
���F&���Ӆ���^.���3��6t���	��øL{��k�\��3X�Eҿ��v+9��I���;���<S��ק����,��[���v�����]����D����] �H��~_��(	�7^p�Z(l�΀F1�o&r[��;O/7�u`��!dţ��h*榟 Jf.��7�;ap����Jko�
���4[1Ҧ��\,վo�f3K9��p^��1�Aͪ���z���k���.�t����[:lS$�t|���&�����&6�K΍��JG�a-"iD=��j��N._y�����r:�ՎX)UKL��-@O��n����;�iaԬT��������i0<�aI9"v�r �Y��X��^�:�l�i�p��㯢v��8\�0�椵�q�|�Tb�Y��1�*m�ı��ۯߒ\�q>��-~ԝF�>`(y��J�O��p��lL�O��ɿ[IbN;�"�^����$�x���Ş~<�# �2�0�rzm-� � ���Χ01��AK�,�8}0<���&q���g�X��qs[��g6;L�0h߃R�X�/�t �0X�����1�C�)���6�}�֢n^�����+!�[;8b��4r�d���n�`]M��f�aE���F؈o�w���L�n랐����*���H[��WE?A��[����e�9�Z����v�%ʹ{*A<���5��Z��w�7?L/h��sߞa�}Ȏ����k@�T�e����$;�p�ړK)M����,@0�*X���-�m����5��,�DWI�;���QX���[��F�;�oә�I\��02��X��*�n}���Y]�K�}�÷wu���� ����-b\p�<����&/ǅc_D-���?�N�֠Z��i�	O~��G��%�`t��0�j�Tj��
������O�>m�2Q���
��Q* ��w6�:,OA�8����	��� ��.��b6�ď�a��<�/p��La�Lw6��c1�x�g/d����+��?�?<���Z{�0zЮ\d�7)a�@�)�,��7�i�������N�Z�Qze.WH@;X��{�^�s)g�]��F�'x����1�O�� ��ma��4��<�Y�+@%/ .1��4y/J:0������%���;���Iv�Ò1)���r$��nH�N^xP.��zߴ)?/T�Ő��Ӡ�ތ�r�G�D�G�+lD�Ҽ>8G�B��coSq�/�(oF+���>޾WQ�,X7������/�Y1M����*V)�V5��[�p����Y��Vs�N3&�9ή�r́7���aV|�Ӎ
��.>��d���\��L��7f��|j��e!7�Gg8���S=�7�E��c�4�$U&Mz:&��V{-�JD�C�Ԅ�ꙅ�m��3��0n����ʅ�~��F#gX�%q�q����7��x�;����m��"���TQ��t�k�Cǽ�����|�xR]��υ�����m�R�����;�=��?`�p�y��ʹ���~C-!���K�w;�Uȵٯ����F��t"�K> b��q�o�T�wqL��A\1A\=�mY͚�+n�����4"O�W����,A��u?~���\8 �[W�2θ�%�V�h^$S-�i*��� .�.��X��A�q��*��k�� S5e�RT��lGi���{J��V�)+�o�
+����wnJ�ӶvJ�3;�]�ĩ����t&lz���&M�]�"8��Q��a	��f�ݮ+ʹgy?��|�&Jn�u����P�A�z��� ��j�M�G�Q�R,��dvIZR7��:N�����.�"L�� �6�7�1�" h��x���V�����Ɣ�c�ڑz��Mx��)?7�]$�EȮto��n��:���36��5�c����$�{E�=��we���JPGo� �0XhGQQs�n�Y�D��(k �r��CG��5��ҥ��vj�,��蘜ʥ+Sڕcn�9&���0}28���A�f�^�uZ������?q�8
t���y��`��<�&�qd���m���Tr���
��>�����s[�XzڜO1�Hn��X��)Ȟ~#�����}��7���@����v�E9T��M�V��g���'u�f����y�h��I��m�����N,Z�ڶ$Gmm�z�a���-��J�M�{��t_f���[\#P�o�lʦUt��\��`e�9�7xT��<������� [�q&T�|f�OT�=9Az����6[��	O{�۴���J\,%�cÕ��J�lE�K���q�S�[-�Na���z�2���L�-��\�����k��Q�Զ?������cs�ӳ��o����pg?��L�mP>�@-��jQ��SyK�����wb�`b<�c[�u���EHĎ����)0���
�j��~18�j'�/
��6P���|-�{��iF� }Un��>W��f���<xkIY)�ҫ���������.���uYm�F_��ܱ�Uf�GePn���㫐���8�aO�>�'��lʓ6}���D����0'��� ��Vw�K��-,��ZW���*+Ɗ�� !x�]��H�3`�y�S>
��tt�[��ť���;dZ� �3ʡ	�u��8�T�v�V�]�zv�N�X���}�a���P�#��Gtق���Ԏ�j�b2��^�0La�5�R��'^↧ձ�zѠ��ΐ��G��u&�|n�=�l=ݐ8��=�z���}'�׺�U��$�<{:S�T�9zD-^�U)�t�7z��B�b6Q�������U�U=��ۺ_H�Z�Ej <6�r��g�,������E~��\���)�����T�pM��.~"�Ɗ�0~С�d}M],��Й������Y�{n��]���5NAvs�ɿ�w{W��]*������m�Ax���_�V�;� @+��`��EE^<U@*P���ȍU��?���?R� �"'�}�׿Xw
����1�x}ߪ¥�M����eF9�|��E�����9�bX�Bl�[#���0eA�Q���]�|J����*����ǱgVIxO�Ϳgw���הs|��������w	�->����ӵ�NM|���q�������?2������{`ĳ����S�g�<���ˡ�#��f�A�u��Z����Suv�[UH���2�zk$R��M_��m���+�W�{��Pc{nΎ��V�:u��B(��' Pe�Nw�swh�,���hD�ip��(�h����`�hҬ�;�iӠg	���7�;���I���}���S�����oKD�Is����S'T�ێc"a0����8eN�gݐ`��xp�4��6�j���Ia"ׄ�B��� e�0�/W#��%��SA���Ix/�n�ì�pеZZX�o�!z]��KZ[�;���=I�g���(`�<>U���z8*�ь��^p%�dR�ɗyP*F��T��,U*���[*�8���=���i�Jzk�0tG�nW�l��d �W2Zڣ�F�&�b�psa5`ޜ��������J�4�_P`�EB=���_��D�Z~�6��:~��{r��X�+e^xHE����-F���n�δ����K��R�.�Ln���3�xE����{����S��IO�T���f8Զtu�7L�3=�|�d�a��QKߏD�d�w���w�:�do5 *�oz�'KH\�|��*Q+8��۴�$��*�ɠW-T�۠�%ʦ�.��X����X:I�}�;������
��0���+��&`�EQc���|�R�:x7��8��l�ڎV���)ULd�/����� Ytc��C�R��x���X�Q�g�	�~��M\9�>�nr�����}����vm69c�CU:<Uy��?�ԝ+ڽ$����&�@�����'3��.%�W�XECf��w����w�?�ܲW�?K��;ĊH�����f� �xe�u����b\y��U����.Kf�ծ�7-.3۰LA�l����뒺NcE��2���?��SM���/����$�\f�l�igz��$O.kg�s�huy[�Nv���_3������[;�s{���)����m�Ί~��W%����#��9�L��W6�4��r��"9�!�P�F�H��_ZP���I`�l?:ʿ|�\~�B36T7OK�u��!���0���O/F��f�^�)��Lc�����R_�v��`�4ViLy� 0+�JZ�z-h���m�~:E�g]�L�ac�רI?2��L;a����GM}��}O�	 ɳb�V��_&�ɤ���(J\[��U_�"¬��}���B���If�I��ӫn��d+4_�Mo]��ږ��.�1�-HfTSeS�}g�H�$�C��v�t>����g"K>�9#�C����V��1��A��y���=b_z~��ߑ��θc͉�'R�{M�s�L���`�*��f���=?N���M7=��
DQe-�T�.5l��80a��y�oC�IU!dzr|�&J�b* ��}_�'�P��x~1� �{���PENC�Վ+V�t:O�] �`~o���x��{��}.a��?;���45���z��E��q��s7i��^�ni�x�&��ѧ5ނ<5�;��� >��Nf�i��e�X�F�G�*�oҥI(P	�,P�3	d&��8`�|U���)��,ػ�ܓ�d����);�����~���� :��Pj�ɏ�7�G�Z�ݔT�.�Ld$��Y�ջ�$7��rR�� HhAW�4�n!c��-� ��Z��j�k�f��X���� �R�=���`ք�b�Y�г⫙.Ԙ $[mkn�r�Zचn��ЭT���w���k�:��[~���by�zyLQæ-�Gۙ7R��R������i��}n�����
p���+�0��]��6i�@>ʲ&3e�PR�j�c��,�1�x $ڒ�鑓x�n����i��HPV�e��/T�Ȗ���19�q=�����0�˽}����nS�+}1L����긽�_���f�8��'��Z4�V��$�W���s|p2Bմ�=�:��/9��'D-z�r���)avi�����$���W@���=w`�NY!E�����������X�����QFk��+��T|ȼ�=�в�:����3���`OR���Jcdp��]S��6/����<n�暔m�I_���Y��r��Ħ�N������J#�����@�`����L�/N��7⫤uڷO�~�]��b-�Q�(	��VIFU�����vx������l'��;�- ����R�,*�c�C�4��G��ý9�w��@{�HDƪ��s���E/�	XdG69�"��]N3\�^
���K���$����+�b�Ɂ.��d���aD-��X�c�볭� ���_H?�#��8h�����i���x�~���?%9Y�E
K��V�T�2RO|zX)'�g�ʶ�M<���˭�+�/� nb��D"prat�H��ȊX头vHGA�q%��}�HFk�5ҿ��~��~
�<�ӂ!0<��r���E�5�-���:$�7�f�&���%����L>�SZ��s6^� �ma�`�
�Ӫ�u�\rN�����1�B.�XQU�Mt��� ��/���<�F#5�-MH��gO��L�Ay��I��y?�>���s
u�H��̛��r��Ƨa{��Ph��o��k�k:'�kt��E�U��&�;�o�.���:vz�Pϲ���&��Ӹ�$͛*7�_��G���j*���Ro�`q����Bj��+C;c�s��>,2[��k��i�DbrH�V���5Yٺ;�u.�����#4��l2=:��Tۨ�v�W�}v�R~a������JÐ$�	�"��62�{tW�G6���:�s)}?����᱄q�r�����{>�Λ�-�[��T���2�p;�<q��Z�-t.]Q{p��L�
�nc�}0��.�m��gݤ���5�E=/}N��,�Ή��<s��ʳ�0�kk2���T4��;S��]=����*^�+Y`���X$$�������@v��E�9[&�u9�m�azr����@,��gI��;o�`Hi̓�����/��#zJp�*�y����¹ �k(�f��S��g;�c�pi�^���˓[;˓-��A�-
7n|�Ș\o�E�k��ܹ;��i$�M��QmPg����A�C���;4Tz���!AW8��Y�w콵�C'�z����s��ƻ�2���[)���N���T;ԅ+u*�ӣl���.�����zh�76l:�Ү���612�ǐ_3CG�drcE�1���ID�M� ;��ݹ�s���-���BיmMcDN=^����Qu$-��:�_Yp�<=g�  ����$_�����R��_2\�;����_�vQ�L�t�ک=�"(]I���5�v�'2�갮���全��z�̧g��4qu:t[�c]��n�ݷ�qp)����eB�i���$�9�O������s���	�B��3+�7���&F�{JP�K��1#�gF�Sid��"��QUB����@\n�쟗JZ�Py2�Ȏ��A )�1�p�v}��(��bf2�Tb�tb�@�ܕ����:o�����r��'mD@�1��Ԗ+t��ľZ�pW
��C�H��|�+�:c�K�\ua�J'�"g���7���i�j��-7T��u}j��u���3���p@�?��Z�7��Y��,���Q�P�~�����1݅fM�������8�����Ș �f�<m���Y��	ƃ��^��=P�^��-�r�fB�����x�'ʾU��͞�^�ؾY���?��G���g*NpF����hRx��R�y��*mh�@0�vЃ�(+ۑ��"!���5�s��ء�`9�)�@P�����[���җ��u���N����J�Z�CB��MA�S�d���&�r�lGs��n'�"j?�Ĝ�&���@`�V�����8c�b��w�P��vk��#�K��F۰���U�7f�H8�'��65P���#��f3��J����oKj����9�Wd'��`�d��W42�N9��!��֊g���A�kF��	v��V�I��ŠF���t�HM�mΓÇ����xbz����������|!���	0���_�u��\�H�]���"F��n%���� ����I�B��h�]Pi<���b�q�^Y�@ v�G���\���n��}9��&L���6B���*�,o���'	�6,����Z��)�P�x�"���U�Z��y� 2hىY���6[�Z�Zn���"��߷���t��wf{F/�űDz[[;�O��+���(T12�u�����1���zYe+�nO3�51��X�9<�W�G�ΤN\��AgM7G��a �N��0�v�����a~�|c�Z�����P�������WZ�! ���|��IX�̖��9��( ."�x�V�L�VXR�`� mNF�K���9��$�,���_֭�v�	 j�%|K�A�P#G�8�x����%ց
{�
A��ê���Cz)��u��=��^�ٌ�V���k�=la4��T��n得ӏ(k���w
V~[�ژ�{G w'�E�=n�@v�mL�PohB��ۿ�êұf���� _��k�Ĺ9zr�$�K�+�O|�[S0�l��c� �@NBm�&�a�;���LT"�ȓ�!F����l�d�V�>�o�::=����L��=�
'�+8<CU���֩(�h�3��V�h�ځ�2_z��>�6G��X����?J��˃�d�������K�Qn�7���bn�S��bNp�T�+��#)���S�j��lk7�5��H�����5�)Eu8��<��]?0A�W$�:�8`H���i��hP5P}m��O�|�0dn�9��}')�=���{��Tü�����U�ǣ�a�,��]��
�!���5��yJ@��w��,Fd�#���.���Ơ��=Q��2�lfU)��s\��%I��سM�rE�.��l���U�����a$-��SBa�a�c�y���Q}q&2�w�z툺l�FV��`���8y����I���5W�k^���j��.)� 6J�`�H
�[����K���o����A��%��L��B*��$<Tx��� ���n�?�B{����I���C,6����x)����������$-�Ǐr/)��<$ 2n��	��{.�9�ЯG��i�*�j�c��R���uP����3ۺ��v�[$��#moR@��=X�t�ΦY~;�b�N$������=L��|{l#j�榮l}���1mՍ�mҤq׾��������<���_�Ļ.���S�Ba`�g��&L������ �ރ����r�!��d�3�	3���\~��q��G���S�j�H�r���NE]��w��r[+m;�a2_f
���
�$/�� �XCv3��<%hnd"A����ou�������#0E���70`�8G쵍�K�� �>4��0�@{(n9�z��T�ɾa�s��ѫ�8z��n�)M���]�T"��ٳ��+<ܠ��z%�9Η�캴��2��E���x �%�6�R�(pv8/A}�x��`����$Xg6h�:�?�}`4|e�Q[f�bDk>}�Mo�_5&�ֆu��4�T�A��.�P*�5�����I���
���<��7���D��ŝ�?����"CS�.�ʻ0�IKS9�����*���;�ּ��o��d�`���;-�����l��G���;i��}�ژ���{m�B@l%yt!'=���e{��V9��qzua��@
zt����oq(��+<_���������T�v��R���<��W�2�ؘ
�N�窸jE��6���F�信Z�
9�I��~s��Q�ٗ	���IRX��83c�?�b-�@a&&�YG�u�η��𺲟� �`,�Ȏ�k�uW8k��6ݯ�.� �uk�R9`ђ����ڻ �����%+#��J"^(�sa��<I�7F���(�Z�QP�SG��B�b�$���@~oZ�A`gal���!_VNp��t��)W������o��Bn�GG�'�sn��GS6?���u�=l]�J�� �J�o#v�H���>c,X�<#~V���M�M�G4��}��x��vX�h4Y2�̓�'A8���/+�J�4� uH�vYlj�A�P�Y�� �G��7ޏ��z���,��z��U�a?И�!�@t��8�[ v����^�N��5Ώ���Z-�U�:K����J]6��he�<౵ n�+�����H:x"�tga�W�P�ǉ=/��4jr��L�g� �����G���rq����z��Dk�C���X$H�3sU??s#~�YJ�
��>Z�
5�@@C'�i���jЍ#�g7Hg�DC�B��������5<}@U������G���T�+��[�`�釡�<4�z"*�
KE�ꣃn;�Nڅ�	��ۦ�v�/$�М_i��ܱ�t�5�[��~ .�&�}KL��J����QS���k"��[�Z�,ir������1� �C_����r��(dD�^�="rI-�Ж�	z�G9A�����s�{��|��/|�q<m�ÈH�ro��Ļ�v�?ԃ�4@�I)��N̒�� r r�t	7�+O��6u�����U
aw�$��/2)��W+�$�[��':@
��6S��/�8ʿ/�x��Ay���~����R#h|�Y���<���o"qs۱��8��[������QtLQ5�^AG�	rI���'/�m�M��,������ɍ�`�߿���U����Z��s��:�Ս��Й���Td	�{fax�%@"A�zi'd�����,\�X]�~�&�JE�����p;�!��.������=d��0�_~^�?��Q h
�ِ�tL\ή
��⿫"dLM��7~:=�U�K�c���q��bw��>�XZ(�L#����HP#N�OJ~zr0���❓��wz:�������\L6��	�����JណP����CDN�s��1��Brf���<C��\nW�/�阼��Uw�q�x��C�1B��͐�F��W�]3��*��2L����=�����H�������g��an)���C�ǖ�,������}9�7��)ή�o���*�ӟ��c�>��p��Di8��ǵr�vw}%��i��R��9�b�X=���y�F�O�n"�+��u�)r|�"f��g�}�*T9�1)�:U�o ,�+�[�҄Z��.��R$�(����	X�N�h���.s�b�_hw7�����`��������zKߣBKb2oX�a�/���V�x��7	�,��=��l*b�=�����M��*�=��w�ީt$A�ڤ9����Fz|�l<��)�9��'�dݪɝ���vC{ZL?vv��C�/U����>���q�Q|_������Ur��tNCH/ �g7}߰7��RlT_��m��;^
,�C�^�Z��!1�I�|CXqb[�Y/�Z�S\,4�w��c��ab��.�;�PT厲5�9Gh��l
���4|�@�=�N;{<&.,a�ʈR��ux�O�]:�Ë�k�n��l����*S�!-�boT~�?�c�%����!z�[By�������p%w���lDBL|���}�_�z(\0\&�?X����N'tɼ�Tը���t��I˜�e�+d��I�+�$�}�Wã*�i��̪�C�89��Qh�7L7I�wK���M��5�կ_�5��n2�b��G�l��LVq��D�����w�.�^a�/&��y: ����25�m�����[��T_�n\�$�]�#a}��ݟ�b�U��V]f�"L2��
��x�lJ����H�[��pW�dٜwg�ϗ���> B�UQ����I+��ᤱwl ��+-`ߠ/���k�:%?��C0%=N�q<!V�dR�$48���%h`�`�Y�TE�{x��~��vT\��r�#�>��{:�b�]�`?�b��e�<�Pxk��h����t�N@���[3���6h�;�[���v��}迸�ז��0��]�{z�{�X�+��J�@����;QvFA,�Ż�����{:��+��7�F�y�.Bs9��S`e�ua�a����O���6T�q�c'C��J�Tg�thw�t��{��e+ ���C�'�(E^�K�7ذ�-�^���,h6���6Q��;��=���2��1�h�Y��Ro�s۠u������� :r>�[]hu�S$8[�ó�d���l�Ly��R��l�0���Wh]��_��U��hk!��2o��/=1n#�xTm��5�#�{�%K�>��s,	������g�v�6` ��i��=a�'����_W4¸b��`^���yR�U�+c���Z�5m^��G�N�r�2�m��Q���!J���#f�E�a�ʟ7�}A���|N4d-X��:�,�>�ᦗ���}�����PSջ��t����S#�a���k_����r*<��WeCVŋX�?�������'vђȰ��5[�F�
;�)+;���k�Ձ?�܀j$a�g��4�F�������W�D��lut�!x'!����΅��\�X"q�,��w��(��|��x ~L��6��tJ O�VV�;L�r����3�mh��:��e;~K�@��Y���϶@f_j�vـ�0 �ؗ�O��^!���Մ��ݍ��f')n*P��í�k�@��T��h��W�zT ７t#��3�e	>��2E�a�C�mE�=�$y�-�q$<E#�^��f��gs���}�]��}��4�x���6�^dr��5ʀa�����*�捲�<��%��zv3Fx�@����1�c�z�@�h�Óo=$:��|��'(�Y�pvE|ޚ<���@Ӌ�:׃0n`��t�Sv�e�p���f�;&z������g�� �q���e+�G�Mڃ����DV6ʵ����L���!i/2�o�%f���Ϗ�F��߶!W��ƚ���/ (�|ANg:�O�L٬��p��,�M�`��M�IJ��E�0�V�h�SU� ԁ���� c(�D��ܞ�ݬ��$�k��q��SD[xlc0����L��eNo����K?o����q�EpY�V(���B�w*��V
�+����32��������bDo���Y����2�~�0W�GG��|��[�X�D�H��a���5��29�a����wڑ<&�+q��w;e��Sk�ڪFq̔���1<p����7!�3������<�Jp�%:�aa�O z�I��|B;ӡ�"a�p�И�_WY��=�zE���*���&C1��4�$k�/pY@��Z
��A�&N��ߞC��c`����`�~�`�����:��$� e�X��fAF���L ��X�P3;�w	���)h�֙;�T�(�W����B��1��f�7�Q����q��cׇ{V���fw .#�Ӭ�}��{y�� ёb��oа>��k8/��?�2��C��S
Ԏ!P$a5No%x��� ���2�����]���a����}�g��&[��<1���T&��A榀�8@���< ׶B����T���T�;�ʬo̅� ǈ� �G���}ƈ,*�=�1��#!z+,��#�g L@��A��)�VK!K��upԀ0F\�Ԋ�Iss�e�Dt��)PrVbთH%ۘ
R���d}�U�"[���I*H��<�`$cp�B0�	�)"D��� T���yTy�q�-��C���@�,�=b[�22�� [xf0�>�H����zl�8�Cs� v�oa���H����T�3�mt#�>)pSFd�3_�\ȃb���
t�����v�;޵괇!Ç�0:�(%�Q.^遞RFP�q������A'\�#������Վ�^ʨ��)�B�`��@���s��p����GtT�|�2#�O�}�e� �nd�����q.�iY�|m�mG�yLr�+elʥ��{V��Ն`���D.������z�Բ2-w��6^qw_�;�p�,����P�[z��h����K�%��`J���"��O)�Iz�������R%R��2#�lX����̥6���#�҇w��9\���� DZ����>!$�W�E&ʚ���p?���D�$�-��d���Y��T�1�|$�s���9�fgw��Os�#`@, ŋ�(pg6��{� �w}#o��{���Cc�)v*�#�;�2����K� ?N�F�N>�A�@ĐmZ��v�A/�"�_�[F.\D0�w�
�����Ƞe�AR���i+d�$��E<�_G�VC��%2Z���'�#"(�/�A�TQ��a`{�WMe��3N$��<��xnu
a��<9Ϣ���7��è�O��t*�^65E�4Zt#�O�^J$�>�q��2�+�r�y�:�R6-�v�Jl�&�$=��P�p�6���:`���`Dǎ0X��<��sJ�<	�O��<j�xp!Ɛ~L�Ht0"婉��aHW?��C��F�fA5��c����Ӏ�"%�y�8��@�/�!u�?��� 3�D�ߙ^S�E%Y�"E0!�,�� 2i O�
�:�Ƞ�� � 0�1�w(�&h��I��
���,2jUh�beK��/aK���
����zȕH�E7cX�����ϣ���X.d�� ���e���$W����FC��A�t�&�g�)Md��5@�&!K�����Xߔ�T�E.� �H'��ü�5HW�̝o�c{:�?�C�2@v'@!�Z���� �^{��	\]{ �h9�pDf�Q_؜b��R��O"<3oDLt2�����e�bd��dov�P$��ԁ����
��G�0�L-PQ��7<^z23��GƇ�`zW�HV�FrM�))aRHN�1B"�@�L��'�¨��D��wg�b��b|�j��b��W6�Ď!����ǟ�D�����ީ?����ֳ�S�@��3��'4�O���1�3����8����02���hw�q!��t��6���FqO����!y59�O���C�i���*��+��`�ίclf�x��t.�Mf��L4�S�_Nx�B��y,�ױ+ٶ$
�y����`W���H�[ (���ETᆅ�}
b��
mbv�f4��."�;���<��h!�8z��ifu
8�n�ȃ)���XkSIi�Q|p��L��R~�;n��#Ѩu��O��dq���ϱ�@Z�zy�I���Q<�N�P�E'�'� �r��/���x���W=�$������2/��`l�!�l3G&Q�͓���FiI	<�G%�G����"�򝄺"���IR��ӳ!�l�7j�p�#�bѝ�U6�N+܅�mM i԰�&�CL����r�J{��e3d+H�g�ȼ0�PREg�M���ID���㲩���C�Ɲ=GH�y��hO1��(�H:H�p�Q�!6Ѓ�(m/���'G8R��}��jB:�G8��z�X�~{�9����ז>C�P�/^0LĶR<���O/HSFv~�R�"��0XF�"@�~ G�ڞA�0��!��a�H@
���}��b9f�y�Gˡ��m�F5��]��^]�7y����ެ�Ԝa��}�h1�ǟR�Ď�l����z٦�b(N��-\�Hu}\&�I
.�?�8�z��t3���El�&Eu��]��%�h�&wm��@i9@ʆ�܋׾��U�x�)|���F�ҳ����V
�h��c%~t���ZW>N�������%�Y���ޣ�p����#Y[D�F���8
�<�̀��|�p��S\�zD��9��b8J��\^1�u�r`���.D%ĠN,�Ĉ��f�r5�<&c���և�ӥ���A�_G�tH�Bfj���̊uM����@���[��ԇ�6B�����2m�A��x��������2��sn�7�����x6E0a�oC ���5��������� �P�z)A�Hہ_Du#ܞ�˗��p/����S�_�l�e
/\��r��/;�?�6RP�D�w�@\�w?��[(f. ��2/KƄ&�_�8��"Ѝ�����'�s�CL/8F�������˰����E����CA����F@��{�4�'eޒ�x	Wr���*� I��⿪#vAv4J"��Ơb�lC܉��b�/Bc���B���O���W�������-['Y�]&R
��
�����o���w�_H��92�����&������A:x"����v:�����߹S������s�%��ضn���~嵭�m�������_���)��'��=B���1�O� զ�Ñ(I/��7{��Um]�I����d�P�9��Mǯ�<��u
9����6��L���ŗ��{7. ����Ȯ-���W��"����RH�?�co+�����m��!�[КqH!���#�:?���0S�=���+��o��>n�P�C����<1������ȡX��T�j�n=YI���U�ւ�A�p\���lk���� ��}�OH�C�,��^�r�_�FJ�ԅI�kܼ�AJ��}��^���L	���ܷ����k�%�g���L�Y�Ŋ_�����ʓ�7�)u��V������� �v�z�_�$�u�����B����x�s�/m���wJi8���=^��U��ϠV,��k���h��w]q�4�?���T���S"�����үo������������"MQ���)x��M�Y�;�^��}�R����C�z��eR����w�4���ڈ���w�wS�����&�����I�m���X�'`{tD�^8�#��ν�N��ǴH�dE�c��eZ��"B�|[���:�h+܂�)v�~������f�4�Mx��"E��%�4���/����k�P�t���u��8$�o�;f�_Z�pu�)��o��|jqu���q�
ʚYfF�<��_'��I�B��R��֧��^���@x�rho����8�8Ga�"�!��)@�]���a�!i���̐KR��1���:��J��G�0;"��6m�eD"��D
��;\�Xpx߾�ࡨ�u�.A�� 2��!�#�]�l0C�n0V�ƺ6V��6�C6��g��&D�ҽ�)�FCNL]��r�=�P*����;$���x����k��%W�}����I���tAl 2����C,��������"��7�{'?]X&�/����D-�� g���m�q��@��R���S���LpQ!$U|��/�����9��-�He�ݲ1yna	D�h'���	��CzO��)r��A����em�(���^�(�Z��6���I��������R��֛얹K�fϥ6�<��SlY�16\�ȥ�%rn���)�I��H�O	�3-�w��*�gu���qNȭ�H��s��!�s��2	Dl}����A�g�[�>)�����o<I#c��2�	cF|y^��6����һ+��_@���ڸqmR� �`�7-�����F�ޙC�: �
F+���+r�cz����ȥ��C3����ja�Q_t�F5A�Zx�7�d��ȅ���c��Z�>R�e9������a1��y����h�g$-LP�ᵱ*�9��}�I�g����wN��.��r8��ys�	���>�m�A�j��Sֈ�Yz}P�Pb=�-�Sp+!�%^Y:�/�)�y�)� ����|a������o�ژ��z�5?�^f�n'�e����WNz�T�޹�#�;_���ij�kn��*}����L�|�V���a;��if�ɥ�v�Q�1�}t�q!f�0n�NGbW����'�:4
~�S�q��L����σ��_>4�D}���w[->�yg�l���l����!�m�� ,]��7,�rg�7U�����˘U)*���<�����4h�&�p;�Q��u;��"�Q�R��y�e�
)��1+2sT��s8f�y�s��?�o��k������^k��z����c�'����
�wz��	q^��{��q��;��yJ~aX�U�G������,	�{q�8�_�>�	mZ���N�C�A�/Ad<��>�8��{Ӝ'q���9+M�ˏ��
�-h:d�`�;�x���:��o;�鐵Û-��W��rMe�r�Pw�Gb����(M������8�A}�M�DԴ9�\��>qZ�VCU:�}/@�e�F3��%�=$�N�A�9��/��t�Ɓ��]�§�4(T������ç�ⴔ@��l���O�i��2���.���!|��%R�HӋ�������1ȋ�GhBѡ�CX�̑�{�S����|0���g��P����8��NQ�>�4&F}t����skP~v���G�t�5MT8^���Ȕ�-w��-0��&L�C+]U����i%_�4geW
��ۅ\����g�;��iAO�=����Fsֿg���iV�Zx
����D1�&��a�h�02U����� .����<c�g낝�v�<�ѸD��&ؤj��S;w�i�xL�7K41����.t+4(S��4����ؗO1ؿ��:�k��v���t��ͪ3�
^s���*��2�����+=�[1��㦹�f�}��?ǜളi�zKsaq��{��h�L�~R�����f��?�QťYK^�!���2��%��� 5�+��PNq4]~���m�f�=���98��&l=N{��Mo��^/�\���t�?����rp�w_�~hv^O3
u^"���siZ'����:m7�:S;4c*��a{��R,�hϚ�ي�J���/WU��h��(�@���K�D,�gK@�~ie��xa��$��w��6�(e�dR�[��(�ʕu�ݹ�F�I�~C�UP�&F��ߜ������9��)�M~�t�s�*����7����=��m�di���ĠS�,��QIM��%����C�^<��e��0�A��L��=�g�iX����S�u7Bl�>p��SH�և⑖��+
s����]�C�pq.����4Ƃü�1��.\H!�l�'�n&��F���(Bz���
�P�,����s)ؐuK�= �U�\��+b��J�����n�y/y8��1��q,��P�S�s��qG��<�'��w���v<!��d���:��c�x���4X�b�^?H��A��Zͷ�����	d�1ږ�֎ �so�*�P~�x���-���Egn�FB�@�B�{���GHĹ���%����Eo?r��t�5��1��-1p�3���F��������wM3јJ�Lu�15%��� ��V�,.}�%�?������W"Zok`����i;)��\]w2�C_��o� ���9�ͽe1�ȖP�s���'1�����wiSϷls��:p�y��ۂtׄ���l!��&3�?w@#�,#��Y�^���-����g8ҧVyh/�3P�yX�e����pO3�捜'�l��O��5KV9��綜˽�Z �������g���Ik�b�[�yp�|���,�DD ݺ&�iM�cc+���6�����ǜ9����w���|���G�g�>c|��ƀ��q{���E߸%�����!��~�rۛ! 5��\���ga^}�+�~�%���>����;�M-�>���zB���έ�bP��a�q
�?:v�� �u��e'��כj%��.݊z�|�X���F���)ߩ�F���p�9�Jl�����u�n�[sP��Gcx%P�B��߄T[�fߌ���(GGg�	.}����xZ�kN����N��� ��)q����}M��KR�ֽ~�m�x���P���N�����`Й�
�q���$�$�� 'TP�p�TH
1;��՛���Pq���N���=�3n��;�kWX�4�yd{}B�.�渼�����n��U|��	�I���|j���k�N�2�ٚ�濃��7�/O��s"?v�]�S��sy�}֠.�ks������!�u�����1�g@�O�����a?�	d|�:T�D1�*����bEX�����j�zR��̹?y�3�Ƌ11@d� fU�"���PU��om]����B
�5�D��~VV��R�s?���e�;F��}�W;�6S���5Ww�g�a7�F��w�Au�oM�� 4�|m�d���@KG+wb�H������AqDU���x��U������nD"�k�َ�"��'��R�q!4�����:\*�ċx�2@�4,M�	���P�hkt�ƪo ��濧ؘ��%|֐U�#�L�r7S��I)Ԅ ����u�_��C�����
�D����3m$��J�e�B0��	{�f9֫�&3�lãuGO�P�w�i�T`�:<oNW���Gߑ�=�����䒎��@y��'ص2v�C�e��E.l�כ����a�ޑ1�29�5��q8?�9�{��{Y���v��9�:�����t��� d�$���z�sV�����L8#GO�!	��vjǿ�?���џcԈ5mޅt߅��Էy��� �U2�^|�g�֎�|l�_��w����:x3�0�ۼ��Ѐ��xY�
M ��(0����{l���U���H���T�L+�lmH��Oj]q�+��KP7c�7��
Π��m�K)�pquP�A��z�nb�^������L:���֬��b]k�B�/�f>��aw?>����̧w��Fք`�Т���j�Q���/O�:��"�5�*l=���g�S�*���cPó�w�k���BV6el�b
� '�,>8�n%���D� ���@XɃpܝ�E�#=��<���#pS�2��2(��N�y��Nc?�W5��z=�x���3�A)���]��
�� q}��������XY\��J��ZY��s�~抓s9\�0*�3�G�F�m�b��%��\�vȡV榱_}\'�]��:�B�ϣ�YI��QT�k&�FP�dj�~��u+{������-M�q S/�2˪���Ķθg]��n�0��o�0�}��7��4�m�k��^��f��*{j�8���P�_�Ӊ��[P28�������r����^��l��M��q��zQ�����bn��19���@���7H��J�i��7��=0�ej AO�~,��	Z�p��/�ȗ���,VW������e��m������-0gG�_@T��߂�oh�U��M�c��
�yBAD
����%�m�_hN9 �	�����Vr���"�� ���B�_��x׾���� �@r���O騷/˛)�k���s�.�f^��*�h�5��!�Й��q��S[Bs�x�u��AUE]�����������0Qsg���be;��מ)9#��s'�:�9n;3!}:���cZ3/�7��v����l^շ'%��k>�\p� ���v���R���_ē�',���} p�Lq�gb�[���!f�G�l�f���	nN���u���G��R����-%�s�����,����%@��%C��C��x6~�Aq&#����)搠CG�i���6B��,�g�	>%6@�	(=���n�ԅ@o|���j�`�7r�κ��c�q��?}�~+Cu|�CN<
��.ݻ�8+<F��6��\����|	gSL~���UR��arR.4٥w)}�-C'��z'<h�CW�ATS�0|���'C�G�{��=��=V,9�d���'P@���������2t�Fq��\���x2��)!&��ƍY�#"��}/��-��,s/ʅ�?x��ѩ���x�μ-Lt��:e�\tτ������2�&v������W0~ 7hg׉qVT=~�%�'�.�s��Xj����P�Pߞx�!	s���-����;c�����ڛ��L���^�-*V8��V�š��!�����(C�^!J�N5�Z���	�p�o��>���-�Aw�h���y���4��;6��5�-���H'� A%ϧw�Oɡާm��k�|��˾�W����	�2�	-�&3�^Rh��g����D�Y��lODA�"�~3S}{T��c*B0��نl�|�Z��;E�T��wlNx$-;�p�)T�"����U8
a�#��Qi'���d�q����$!���
�*��m�B��Fі@�\�\T��U��wd+w����<
HzڛD�h# 諜J���(��>t��*�MW4D�agbM{�6QAX����B}-3�|Њ��)�;�J�8 �bu���̕�US�m���+��âa︉�C?C>¤�)�Lg�NXXY�SK��7X*Da�+�.~�n���O�1񉾣�u]m��Vݯ;n.R6��u�w �_�bE�����:�Q~��sk���{D�Njш���R2��s K��Oi+���mG�y�9���A�a\/0S��Pk�����O_1��;	.@��W��) ^�����{���"2;*}���� ��a�둩]�ߝv��s]����.�o+D8�ތ9E��V)^�nѧ��18�u_s��W�Nޞ<�V��Q��D��a��UC�:r��m
d�=���%Y=���	̡�5e(0���?A�E_{�XphvPmW�KP�G?oݢFE�?�3P��������6i�cLw�Oж�A-��w�*�����
ߞ`�5�*�Բp�0��#1��(�p4e�݈Pwn�*��3����X`�d��w��0���4�=�-����
��k$VVoβ�>�����db]�y����2�o}[a�/�j��&�y��`�����,��]Ti��I�ɀ�Ѱ���In�����4�B��ỷ��������(��uB��%����9��-�V=��LB5*���M���<G��A�����55���rQ�ZyY�,	E��#t�%%Ie�d�.�i�'=K���!�'2�i?1xW�2׵�ݰ�����EV���)s1�v����ܩ��Z��Q������u�G��}�̽Ry�%+c�y�[N9x瓍�^�����K|�D�|�He�G�'�.��_ս�AG�EP��7=e)�2W��g��݄���L{]���[�2y�<�`'�E�Dh�����*��o�h��
	�SP����p���M�+�N������b��d��[�	|�E+&;꿧���9�����_Hg���	��W�x��DM�Ʊ_k�^�T/�p[�{��8rkkv� p���z�*��܌�٩�in��M�2�Ќ�=���N�	�O�K��5ςŕ��[Ύ��[�~wA��F�W�
H����A� 0��ɮ�N�R������©�l�2

��__�"���E�'�9��*���@�	0��C�A�pչ�>s�I�#�����zC�)�:JE�&^�L��V�*詀-I�jE^1?:�_Z�5G_[��}��$��$q���R����3�9S+[�V6�H�*�"wԸ���u`�@pnV�7T)$��\��C v�.t�UR�����W�c�J�ߍ�؄2�t�;��$�v��#�X��.���߶���͒�'!��љ{FP�-�q����M��8aޙ�νX����r���[�mj_g�KV������'=.����z�����e��/rRD��O��"	�)�����w��,��{�z�*���~���;��{)�iٝ��2�R���&n�]�\�IX ����	���J��J�Q��ݻ ����A�W�g�]��?��io�jm�G���� ��Bt�(`)8��G����o�ae�c�[f�?����Cv�I)|�SW��O�m�Ơ���G�߇&.4f�n^6�����[���낮��֏����j���"��4�7��F�rɬ[R�"^p�պ�n<�����a��|�N�ar�cIan�e���V���6l�&����?P���D��7�x�훥
��Y���T� ������5�z�ͣ$�C��l�䘞�QRŇ%j�cn"�L����B_<]y��6T� 5�`�v���͵[n{�d\�uefU̒�����t��b%��6o�l���� ���p�l6���\r@F��Hs�b��G*�4��̬_;G�S���Zْ�n	�d��R�w�^�WD�[�o�%}�x�����9dp���sF�H�֧ͯJ�n�Jզ�]fըйH�`�����2Wo_6��s��Ѯ��gC�B?�;���V�
�q�ۊ��M�9�q�O��	���q7������Չ���Ƃ،Q��}��1S�)�쭍f�O�\a��r�'y�=��*6*���]\��XOb��Z�!{�s]M>���x?ng��G,@e�b�[�^
w�;�����+O0�EТ�Y�u�_�����3�&ۚ��l2<��8�XC��	�2nNԆE�]�2���uA=�~��=7�������T�|�r�B�8��rW���`�bw=Ц}�~��jI�W߰�;2
]��N#�'d���q՚�aA���/�-H�F�kV�+Q�����%f{���*9�S�8�)0��7[�(p���R�0u������"�����V��ye�y�Sn��ݸ�d�~$U��<R�mL5�]��XoCm&�7J���K߼F��(�b�+y7�����IbCR��^kuo�YF�O5�S��-��f�$�zx���S��`vu���w�r�S���Z��dOhy�l8P�����^E:oJ
�t�[��Z#j�5z7Y�E����t
�����7"�2�5�4�ݣ�[��%-3��e���2���(gt���<��O F�L�Dj�>JM��=���8j`�/h����hb���R���%���*��٦�t��oq�D��d�n� �p�"�b��W��������$��qRKfK
�+h[�P��8�VV�Q��
(���.m��k1��fb]���h+�(߀��Pl��#\	�1��βh�Z�*�r�,��>� �6ϙ�.����\��45M�-`Wi��x|�w~�-� |~�p&�zb�o<��H��KΡ1cbm���QC���6v'�����J�++ΓN/Yɐ�%r���-�`��=�;�ԓ���^���h�F�z��}_c��a����^^,fe�S���@|�;�ߖy̽h_)q��u� ����%�n���].�w�L��)�y��m(ÿ���ֈ��
��:fOg̭%C��:;$S���N\�7A�-��i~l"�*�㨇�����N�j`
���Ug� ��:��f��1W5�����q%@)r%n!Qb��'�
�;���`�IXK?�U��YCT�N+�`��[�K�����?8����͏�t3� ���n4�M�4�ajLAXK��N��K����KU㉵%�I�͒3tx-������z���.��Gf9m=��x-�pO�G�6z+tVĦܚ���\N���r��p�����`�UT�k��![�>�<ɛ�E�W�|�n�`O���sf�Ւ}�T����C���nc�쪦�����Ϋ�%bvr��~=�엷O?�{�Q���8XK.�W��[�B�r�>h��),��xx�x)<?���Ӯ`~�o;J>GZ,���Zm��^��O���Z)���: ��X����gU�%�r����M�I��Y$*���� ]ʿ8���]c<��z��2�����՗t+Eg��?�PZ_�dۘ>�v�hx�i���)��o�
� ��W���r�ß��pc���}�}�6�%ǅ6�hr���{(��Ǳ�r��2/��K���`cR����en��ѼC��i��P锓���������0��*�)�dD�-���e���-M���G����.r���Q|['7�QG���se���IoإAR�xy$��0�k��!7��֮媴�Q$F��"(>�|>?�c���^�����~V7d!�����*�	�3��'� y��<��7�}su���rq��[V�/�����w�d���j���?��d�ѻB��Pn��^��_�F�:�BqM��~uS����M��:?�sCݷ�*��)�����s�>�e�{f�§d/���~�c�{��x�88-�ÃN����n�#���U�fE�"��,ao�*�v#��W�g��.�4t=ϐ8��P{����@�+uSn�k<�p�,t��ǜFJ�?W�иt�=�)6CQ᝕H1KP�����aP�J��oht���T��\ɪ]6�p��e���r��o���Bث�������4CϨլT&�U�C~D�0�B�D:�,���7�9,g�/q5�ѷ��%���p�MYI2:�ZՄ������,�N����m3�9.��>}1����wjm{��r�b�+Z�É#m��������f��h{U�g��e\zH� ��$�LG�1�AI�vQ
N]�^�٪-��*��N29���5�%E�㼟��cH�F8]_����Ӝ0���v��7;����b�d61̜�]񌔟*щn�����굃(��w�v��;�������Pr��+�mIܭmkg��ኍd� ɠ$�J�;��m��x�lNl$�l�'���6#�O,S%�p�S@�8��Â�!Hw�
�1�0���?��.P��Q�����WH����\���\���w�!z��Ǿ�a��	�#-Z޿T��O	�Ip./.*Naն�E��H~���j����5�(�!��#q "�!�00`#�ɻ����H�1��>������*��C�������цj���J���#�n��w��s�v�L$��g�Tf�o�n)�<��w��)�Z��t{2k�A[��
7K�!(��P�	�B]��eu�k�|ہ�%��I������?qw�o�U�k�Q�����c����j ��vyWOeq��`�Oj�}�&�:R�M�6 ���a/�b���_��j��U5Tyt�]��a�H*ܜ�V�X�E���2@5��T�S������\u����1��8�G���"d�V�jGP���L#!6��Yt��­�}p0��]Ҹ\���F��J�����(�o���u��oVS��O߽P���5lh��u`窋�)�(1w�(��*lݍ �ƎXȼfo�ofʂd�":���y+�XӸ�!��Vg����S�"��_A��B8�4�i�߈��ui�e*�1��7t]lMy����$٨B��=���wR��:v��V�,��x�m��5@	�=Ym��O�ǰ֏.�i?�d`x2GV�z����~܊rᴲ�Υ�&Ou��D�Mn,q#]Je�"�%�g�IX�K\����U�lyDC��|��s;<��ú6D�S.��9�aϪDH��$�����
Y�_lM��$L0q�:�����C�Wn��c�8�M�2�����;\�zA3��n�H�����?O͜x��N���Sb:�M ��e��k|�N<����1���A���V����F;��y���-�\ӂؐcA�e�dS$�ʠu��r����_P	Z�d^�a|%�d0�(J�'G��FĜ�m�b�STG a�^V��79��z�W�2�<>*�z#�q �m�_�q$�H�j\��E����>=/���w�	?f6��0se�ڸ&����l�����P$�	6���'����^w
� -сy]j�[����+/z݌��,�� ��%���|�M�Qq9^��|���^f�ݮk����x>��!
�JT�]����W��SHQ��+]��qK�nޝtn�7�s�K��Nc2"��])�S��A�����~z���?��K�rm� �����ǽ[�M8v*ˢVs��Pj�N�	@p�����J����Ǩ6v����mH�Jh �kT���z|�� �lkD\�"b���?Z?��{��qӟ�`$�h��fʪ��-&_{-F���rO�mO���ż�ǲ�J�����&ܷ�'�z���b ?-9]=+��[\O�>���KC@c%I׿*�C�D��U�~�v9(�ռf�
�Jˑ'���"���H���Ӂ-O΃B��C;������n����V6�jh���S�z|�h��Ⱦ�q��x��)���A&e�mE9ւ����U��������mK���At�"�Z�d�_�gZ,�7�8�l�Q2ֹ����h�>ԑط��z�qcU2�{0���a�lR�d���@.ʽ�6��Wn��si|�@��Ÿ�sʿ��ǐ�(1]�ġ@�;��j�y�Xr�2v]<�n�D[;O ;�lC��hAT^x��z�d��P3��R�t}���<��)b��$"� t��6���zF��0ᭌ&sD/��,&,��A����N�.Wڄ�"�N.q2{�庢@�����i��F��ǛK��ֽ��Vp��nl�!8i��k�nl����z�?f���@�o���}frٿ~�oW������P\��� ��>K����^&���B2ŦS
ۨ�WR8��XL�RS|a�����q�(=���/8��*n\�# /e�d$��<&dA�xD0�hbz%h�f6��Q	�=p�i>$
g��b"�����qI�j��H�o�h�T�qJ�)�淏$ed�!� ňY��ٞ���*� 3O>0O��yqC�����V
�N�xq2�%�����Ґ-�k�p���b!�SH�9��xޱ�!w ��!A4� 6��k���G/���RJ+f���V�~]h�6ֶT�����@ZzD��4�#0!�/��m"�����ɠ_zD//X���*�U���CM����\� ����?;���Ҷg�]�ø.�s	$�)/������\�p�IM��u�\|W��
�d���W>OZT��Zn.�7������N�����4�fn�)��	L��C�ب� z�=*�C�u��J����[drQ�q�Z�_ja����WL��UP�٣�:k�%,\������!G3uK�8
�t���Mz=��,�M|�Hdi��7�0�%��}�*�;*����U�5 L�I애�fsC���]�*���AIqFrN��+��I"�*����J�2s9�l_�F�=/���x�5X�b�=�V�z�}�C+䓳W �o�B+�Č��l��~���Y��ՋӋ�S��99~ۅ����(�bG���/�ZUQ�k�@��Y�探��Il�&�qx��=��'dq�|�V ���D"�6S?IZ�.W�vi*�J�߅d��V���/�d��N�f��y	�D}S�< s$��)w&Q���,�85���X�E���`SJB��th��JJ�xD'�ϫ�� vT6�	��I͊�M�D�V��l��+��_�,���5�_��E�Eu��]%őn!Dm�����Y x����mUYQl��y�J����(���H���5��tz>�X��x�#�>��j��4����O������g >8`$���yj��_�^�3���>���UKnC�>���� �������l�5 �\T�bzv�M�R9J&���̆���������w�H�&ED���$������f��L�����z� sM��A�804ҏ"=����ne� $�9��\_'`�gdj��\\����6P��u�A-��l�#�N��5��3��H嵸+��BR������]H��za�B�d
����u<Dšn@Iw�����>�_���=oPB��:��� �ǟ�P�)�ei(���d*��}�t�Tܿ�Vg0BO ��\e� �w��&�t�;���F���,j?�Nk�$➠�i���7O���Q>���qlE'�&�C����/���߼��.Ȭ��t���L�L�r�oDM=����P����lA$�~���n%��J�:̼G�W�7O�X�./�7Xlr�n�x�d+�_�]��[ǻ�G��2�k� Mm�?9���f���b���a�I#Ձ���G��2 �"����H�nDch{g
�T�R��"���g���V��t�׳0kH&`_�k��G�hp�1�X��h�0�&���h)�:��XW`�I�|P@���~f1D20�}J��S�+�w$���q,(p� �G����w��8�uPw�7ˌ���ꅊL���N-/��y�R�*�y����gl��?t�!�9���-����$���G��x$���!�0݋AU����l<��͉h���-h�p�z)��k�	���^���B(��/��@�}����C+��8M�G���_*���L��ߌ� $��pp6�y쬩]�G�o�ְ��D#���������s8�S�*kq�KC�S��q^�@��E�?�I؛�.S����R� Ͼ�����_�1�N-����@OV<Z��C܅!�쯝
m�k��ib�#�ŀ�c�&I�?��
�,�-��C�rc���@����oh����a�ot���eƟ>�T��j0t�<�Q=��#�ߦ+��t���W���&����z2�Fŷ������j<��?>}����h��łt�	=�p�b$8���2�5��X�f�ˉ��ANh�X��,���-��X�(���FHnɊr@�r�����@�LeP�N �>߂�Q��bf�[08�i"�������h�����K'��L���i�nk��^)����X��MwR�>w!6�8�;XaH��ʡ�L�� �<�}BS|*!�mD�.!�5�D���̠)7�y��b�)р7;|i�΄;���C"1&�-@~����1gN�ԡvp��c�(���[�R�á��Q$�&�Q+i��>^�i�� `�` ��^Wt�^K@0�xi<W�)@o���-����!�'����Ib�2�p8P���
YR��c}*0f!��T�X�s�b<�Z���&bH�"��46�]vQ��D0� � �}�"��wz�,sj�Ha|y����(F=@����ba�i�+��C��+��d�?��]O�m���r�lJ�n�A��y{J�v���Y�J	�����3�M UE1���aL���uzz$7���� @l�c� �y�
�[h��Y��Ñ���O�@3���v����o�X������<��C6��{^O�j���~�h����.��z�X|��u���Z=�)�xr��n��6��^��A��)v�D���1�}e1���U�I�F'?�B"���u�*|�ST9�]/��G>�8_~��bTD�D�ywqڿ`�
8�W$Y�?�Հ�xf*+��榃�0���{zy��\�B�{_�v�F��+���at�?R�/q�{��~m~*�E*9��O����u@����{�9�Ը��GE���p�N'K�ݦ0"'��,���|��P���\D�]d鋏p��Ɔ�Z��S�xװ�0Uh�@�B�=Hf�d��y�pj�u	���(ohW��º�0G���È�6UW}.,� }��Z�0{����Ȫ�s��+�S�	Vz�q"=�������i9��+�.�C�z�}~D�xQσ�� �V<U����c2�&�ޣ�*v*>����DbC��3�#^!��o�DV�C�I`!��O��t�zg�0�m
&�0k�&/Q@��g�e�~ya��|��Ob�S��i�]��Ǿ���������y%j���YK�R,!��w�4n<���ZFd��^Tܸ�앫R౲�c:Q;���t�g�^D������S:��E��}ȕ��,���(G4���3Zͻ�E���X_�" ʦ!�I�5c@W�y`1�(�cO?	���iՀ�9��C<]`Et�IX��0u5#U����N,�+0h�&c!��D�?;i"H��aj�>�\�2���w�3@��������q �R�^-��i�/<�������B�Z�ؖ�9��(���Ƨ�'4��%	�
��q���΍�hft��nR��z���$<+ E_m�_����Y�p�F�
�h�A�d��Ī�w���uђACՎ�ߊ�5�S���ߟ(��=�@(��� 0�4�E�I�eʅ� ����$]���T_��/�fPj]�jFW
Qӌ�1���m����w�}��kk����P��Õ\t�K9��}�N�ߓ�NR�#T��3|��S�E �����H�|�_�d6* @�3���1��]	�u�g��|��X�^a�|l���W�7�s-���o
���!q�m��o5Qe �x5�"K ��W�A�&�)���34kj��[�늀���L6y[�Y8Hr+@�t�ɥ�sN�C�.ƿl����d`R/�B]�B�ԲA��������Ut�[%���r��R�̨s.�t��2�&�����Ɂ�rx�8������-�P���������Y���p�5�x�\)�;;ŀ��8��e�Kp����%�"��y`�HX2�˸�2d{Tmx?�G���"�� ����{�T���M1;�m98��&'�1��w���	�fH{��`���O��82Sۈ
`��y�gV���){�/��f�I�
��%�*�~�6��t�byD���f:��a2MB�ɘ&���d�ҿ�y]f���n@���� �F�ː�6���;i~сnՄ�Y�10��Qݒ�������Pk�
�J!�Z�<N�ޕ�Fw�*�Y,vpՃ��'��MQd��:�F����ѱM�5�˅�'}0?�,|�p �f���֭1����z
K��FM_�M�h���a�0�����A0�3��"���T�HN��5� ���ü�Z��ֽA�mL1so��Jt��.��=�hb<�7���ܓTIwKB����\%��9c�lSi��7�<KoX"�m��h2����(�N���V�8b/��H%;������14d1�q:�N�Z�T�aW�k�7B��� �_��ҵ|�����c͊ze'sv!J�� �@��o�2P�@���bxA+T����{����󼨴@f�@���.�o����SL���]��GW@px$ू��!�80���=:�:Mőy�9Q��1*��i�]� t�g��ߥ��y�Kb�-���C��@�G�x�S��!�����7>�Cܳ	�I�{�I�$Ikc��g�}��X��� ��Ґl���F��vᛆZX�J�W�z�q_����X���K2ʙ`$*В�w=�d���<�����f	�v�1��E�@�ةS9C�%8IƔ3 Z�i#is�!P�gm���\������;�#�K���P�K\���� �H$��,�O�
���I�X� y<�ŭ���0�#\����]�qރ��|���*�K2�[�M��O-a5����c�%�����}�j�������aQQ�x��U�����U����q�:(rf�B����բ�S��/�x��P�&�r�9��++Pa -9�|AӇ����coM��D��q�����t]�X�B�����e��[t�T6�
@����"<s��9�t3&t�R�Ã���[M�K�֡^c��8�5�v�����I �An�y;�XZ)OgAQ�� ��+4C��mS���r�^yA��e
R��+qv��5��0����L.�d�E@:��2 f���o�ܙ�#1�O��{��8�3�
5
���-����6b9���R</���0I6;��B9�^o3�`Wg�`}�4i���.� oc�Z}Ŋ\s�+5��(��d^�`��,aC���;3��D�/���A.�n$I�F�0"ܭ3=ZAաxW���\�?���#Ti}J��� X���7������-fM�hրFk�>"�[�Y�A%��?�.���	�$��؟EK���Oht�iX<RFrE/���]�a�:*�~aت�����cH�E��:�# ��6�S� D<d�gZ���P�!� ��R2�4��e1Ȩ`0�&������ө�Cp;����	��J��-�o����í�z���fFRF3���&�)%�,ҬA���@;�� Q�ZC��㼅�X��w���94l����1
�l&�V�J��9�A�NA�+�L�����b�]�--� �2N�0�J�E�^D��1-kD�K��|ʁ׃�,�ݖ�H���C �r-��l�����M��<Dp^x|X�8�W�[+�A� >�W����,D��g�0~����sk#�5�/���*g�ܲ~���~�T�*u��I��f���D�&$�̬�RslcZ��GyނZ�KҮ�$	�So��yJ�Wx�f�xĿq��� YnVe�Zka�c�@���}U�8Pv���>zAf�:cif)8ٖ[K�ؿ�f_پ�9��[�p�r0�P����jB�]�b����'n��!��"u�K	��*�+SUL�y��ln-�>�^���'+t)=!�_�j[2�?ڦ��	�����dC�'��I����{�Sc	�5��l�wG:���� �n�� �5!��옒�^�g�iI�f�����l (��{.t�.�X[�̫)9�o�����h?Vt�f�{/z@�BП<�H�R3�^˝�E���D��zW,&�U��-5�
-�@�*� rc���^��͜����laD��9�8����r_:�\s��3��$h�p>Z���v�	$�������E�I��4���S���_�5CL�L:=����m�dr ��T�(\j����h����6�U�C�="�c�{�����rU��0��t�`�6���Zs�Y�Fab��-ʻ�;�R"�C��#,�C U�ס����ȖG���|��x�5-)DE0a��i�Y4a�|�[m$헌�~]pY[�J#�l���mR�Գ�a�*%���<p�T���$���e���]�jU�LqX3���l*y�-��mi�k�XY�%G�b�1'<���m�D1)
Pڶ`5�Q��L��]�7�{����x��>֯<"QQ 0�_4�]�o� qϝ�/ޘ�-$�CȲ��f�`�^����r�#��ۘ޾�3�	ر=,��{��%k�G��`[��V@J���Àj&����@�J���e(���l} EU\�c-?�;�,��2,8�T����Ls�`2����(w�R�2p�u�
|��f(�mf����n�C4n&��y}�n�-�J�n�/�ɑ���B.�k'�@��y"b{�R+_9Cm�1/L�	O��n���u%F������^���D����Ʌ���	��ͻ��Mͯ y�p�P�pp�kE���D@� %���T�*�c&$���<boU�98>�mQ$�[u��*��k!�lڢ26��լ#vQ��1$c�(�U{{�&��'��*�#�j�$������� �v���`�w�-p2ך�)	X�� h�a�B� *�F:�+�2xT�~�{�\A����&.�[����J6��)0�=�c)]KOy����ur��?�㲜?�<W�:�8�3Cm�������E�Ó
n���&_1F+�lO���t�ߣ���QJ��
��(���j\r ��.��L/�G8M1�ƍz�A;[P��U�Zy��3p��J��$a`�3���1��߾�˽�I<-Q��xj�{#(^�R(�M�^�L�ַ]����j�����s����A�V������g���o�7�.�LE�/��Q6������7řN�1�;!����{9��Mw}R����v~��8�����V/p�CU�X�~�6_C��Y�YXX�d.�O�
�6p��V�'h�n��P;ܺ�F�0{Ŕ���*�f?�+{7�a� �bro�k����~�I��&�GW�]�t؏����3x��x�C]�/���hY����D�4�E%~`��V�5�Ê�?�����?�'�΍�����j�T��P�a��ur:��v¼�@��$&����J�Ŋ�Y��xa�����������w�=f���
D����@���O@�����'��"�^o�E�*)6{�%��R,
fFؐX��Z���
ϣ]���jm�V��!�K�}�d��%qf|;t���]%}^�@����v���u3A>�!�^���:/�*c�f}T��E?���+GP� �� ���\�8���>D�(���d��0c�5�U����E(��j�Nr�6v���-B	��4�;�����)hu �kW��g��I% ���]H�5��7�n�V,X.m8�5N�I ��>����΅&e�d[]��[�mSѮ́�L�� ����j�c�
�և;�]+����qv��t�$�����h�u�� �t�,�����(��GO��^��"�9G�X)>����V"qF{+PA� 9i�Ď�?� V���M\ eR��?�E.�wR'�s�R�'��%��lmy�Z�nDp"J�a@\����Z�*�H�iZ|�����=�-2Ԯ�re��=�u�b�F)��x艹�,�k(�Ǎ�6�_#����8[�َ �ɍ�MO�XF��,��e8�3!:��z�N��U��0���K[�]�v��#���uڄԟ ��aٙq@gZy&��#!��G�ͭ7B
E��?���Nb��9q�����s�q�VL��ƛ���( рm���5o�!6�xߍ�j��q��X�ՠ�<��u>��z�(��W3 D��\h�~�:���#��ͷ:�Zf�+�`Da���yz���j�A�񚔈�P<�&|�f��$uՅ���m+6�m�k�{}A���O����]�J�V��R���]?o� ����d�yk<�^�|D�?�%��Vq9�a?r[���1 ��c��l���G��"mYEԱ�����α�(3{o�2�E(rd��p�޲�At�2��u�������u���yޟ��s�羈K2k �qw��.�C�]�Q ZL��RVeN���4m��ԈA�]���K�~�엩u�Y7�8;�Md�}�����������F	]�KeH��Uz%g�T�2䀠�`�;��D�<��.��j�f:�u�؋� ��z��\�����W�T�8x������`%�-���Jcj�Jq�y�	��X��S��?���>n�U�'�T����aaI3��	�悜R��WIY�qa>
L5���?;z����y�3+U�AE�_�%��X���O�������j�'Y�����/�)m�5u;�F�ֻ�E���H]\�r&C���D���ŞlF�:����"� T��b�{2�S�0t}�z@�3�&�9܀D�-�@��6�m�}�	����˘�nw��ƄbUE����ڒ��%�T�9���ʋ���WD�>�t��c�(|>|K%e4�] H�԰,,�����F�_�x$�ܹ�-r�'ka���nU��7V�h~﫸����%�8����/V�,�hq-t�w,{��{�m�[B�U�t�9�n	�]�����|��Dy<=��f��~�Î��N���-nǼê��S:vp�L�<7�m�Nu��7��/L��˜�Fvs��_�L���N�|��<`;P����G=��v�����:hG�q��K_���4��bj����@j]Ԝ ����Kl�e�J��Np�G�xnu/�IW?��8��I��,%¼�6Ӏ�~ؔ�@4� .��\6���=vwxM�'0�O����ƴ$D�rc��  �Vੵ�@�s
#VZ����35˜t��!ᛅ`�X��������! �q�I�"u�&�z��Ѽ1].<Y�w�Br�2U3������'@k/�[>�iu��X�)��kjTڭ!a�j����'F CZ3Պ�tȞ�sUzl��mW�����QY}"�PIE� o�\t1)F	�{�8Ib�?9q ����{�YAǱ�r��5���/�0� u���Ty���+<lSG=hp �O	�P$�Y$᳽��n����ă	$Fu�G��TRF��Ps-kы��CPaqYX��@<഑��s�,���ϫ2�TFö�$��i�C�P��E� 
!��;5�&�����\�6��)�*� ���oq-�+AO�i����zQF�����M @�l;�3t��+7۫��r.�����n�MN��9���R�A�L�:�?j�S�W99���c�l�v'���ej,t@^H]_�IĞ�m֐r��im!��-��~ �����Z�+}���������!� ���,Ҡ�/��']��}�4@7��Hs���ŵ��b53�y*��}cp�-�&���������� �f��n�����=�\(����t�]r\�7����w�+�_�k���qO��6�b��=�,�.�htťD��M���-��5�)�ч�M�mSu�hɕ� �ˉ�|'�,��M*	Y�3Cx΂J��n�᪓�7`Hr9�kՂԺ�i�9��?��z.�{7�!�o�mV��o4i�D��#S{�A�L=
�g���1�[nvRƿ��.���??��+-��֒�,T9,�L<���C M���z�̷�"�!�T�A3�yF��U��֜��0@���@��vYO�
��C��LSǔ�[c@g�z��<�&,kr����y ~�T �Ve��(((�%5nF�]��u��x$�K���lwdd^Z��#�J���g�Ss��P�6}�;'�>�\&�]����}rfv�ʟ��>�������"�-`�ږ�V����)�Ă\{�<fG���.P|2�_�sA8�nAخ�(({�>L0��f�o�>6N�+�2�O�{�E�����U�%}̻�|]\�;	A:��a�2�\�����fL�EZc~�ݸW�V}��3Y���7>���;a�V0b�!�l.� �_ר�B�&�7�&1��PGm�P�����YԐ��O�[�\Y�A��s��=6�Z�������L������Lz���%���oR&��K	�U�~ـ*~�I|�n�dP t(�X�߆��f��a���:�l�Q����?�����bVho��[�vt� �`j��49�դ\�+�l�����E�ȫ�<W˄��Ͳ��j��d�ͷ[-����$�E����z����O|������Q)A>(��K�T*��"��mt&cV���?U4ڣ��.��V@կm0ކR{	po9־B�v�щ4{U���ƀ�֘��՜�c�}�y�Ȍ���6�9��ZM�-p���Q]�\��
��tT�"���\��Jʍ���H[��c��vpd��]��R,��z��ex�?�L ^&;�540 4g��Ut;}�E j=h5����ID�f'���>�#9���ª�9��醏��[����}�Ql7��7�W&u�y�]�M��M�� �g�w�j�= �w~L��o0�^Ⱦq�Z���[[י)��j�"�R�]�B��2��C�L�Ε1�x������]�3����cSu/%}�7QYa�ՙ>{��42乬����h�g�Yd�����(�a�H�&�F����"_�K�!I��K�R'J�'`�K�G-fNH8 ��E���6`k5S۠����*t�! T"*�y2$�X���7�(��0J>SJ1����]
n4T=�E���}Q2?���w�T��A�EƗI4�L�(Є$�}��n� @e�7>9,���l��(?؊�����7)#��T�X��>�lX��IhC���Ę��5�F�~\�����@FP�L�ïQ]�s_�?��t���T��p;+��Url^��ʣ�>�N�����WP�Q�/�^S_^\��k�c�&m@��*��>�����÷(4_v�B�o	�+[�ҷG�ح����z�z��Gj�]/)��n�Aݰ�)Pv#�K<�Ŭ�H�{���ޜ����Gؒ��6�R*E��4�'
��.�O������S�Cgg���u*�b)���v9 �q�	�cev�=������"�� �3ՙubw֐7�q�GX/���$k�(X�������6�-"���PW&B�{ *{���l�bLw����5q4؀:vW��E��1b�#�f�5�����=��n�5E;n�_�zJ�rD���ja�KCQ��e���%��V	��Gu|[`�x� ����n��W���,�v��Y�9^�6��h�G�8��O{��$�Ss x��B�-�$�$���1��ґ<�7�r�'��I���%ʇ���V2{��I�D �6T>�W�5��*�PNb����,�� ��*p�u2�u?C=huh.��-�5f���R~����̙�R���V����%�+��;mл��-.Y!~��X5�B`��x���J"�0�����:G%m���zsZ�u�́���w��AX�e/ʁ[��ևv^귺|�k�
,�}�n�	a���`6A����Me�:F�.����	Oe��>\Ȯ@�U2�xއ̉
��zX���yR:U���#��Ty�S5y@�X�]&;Ή%���Iä8�O��C�@��$2�a(*��&�mYt��]���@S|/�@���,���C����ܔ	)m�àn�ؾ�Q��..l��nG�2@#�e��}�fa�R�D\�*�3�,QBxl��}�M������i��Hb��!Py�1��V4�v���F�HA�%l��v�ʁv,�ێ �K�_u�9����u�U=Ri���	�ЦU�_saJ��k.w|��u~�W���BQ�
��k�r�|+ ��7�)���$�U�Eǌ:�,���1|�����u�5
�fhp��!S]���mb�����w���x���U�=l@
i8�V�=�b���l�|~���3�ݮ�[�hp2�,9[�=���M"��W�U���� ��t��41*����d�{���n/�v���Z���)_�*@��OF���\���KâI�����x�.bp����i ���ͽۦ��]�G��z_�ڡ_?��Q�P�H�g��áEܗ!�(��{c*`�:K.�V�eN������S�fc@⃀�Y#�=���@~�]��{�6������Dwq��D�441��7���D�U�?�@�)9��|����	��Z�ċ�r<�(�s�Dpe%��b�z؍%�-�PA
��F�t/OFLCp22��˛��*��NwVN#�J?�zC94��P�H��c��xsb��]�{��%Dɍ��f�+n����j.�A����qW`�J2�l4����`%t<���PM7h�Ȍ�ap�"���V2����1] v�l�%6%<p
�ga��ͦ��G�(-.2�.��A�gZ����΁�X�4�V�Vs�T�*���699�T����@�=t�����b'�s~����[c�(��o,�^"�ӎ��ǜ7��<�����$`���#O�ۯ�u�����-؛H���ɪ�, K�"w
�(a��;X��t@��Т��v��d����6�&�<��#�� v�q��J�@�#`ŝ���CLz��V�S�)?��f�xӲ��(����J��
�L^�9�.@A�i����6�m�ݺ�+��K�o�_EMPϢ��q��А;��c��^��vDD/(.�"�޿z2���@$א4��y~������^m��|ġ���C��+f,�U�b�d�t�g<�p�- У�����~c�j����$Pa�L�N�;���6Ga�L�7/B<_:C6=�Xa�_�f�r���?i�?υ)�2�����T�O*�R��llh�,���f:�dVo�����
���ZK�ϔ���<o��pBv���<�G�D�����r(��a����7\�N%�y˽'<��hD�A�N6�D5��n���j��Q�A[��k��qF^Q����Q��y2��s��I�
q�Q�B��"�X�pQF
����׃���Hh��T�'Q������u%W�of<y"&P�2��$�Q]j��CO>4��"2���A`�������)�@>����A�G��,Iz�&G6'�Ǝ���
q�M>�κa���^��͉sh"�[�ԭ�2>E�����;�Oʽ�?Ƚ��:5������b��Ba4���H�S��k���(��A7��^?$��tH<|n�'�|-�t��	��a�O�a�c�j]�%�����A�n_���o�N��䡔��y;��hw%P�)9:�^�&2s�y�4D�t���'���5�n�|�xce
�5ΩL�Tu��Mumk����/uQ�JBQ�1p��= h��yuW��b=Q��誕�D�}�O躎S}���ҵ�� ��4��XRj�I���<�]�H2aF���'�`��Q���/V���n�C��#��c�'�	5t�bK����7�@�[���!��Z/���&{���=$�[��ѿ��֏ѩ�����r�#>sߩ ����i[_�F� �`C<�9��q��gݹnվ����sv��@3*���s��|�Cp
����p���b�׾�Y�,"����qz�3���>��X�t\Q6z��$2����_�6���7����Ie`��5�v�j�<b;F�S�ʯOf��5�.}�w������
�gB��TuL��r��U�
Ox $�/ܵPa�c^O��k���^�V�k�/�B���2�Eђ�9���qb,�������B�V��580�Hs��)ykCU���0:�ݎ*���W�ƿ�r�_��&�y:��wv-�a��:Z.	ۻ�&Uz���cWp
Ã�֨	<\��xj����`��s�vC>Y��T"������F�`ܯ?r�V�6k�Xf�6�K�6,��p�Y'|X��eOU9'�K2�e	֭.폧a�6�2�K/@m]8	;#�ӳJ�.��Yʂ�[g���l����L%�T����s�r!3�+ޑ"�Y�T��O�^_�u�.e�Q���{��g�w`��v��-���T��{0�'鳜���Ydv[�|�.����TnO�٭��]oP�0lx�
4t�^�0ߍU{��Y�5nD|�����@���&\Y�j��{���,�9S\�\��kž�������\���Z��n}����3S����]�X�'��������Q)	3����,�p�a@����P#N���|R6}�6^d#�x_'��#F�?�\\�t64��ȃj����s*=��m�$z��%��?ܿA��>�1p�!�c���2�ׁP�5���
�T������JD��rj�]rc��N�e�)���qt������F�j�9���|��I5ދ�)�=�S�A�&cc+�w�$�On��Ҵ!�u��`�������t%���!�d�w�sc}f��Մ�3��0:��wY�R���-��/�� XJ���u&O:H��:�m�]���l�A������{
��6��(yj���3C��t�D4>���Ŧ1d3+���+O<����~�k�=�'Ta�}��]�	f`m{7 0��a��4�O�`uT�R +out��ʚs���e�Tq�{���à@P�
�Crm�A��[}����)@,�� �u���z8���C��J��1܌nN!��5��E���5P��5b&z+A�;�f���݋��)�d�;}x06b*D=�4A�ֈ-d$�f���� �b$X����dV�T`x4 {�bG�ء���"�GV�;/�Ke��Y�M��T�Ԉߋ��z@�d�v��y��ő,������'�(G�4F���p	�l�����Rw}�0�y����0�12�=%����O�\� �e<N����-^���g��h1�*`e)�Jm& 5F�Q�i���%v�7�/8,�� F>g��'r֏�ܪ� ���Ō��mS57i���Ϟ�Z���:�_��P��B��RJ=Gw)��_c�@�5�$;��Y�{���j��������%Y�L+%⭆�����y���T -wϴ'a�s�Y��0�5��*z �fI25�U��]����借����}� ����-%���-}�����r����/*�?�g��[4Ma�G&�ܜh �5b�ň]iD�q9�t(+<1��]�x����.�HZ�X'��{$\O-�	��.�]������\���C�!�O��j1�fW�J��2�%�	����0�u[��؋E#�l[(�iKIa:l��;ӊr�N�����k�ےr���8�E܉�,�e~�g�3Rr��#C�.-�G�s,�L��1ѽ�8��}��S�p����,8�PP+��rP���7��b��A�^��cd92�]k�D���`�smMK��U�����o	aI�	�{���$���=1�0��G��[���EK�?]�$V���U��r����16�.l�c���b$Mؙ�+[{��,���(J�G����*�eCA]0-#gX�>$���Y���e���g�KK�I\�?�ؿ��P�q���̬�w��F���P+a����l!�%"u��w����S�N㚼YkT�Z/��GU`�K�oJ��g����XQ@�����K���������W#�����qKH{7��'�j1J���O�C������}7UJ6nln'�������^�9�:+:
����[%t�f�������误��q�?��N�L+�I��E��j��jG�$W[%���+�hp�0
3@�2�IRO���;Z����Q�(e6:%�ܓ�
�EB���L������fǸ�V�n0J�����r%�?��x�nk�6=����9�1�X�����C����~Y���f0����*Ρ#�0��{�j��>�����([�=C6H�V%�_X��2�e(�[��K�;��X�vK6*��Ҽ[�"���c&G�P˿x���.T!oCS�Ũݪ����7��@\�vP���e_����@�%A3��1�3%
"�.pI��R Ǎ�����Ի��o�K�-[�jh5g�K��$���T����T�< ڪ�9N -�\��@a�Vt�w]��|#������=���|����Dn,<�.��h���	4���64���ay3����2k�����Y�<�1+8�U�@�"x�Q\`c��{��9�U�uwH�d�ә�#O�W~�xX^�N�>=_k�v,�W���Ty���th��$!�	�੻V�Q#:V�
�f�&TYJ�L��
FLr˻���pA觪���]����k�!ϔ2^[S��L���v�~,� 8qOB�t�L�ocԭ�dL���_Ϩrks*/V_e��t[[�v�����Z��7P>$
� ��t��J�]A�UJ$�6�4�x�\�j�9^V-nf����)��Rv���^�_ƪ��-,h�s�.����8aD��Ch��.i���!�g�֬tP6}9��h+���������Q4m�C�6^6h��V��N�FJʛ~���+^� �q�"ba�!��X"��W}iا{��.��J�Vwi�WJ;��n����eC�+�wTˠ�\>+v���`9�s������SVjҋ�����<���bl�G��	ǙK�J�&��U�).�A26�R����@��v�i�e(:�$D�c�e���M����p�km3�FW�R�q<�p"i����A<�ǉ	���f��\i�_���e	oY�`�r�,��,)1P#;�*�<�>ػ�����oM�_��_�bō��L?/ʁ������@�R�{����A�Is������[��|�r����n۾�z��c��y]��b�c��}f��-V����p��ķ9h��b���9�zbj���ʑԐ�ۮc��һ.��`�О"�����>����u���N�~��>���dV�5��� ��3<�W��t�s�{�?���,TaN���	���,~���ob���Y�Q	�6(������
�&�>�,��������A����t����#)XZ_�f�Y!z�'W�?u �n:e�p�}H��Y���&cjA<=	���g��tD����wy��� !��FX�v�b��Uf]Ou�
 �Bb�U��!�0�~�pB:�*�������VN��8���U������O�=K_��-��\����E�p��Pe�of$~&�g�K?͞ �6���)c�s�+��]J�"�V+]nd�Z:T�SJ-yrN���}=)/u"-�tߺ��<�8P]B"0
��c��2<I�%L��UC�N�62R\IW���r�|�xz�]��<�鏅��lˆ0��sy@�����q�]>+2�2�~����;���FBHh{�c ��^��
���^-gE%��p������n?O�,��,�/�2�W2��2�].�=�����y��p
Xѯ:,��i� ���_q1i)���6���w��P8c��̥/9�}/���d�C&~%�f<�cJ���(���Ìh�dU�m>l�e*c����@�fs ��M��f�LmI���6z"b�dp�=��z�RN�� ��e@}nZ�y�a�����7�#�[%a7��󴯑�8�1��Y���3������x�Jמp�1g�Co��@휁�Mǵ�����!��d���&[S���5�n?$�V��E)��R�� Z��.}�N��+Y�(/ӱ�co���H�|U�^q�)�J��Uy�%﮿۪R�u���>VT���1��Z�T�rg e�g���>y���J�c�"Ց��Y&2+����bk2rfH�y�HM[�Rv2w:�S�A��u��q�E'�����7OllՀLӴ 2Y]%G?\M���'9��|��r�C����1�߭������lX{.e��p?�Q(���RV�`�]ak�Pao�M�,rӟ`�%C�M��&���s@�Uy����\�cu_m�#�2�b ����� >�ڰ���t�TZʠck����Sd�vvs�7��t��[��(��K�F�W.�+x��wC�dʥ$�Van���E�M|�d\u���+{���Ŧy���_m���b�(�+�����=�d)�l.$߯ˑ}��~���z�h볣+犬���ݴ�}��{������y��L�W"2;�3a&j�U�|LH>���V�d��;(�K�_A��k#-�,�G�W��0w�6��~*�Y*r,��`�&�iwCX���p�7�lfy�Ni2]�]~> �6�A��OU�̶�[\���c��:�A���^L���UoG�� ���-��3�ܕ�0���|MQ
�S?�T���=���[Բ�{ð̦��|�:cջ��nDZ��t������؉�}w)���ó�q�J�<CX�}��s�Ś)��/�T�*�����<�;�vO��Mzw�S��L�z<iȜ���泐F�������m��zI��!�TMh@$V6�gK��~��H\���TK
�ߌ�'"��C%So�)1$+��Ce�^F�o��Oo��I��\�=��n.(j���5c���(O�a��щ�BޤE��D�Q{�rV�1�i$���.n��w1�v�}���]��9�֕��/��h�ĵ���"�E3��R�7@nLw���*`g������c���t�v��E6:&D��\����O�y|:��]��ub~��C��&!G�m�S����ڽ���_�>~)%P�d���>��u=>W�%A��gj�.���2��� �͙`)������n�9M��z@�Fc�=��`p4]W�*��8p�Fuh�쵩���؅�P�������߉A�6ҷlc-8&F�x�6���t����P��V%f�N���V��Z��H�x�!Z��1��\rA��%4Ϝ9S���_�j��Ѱu�j3J�)���w�W�GO��Ȍj��k���>��?��[��A<bP��&1^ir��;1-�;����C��o*
>3�6�����O�E���܄[�P��g���"���5[������q3��B���ৼ+�C����S���{�M"N� �"9��,�|$]���7U┎4�#}o��u��L̐�K��n�If�O�kW4WԢ[N��J3�k�g�����v1�f"d����ld�=y���q�iW̊���Ǽ�S"뛒*Ν�/Q�������~<tp�Σ�pK�{0����P�,�f��ԦI���3��K���O ��wnv8r�,�E��?uT�w|!�E���J�bQ��\�����wٷ1L����tٶ�a,,�A���]S ��������Z���b�!�7�J��
�0�Q���[-�P��"�[Taj'�6(��%?۲�$���kd:rA'�J�� �*�|p�^�P��C]z��a	���>E.�S�t��D,�w�d���ج�0_w�S8b�&��V�Q��0��&x}�Eޖ����>�ƨ�ǛN�0}�ѣ�h�ȓ\�/��4�2VP��x�/֙��~脜����3�ñ��f�����7h���\A��rz~��<���Ll:�-��w}����h���>�ꂫU���|��<�?3We���<SA1cꐞ�D���ɬ���"�KX���5�؍�;�$J��:	�"W?�M0��~��8���ۯ��O��?�l��"Q��u|$�6�غ����Rd��;G$�s_�Gy*�*� j�B)���3m��\ss۶�ta�d�.K|����" p� �Ù�LT���JDE�k/�#oJ��4���N���U�I!6�T�R�b��~�L��6����K�����ۙ�?�)�[]f�!\�lX��BM����/<(e�gEQ2�~|�#����tG�m�%T����1�w"�S������'��]�.�o�앰���ퟱ��h$��Y^��0�{�Y�e*�<��j��߹�2q��f�`���~�$R��;��r��1R�JO:ǭflF�2~���`m��4
sr>a�쎯�R����|�ʥ�p����������	�u�/e�.?�����9�z�s/idi���)t�tH�	�P�y�X�N�kj[~)b���
J���ǖZ�EO᫄��u1Ұ
y#E::X��y��m�X�H��T�TRF�ԴJ� ������~e�q	�x�Z)E"~�ׂm�4�� ����Ö��:+�5ϊj� ��c�l�F��9��v�:{f���t@L�<.��韻��}V��"��~b�M�D�p[� ��U�j����us�W+���ț�g[������,��U �|Z:j]�Lb욭��m��)C�7��%����dj��^��;~��}ULԭ���<��]�^D�U��㸺Yk�� F��_t�	������dW��lZ��Ҧ��)d�K�=����U�;�#�MJ��k�M^cs�� }%�� �(�I��*�y�=�>�o����%����td9��U��r�ǃL@��>�R$����7:k�ӾN�B?���T�SJ˒�M܇t�~�o����|���f�m1'��e�G�eϻH��o������w�(%PQ,�8� ��^��Љa��-f�ќ
%ibe�t,�iuDc�������{�E1� �Rc�ZQmZ�`WZ��ۼ�W����*���Jm�
�V�[�.��5����H�)�t�~��4�������߻�+��e�1턃��.9X��a��T�1�^�@�����)ɳ/�����|�o-21����w�ke�P�^8`��:���*�G+�:���ɨ"M��On=�<`�x���9�߮�T��M�� ҁ%�$����q݂Q|IgѾ��n7�Vd��
&�����q�}��]��b�l�Qtr(i�x�/��/[�j�i�y���IBx!b;�鼞���'�Lc�x�7j`^�}_u����SČ�+��HYm�GU�!�'�9���KE�f���D�ߏ�U��O�);ޭod��f{� ��7��Y��յ���y��_
�f)�O��͟����p���� �SY�0����i�-�ԄhY�L߽���e7B������kPu��;�����{�{����7��Gr>�Չ2�!}X�Y�K0j���*���VP�dAַ�&T�g��Af\�'N��Cw����:�6�"$�L�
>ۜ�?�n�<:gJ���G�?v��Ǟ:,C��2Y�#Ȝ�H�F�߅`���>C>K "�U�WҶ[�D�g'�Au0�{;��#�J�#%�o����$yx[�x��o\���]��~�5w�z��8�R�!׷�=��PG{�*�Ըd<+&8�ŚQ��T�a�̣zTa�}�$2��������w�؝�Pt~�9aq�}�j=�,�^��',,m¤3Xȿalk�hb=]�P��p\�*�:�+��q��%8�7����>�fm6�4|V��m�}4Ë���5����Cc㳬o��qzK�M�HL�xV�?����uҭ'�S���no����Y��oޣ�|�g9�ΪWp[[�l`R���럏I�*�
iG��
I�A�Z�=�(��K(�(�JjV�mj��<ڼ����ה�bO�}xF����B�O�G<qe˵�`8�1��3����z����v�����Hj�"=�����h��-WR�;��A����e���;M��D�嶥/����P�#��T-���!�?ܖ��kx�p蟨�K�h�P�h���>�wu~s�%��=�c����G<0�����攍Y=Ґ�xD�Z6痬��D��Ű�J?��"b+�����Y_}��Iy_���{��Ʌ?�1�] �U5���K�w;�KzgXR�q{L^u^�~rP;�v���vzB����V�i��n�}Z�0(�>k�h�[���= gZco{����%MrqL4� �7m@������߉��v�y��rcleF9�Hc��zo�Ŧ��9raG4�ʝ"��:+��Z3�6ہl�%�#���ީb�[�IldPE3г����pi��/�Q��c��C�b��G��������}�ʎ��,�f��r�����i��dF&�ׯ����9<WhT'�l�9�eo�>�|.��,rUuHB3O>�#oB��9�zf�i��aw�Jփ���5j�yg�lN-��Ʃ36T~�Sw���)�K(������cO(�vNH�]hR�[�X06ٯtm�!��<NK�i�W�p�n�배9�%���#�җ�&qXQ�D2����A=��i�����:h�OrG�N	ߕl�$��$�o9 �����w8���k��P�/��XA�8�Y�f���H�b��_�ү����h���Б�����n^
f�_a����/N_��"���.��:���\G�0]2��^4�Na��-����^���/�x�{&�6��m�?��5���0����ȡ��Q��EL��(>�ٮ`(�k�4�TA���t�w�t5�,�&Y��⓳��.������f�׾�C+��Sd�*rp�9,��nd{4�d�C#O�^��P�v��wO���$S�������~U�ݿ��t�k������9�hD` �^q>�q���rd�wV��(E�.".�E�`��Ĭ(�%�F��$�~ʐކ�?�tn�+vVQi�W��h��I��Dx�|��]}�6�|�jhmnc���N��E���7���$c��݌�(�_&��?�׋��@V����is�)�N���O��$�.�q�)�g��٫��S��"�&O���^RD�/l���?�xM5ە���g�n!�\�@!ͩ$�?V�Hط�;�W�٭��π~�#kp�Gь��5X,�6���%���D��6�q�t��S��}�"���ܡ%!B����s����j�<�Q��_0ڲԴt�n������80N+%$R�z��MD����W�C����A�n�AT�O7fL&*��W�L��ò�|��,/js�e�/��||����x�v����B_È�'i�9�z߶��Q�ĭ�U�L~O{�D�9�<ˁUB�}��02�䗋�Sku��ڏD%޼�Z(���g���['b�\���IC+�hP9"��{���8���qTϧ�:�7{��[V�{�x�"ׅl��:���d_P�w*�XX��3�8��2g[���=�mA��$���}޲�H'I�s��e������jیY�ߒ��y�� ���S�0�*����p�q'���R��ހ��z[Ƶ�c�� I��*W^ ��x�y��J��%e�K>n1������\��_*.���C������];$�_��_�h��\e���.��&�eM���攡*�0��oh�i�!Jx��&2e�;<S��;Q�� uS��������[�ꤠg�C��� 3�����w�
��]��\�6���T-�.���$8B�\v�����*%yJ[W6���~W�đE�E�0�*{�#����t�
��0��F[q���J�ز$]h���PĮ&Xa"�=�s�(�x�l~���Ԋ���KB��$��F�D��7f�vӅT�Xw�&��7�>Fli��@�;�N�~T�k�"���L� ��Z�[gk��#�kQ��^E6ߛ��x�k5�f�K.�~����(�,ir������P��%��I�\�A
ܳ9�7yB~��4�i ���c���˅f�?w��&~y1	�{��w\��/)�iA����j\v�Tx���?����� ���t�����8��?D��7�=������k*�W�˱J���.� z��V�Vi�zktq ��N��(��X��S0�LY�9�a5ަ�7<a���#6	 ��Wb!5��W�=5��1�WP�a۠�?p�n�x`�)��h����V_֍~�4��0�qXZ����Iu���>�7���@�����6��V����7ը
_WNq�w���z(����+�'�_.�����E�O�`ׄ��j�ʟ<V�G�
��N=��J?:�9�s�1�78Ԏ �� aN��y�${Se���G�u��Y�I��#jW���>g`��<\��P��H3^���,�d���u�K�
��5d����t�?� 5ӻ.�]�U���I{�����{��4��Ůa*y�C�׽�?���o��;�_�)�R�yKAvkbO_s�zm{i�t�ě~�
��t�O�]�&��*&w���^G��;��	x(�}�}vv�<Ir7q��/�߻�t�o�1Vs�����̃�b�~�l&C"r�����W6N*�vٴ��� n����y�Cz��}��\Z�!|���ƟgHH�TnK�X��*ԭk��Z�`�����#�τ�Q}��(�pN�x�u�u(���b&/�!�焰zMT�$�qBǪ����4�[�,][�E�xU��y��3�jL�&��D~���23:8�oL4Uh�0]�IҶ�
���M����o�<������ýz?�d.�tmZ�D��&�ԝ��{%����œc�� �uL<g���;��%i����E�ҡ'<sMX��#��P ��:O����KA�}��b��@��v��&�1�	�C�f{�e>� ݲ�_�[O�~Q�",Ϗ�\�I@�����d��5��5س���{�.�^|/�����R{����78QE}�%��n�a���a����`Aj��Y�v`�B�.��a'&l���F���$��FL��VH���_;�9vpds��muO�]��TϽ�)�zW}B���E�3�� ��o�q=���|g�d��������IЛ<v lo���
�"�O'��D��w� \G�L��ebr
���ʜl8q�ԋq=�g��k���6��&]�G� �f���+>mÆ�b�OBЙ[�g�8%��Fu��&0=�!/o����{b�vxIh����wc�dҼ@w0/B����']�@P���.�=��O'�;����c6S�|��|�OЄ�@Яp��{�6HIm�or��ؕ�Ҥ�'	o��o=/��,]��{X���Z��P�oԪ�2������m%3�y����O��I�Kb
�}ҕ�y�EG���_�������ū�l���4HzSON�*�eTk�!j_�X�����t��b����So�\�g���M^~v�l�z��y�Xp��q.��]��_p��
E4�݌���2��ӄ�m0��)SY����*�D��D����$�ƕ���֞�7���CFn��9��9�#�TYN�h����头�y��I���`-fhϳ��@H�Q���_����{
�Kd4�R��h6���{�;�R,�x��?1�8�t��C6�w2�k���/�bΣ��Z�}f�L�Dz�T�ꠄ楿��eu�3W�k�L��՜���`�N,�t���ӓ�C��mo��k�����#��Զ8�"m�J���Ȗ��)��8f7j�nեh'��03N}ѫ�{�]�Y�}���P�4�^���m��-�<�9��i*�j׮Ox�̸W���'���&	V�����k)ׯ�o&��h[���fr�'d��o�h�Ns�/I�����*{%���lǿx����QW9�l�8�q&������Y��E<󉓣�O�[���A��"z�<�'9T�����`K��;��&���\�i�
��N��OJ�W�<��ɡXkCte��2�D&�SכQ�i����#�V�P;.�Eau��q���%](�(;��]/�r^Vg�A���F�s�[��Xv�+:����w��Ġd�cE��h��F�EvΥ�Zn�&�HwA�H!ӮxVg����|����'�5ٷ%CVi�WQY!��v�02�rK��N��/IK��]���d~m�����a��a���\#�l7G�֭��w}�n@� b��w�x�M�8�9:Z�>\�c��J��wOS��4\��&���V�KڒB�4n�>�l����ef:m�`�k�(���`B��fQS�~Ua� ���f�4S{��g���CoT�������7}+�6��oxo����������W?0WڔV�/t�_IF7���X�V��(�
KtN�|2z�h<r���d�|��L�fRϯ9/K��)�{_�Ƽ(��$��ܓ93��+���u�O7y'�s�s=��<�G�,7�1�'�r��?�K�Tzq�����$q��oy^�O��Ə3�8�L]Q�
��j�j��0"�z������-�\���A�9�)�Đ(  !]����0�`��:��R"�C*�8��������������yq�x��k���}_����@�kr�_z:N"���� i���	��-f\f4O��f�ɏPY@I�'w����zP�L��u4K��F��b�*>�iX6����i�B<Na�b�ϤwD4�/Q%��PH�O�;����)��RnԮ,����Fu޳��1%F��AfG�T[1�}����y�a�r~m� B[���؁¿{������$��2Y�uz���w�>��1���������-��鍧�鿱��y,E	��5H�;6�K�Trum�Uű-Zhy����|kS���Y��d������9}��R�V�7���>oe�]�`j���͵�F�`�lR��R������e�4����1>^Ĵ�_n�C��H\F~�}�JX���i�tF̺���N�3h�;6p	��誵�o�X������"��D���e�t9���TLH��Rw���O���U�C��;r�xC��9b���	�\�[пXC*/����'&��_
K"�'�\�� 8T�iS�E�h���n�ȗKϔ��q=�sw[�y��fAi]��B��+�]��vj��&G�^L��_P|�9Q�I�{+�_��In�=Y�{�LzT|�]����>#VL�ںy^*��JT�TΏԙ�=�l�t9�?`�r�w����	%t����`aa]�����Ăv�V����5/~��ۂ)�C8�t�a�tɯX����6��-B/�]�v\~�#��1�Oe$��訝�Ӓ-뮖�h���b���&�j$c7j�ў��ܑ�c��1̬��6p69�[ݭ��E@��������kP�5\��,uұ\'c�6)����c4=�L�e4)sBNp����Ғ d����������������b��d.�$	D�)/����m�	��#�S~oi�`����$d��)���7���3U.�!�*���,���������4��oE8bzG��󷷨 L� ~Ar-�W��c}>@�V���\7r�j�H�[ �X�ʥZs�VW���B��R���Q�ޝū��l3�*�� 6L��A|����K�����,{���c(ٰ��6)�~�+�?L�AcU����2v�T���*��40��U��C���R�ʄ�v����.K����J0�ɫ���C�ˈ�����/q�D�{te��/�L����wk���?4�Iz���&���g }����]O�\"�W�B=�H�WR���-R5	'sO�1��#��	�����{���U�|��:���042���Ux��2U7*(+wP����mߖ$w�����:Ԗh u���)��.�3j�q�deZ��'��f"	$������w��o�R��P4r^e�2�N"��L�L^�Q�D�^�׼m:�{��\^ݻ�CzZ�ޫԂ\#��T�@wc��:|FUu=%RG_/Ap?<z�`�l�S�4w_�Ш��$e��&6�YX���&�m/��ЫMz僫�+g��"��$�8-*ڠ[���Q�X�WI�m>��C<�-0�*�0i�^���ߦ����X�{�)�^�6y�YW'>�L�#���p0����7+�뻮�,8�B�9��T���́�\)���q��I=�Y0�d5�#�G�tp@ɹ��Z���^��L�g���u�Zu_L�����|E�6�Ț���T6��$,�B�U�W��b�ѓ�y�������:�;��Km2�����?����+i�(�O2q�Vɖ�A,����q���co%��Ik嘫�;�'q0h�,W,ʩ��01�8��+5m<T�t��a{�g�� p.nZa����V>8;�� ;���'�nrQ��܊0X2���7��
m	�"���ܗBr'�|l'S�V����$�H��^N��sǩi��*Bqח���lG�W;�^�}�r� ����D�{�B\~q��D���L���wN��� ]��g�q	���v�vܶҔmL�̂d`��HbQ�b�o��_"�_-��q�?�U�Mw�z4+��V�z���0�^�d�q��`M��SI� ]i{�y���#}5�����/sz����ܕJ����z*��ԫ���\��LU���8I�b��$d��i���6�g�U����[C�*9w�O��-�⇋v�8+ �f�����`������8���E�<����U��L�O�+߁)<E�j<]߱@�z�c�w�&۝��_����TzP����kQx_�p��&`�� �k���J��N��@ԙ����b ��]F�*S��G0��p�"�G1�;�.�:��i���Y��g0�'���(,�V
�c��h7�Y�.�k~�Fy�?Ã��1j�(�'��R/|R �������;%I�n��T�j$���tb�ĺ�����4e����a��.¡�3>�0tyxw9H9�Y}ǛH�0�:E�!��nŒ��B�S��mwj`"���9��_u[��w�l���R"�%nW�s`�]��P�'�2r��^��+�vfMW�a�%J6Z�h��{t��n�\�B�<��,̆x[�WC�CՕZ������*(�G��i�	)�!��"��f#�}����y�=�lM9�V�W�q�v>��[���HC�@p�;�U|P=	�1����@�2����h�yeA!F���[�)�O�*�񦿏\d@��HDD�� ��d��O�:���p�piw���k�᮸�v�&4��)�9�a����ef�� ��ᓹ��i3�K�\�¥]�ժIc����^�Z��R͋9�+���)xwc��j�����X�jZ�s�����j��d%u����HJW�]" !���p����1��%����`P����3��^�X�A	}�Rc�������'�ch����z 8���T�� -2M�k��LTbB�F�����X����ᘕ}�LL�w<�Y�<2�`���ݠ��Jk@��{O�˦ڰs�u�].��á�]��:�^�f��\�w��w�=�t���s8$�|^�G�sw�}D�*Nj�|~�@�>f/Z죏|�Te���/S5����eGp�~4d7s���e��'d��8��O����L��B�DI�IK��l���xwo�'$�\+�j%{8(��{������7k�K '��C��N�?��}�-�.O��byQ�6T1;x����F9e���Ѷ���L
�����0<5F�������8<��VւuѡI\�Jt��ӷX�aXO�r �;E2X�;-�I\�2ֵq^��4)�ߗ�j���;�@&F* ��1���ss<��)��AU�W$�29'��1/�QQէ�MЗ&����U�yC �1���Jj�7r���X@��Η^ݎ�X�~U�r9Q��R�n������H�,��ƁKџo��"v��@�K�7!�l�:~b-����a���ez�J��, \��^Rjb��H����W�Z�0m$;C��`�8X�?1w��
��zog^��@Z��c�C���-K<y��c ��N���I��Sk��Q�׃�No�h�;ѽ=M�y�j������3�Lȶ�A�j9Sb	��M@����],���0?��{��.��_
��y#��A<��I���z͢�s[<��G����?� �����˩�C4λ��ݯ���έ��.Z6�w`>�Ƌ�I]�㌦�����
:�p���ʮ�0E�[��v'�Eڝҙm����́��p[<&o���^�y�*W���	�Q� ����?~���@�~nq��YE�Ηg�]���I�,�ǵ�"�M���ۂ����um͹u n��_f(� �!λ�i�a=i����
�-�F�W.<�_���Q�*dA�0�&-ҫ`U���g`y��zfMUlLC=��e׻��NH���8�T�����N�s`�HԎO�i�{ƫDZ`�A�'�ut���~�OL�k�,��n�G�� WC����%#^m�Qְ���n���4��'������Ԟ�L�($�s�_�4|�XR	�`�2�U�[AY���4�d;���S??9_l8�$���U/��d����ś�\	��/@˔��h�j_�~s��y�2]7-�g�>�`	�~7h/��!��Q��w�>m	n���f���U��@+��K�*\9������_�G-�
YsU�s;H�,W���7"�pW'l�܌���;�s���������oT��b�@��'��"_S�y�)�����H}V"�F��M@w�(4���\6D���B�jxp8��	������rh���mN�i�o�[��ŉw/F�.�]��:@𡈻hq����h%k�u���@�*�N �����{�� ����� .T �J�8:޻F�7Y�n��0#8 i���B���)A�M�[��ѫʲT����_�f|�95�=K�l���:%�)v	�۴;K�J���NE^��\���"������FC�oh�@&�\�Ur�s�X��"@}DT�u%��ݨ��)��k�Vb�*/��pD	�{�n�N����U���F?{+��?	ζ���d�	�/4Q�a�?;�`3���x`t3��<_���[T��2 �a��5��Ͱ��_�4R��3r��������ݯ
�z �e^��dX��oZ�t��
����![���2p�WQȊ��ʛ��D��&b��q�[��;ڤT́ݓ0Sj0iq4)_�\{U
�W��yR�2�
�S�e�W N{&��l�#�_�K˓ԿX.��6���Hy�%��y�Tw�3�÷�D��Gž+gn_&�*�a��cR�=�w0qI܆`bX!bZd}���}����F|�eQY��qt�Zm��]+^ '��D��o��y d�3+��qBP�C���s�ΏU�T��U�
�	-���8`{��lU7s�� ��:��
�+=�ò+?�`P���cB|��}LHؖ����o}�)r!���B�AٰB��3�����8���'ڢ���b8���p�V(N��#����=���� �7�q���dQұ�q��S�|��9Xt����֪�yXu.�m
�A_˗���o�5��o��H�b�x��Y�O� ���v��dW�i#��6�o�R���{I׽k˺�VfD�!����u楒N�C"��+������;��%�`d�����bm�~Q �����X��@��ր>��ĳ@Čv�}t�`���B�7�m�{,:�֫[�Ԥ+6ʩ�����zx�1��3,��M���/|t�6���w'�V5E��!���>����n��ޱ#b:����A�����<�C^���[�"k�Y�������Q��z=kH���΅&|�����9�����ٵ%�j>�4'����V�Yws� �v���s<X��Q�5x����|���EBk��Z}���ʈ	�9ސ�Oi�J����Ψ��M���3`�U5�!��l|�זb��0ӻ��ĤS���gAŬ�.:�Ǹ�aIUl��t_��\�Q ��k���ø�j��v�i� �s%��4���/iN���>���2�E��E`\�7��K}�\DbI��0ay>��:��+�#}�ڛ�ê��C��҈E/|�W�#�����h+�N�Dn������s �r(R̆�q"�[��Ce�����[4�t�3�Π�[�CJ�Ѯ:�&٦��xWa�5���F�YÐG���|g`����ڸ��_ː����jܾ��1���Eߐ��h$�TN·.<r��l�6��v�kR�i���<-��g���D'��̸f�������ϟ���G������o��ock��b�w_�#C�����׶�Vr *��R-�7�@��ɋR~�8$�$\V�=�,=*�����\D�Z�D]v���N����7z��Iz�������9"����(�L�R`d�C3�ܖ�5}�a���;��> ��۲���eˠ�@�t��O�h�10����35O���o���vG�$��ص�'�ʔ&��hS��P>x�ќ> ���8�)��u1�y�I�s�sփ7���( ~?]�Q�Y��'S���v�Q���+2>����=�c���iba'�;�\0�񮎇�R��B���Mk�����c��Df̛���������Ń�������X�e����MNa�UG� ���'3d�!o��e�>MMbP�T���F10�a��_qZ�2r��Ｆ�����-삿5�Dr���PW}ԽG?_�c�<|�`]��f��J���q)���cR���xG����kuo�O3�z{�J$>��NL*��;��=?L���Q�������WSC���^�����y�>ͳ��;������H���oO�IQ`�)gD�mo|L�,��\��1�XF��a�iþ��֔�y+,�{{�q��xe�l�W���6 ������Eus3!����$�;tBI��?j��pS�r�~v'L ��Ӧx�yԽz[��}��R �?�4�`���t����)Fŝ6�?�M��
X�:��u̜X��(��U����1if.U��`����@M��5�� �6P����)��"��se8v��������ڿe�����L���f���]�V}<�ً֢�=
~��`�S��zi{��3Gw�F���2��{�s��Qp�G��oc+!0����hfl�}����� �X@0T'��4��ϫ`%�k����7T��b��Ԕ����n���!��t�
)Җ����sUNGs{���ܞ��r�F����C��+B4�O�LT���Z��_��!I�؈4O5G�$/�_I=)�]飖�,�Z"/�$k���Y�V~H��>���&D�k-���@|��}���W�.�B���NK���U�[$L����B0z�H�{�H���g��_+B^�h~�R�WOGk!j�:R4����I����=�ŭ=&��޲Þ����[����#��#�RAe�^�3z�:�+:�u�־F.B%+6���������o�i���P�kJ<젔�ΐ�O�1*�Y�n	�}�P���31�aJH߸k���1)���Iآ�C�Z��0���
��ڬ]��M�J��ƶ#c�M;+��«�Ljv���3�흛)��<p��?��=������T�������^�^����V��C���P���8�Yy��g��L���y؃+f"��*RMbW��aN�Vu.6��OW�Q4%p<��rD�R%���T�
�z֬��o�(f.���[|�oX�E/��v��ga�p��%^/�|��W$h	#󏞫Y�&��u��w�ƽ-��gk�s�i��-؜&8:@��SѾ�xp�P���UjC��ꞵ06zְ�C��0.�5��3 sZ߱�u+�w{͈�2�p���2H��p3�}2�@ȅ]&���]U[.�2���kx�d�'j�e��K2u)�tCb�	�+��s�+���dv1Z���Jme�E��_��S6�z�$��������$y�1٭概�&$��!�W�pv7%�p��<��j�ER����pe��4: �����f��`�� '�������q�fMb7s��+b�5n�.�dm"Պ�l�;��o ���y�l�ƚ���\�W))��'2����E��Z(�X�F{�^3q�豺���,)��5�L�8R��1܋���*�@&�j��5p�_�,���8=�s���"� ���lqq ����XNL(�h����sk�_���v���I^{�7�Oy��O�)#"y\@3���\�B}ݾӶ��P1O��|�XF��&�Ä@C���2銞X}ް�2m<��ئ�[Wv�e���!���E��.mW!�]5|cA�70
��9�L����z��K�x����C�sK6WT��V?�	c%�+7+�*���C`�vdoL1sO�S@ƻk��W��V��~k��ib����6:��O�������,�R�_���@N�/��\�w�/|��T�����]}t�Q����5�ZY'�p�J��6�-��Р��m�Tׇ�y?�15cPRT 3p�k�o�y�Aq̲w�'I�f�'��������;��SԳ�W��p��wX�ʷ�Rh�^�t�텠��(X���:g�Hp�o���mym�8�� �	�=�����x���0�����ʯ�M�t��|!���=�_�>������/C����nm�O�}|�,��Kާ��+|Tx���M����+#/�^��E���uA�%��r`��s�.�U:�by.9�54�r�ɸ�˼�Kr���}_�܍��Np}���cy �V�����đ<F~5�h���H����>M�6Ʃ�3�JZ�?�����(*���}<T��|�vuv%|{4Oml��-��X.�9?MQ������/p��'V����>a49���V�k�3D�"�uEŶ�C�l��x�؜V��5W�S�w��F<('��
���ʒ��W)wR�����"�ޯ����/H�ix���X]]�Y���ۇ6�W�U��{�=	��^������1^�)?��%�&��Q��&�$�n��F��o��M���AL23v���g5��g�y�-��:�&5����!��z��!<�Z��`���p�?��~�֓����o��\s�@0t���pX ��L{g��{ŝީezB�߁%u�|���l�2lTZ�H�ٓ4z����dg*�Dh�t.��ܭ���!` MB�.�w/fsqk�����g~�-�uB����.�U�b{���"�v4��=[��1�5��A��ے�/3_�=>ӸGG�{�j|���I�T�^��-\����IӦV�F�b�����V�g��+�X�e��u���gW3]��i�5�O�A1��ES���r:��!z��H���q�2K��(��f������G�S5'����N�I쏱U��v�@�&��@�7���a�s���6���|+]�y�a��~�3܀�ڻ��'�}�'�!uӍ�Oy�Qل_{"�a�^��r���,�Nrp�}D��F{�GOZ�A8�������/)
����\���@2r�e�2�)�Ec$�,� �������u~���؏9[���S��-R6+���wm�&q���=������VH�P�?1�+eD8K
�bhrT��a�&�_Mϭ�}H���̫ݙ-e`�s	n��ķ�e&���x�H���E���/�����%垟:�:�Є/��_�C�>� Ա��WcI 	r>��ѫ��`�������#b�
va��bX|��T��g��۞�ڀ�$DQzy��9"~��v�l̋��ů2����Cd���>C=�1t"}t��?1Pa��/����v_��i#���	%�`�~�;�����VH���0-�j��������G�a���?������G�N�N�����{�|K�����c�o+���� �}d��l�M�؏��<�
$���{�+�N��ȇ�أJ)�r�[ٮXF�e����w䙂r�VOĞ�Me���^�NwV�Qr>��~*&�|"F��`* F�'�\�ri*1I�G͔������������)�NsT6J��h򁋏r$����8�rfH�i�X������Վ��8��ޠ�J(�Q��M�\l�͈Oߣ^�Z�&B���E���r���Ѡ�I��D��A�l LƠt3��]�r�!fh��]����k�=p�K�O�A�%Y�r+j��ݸ�������[D݋�pǓ{����Ӯ��e�S*�7�i�ob�?_C��7��@[²WշC�_��oiɰ�l�����>��B2���|�	��X�Hqd>3qS�©�����\�
G���8�E���3����z%,�^�����a
���J&"~�tV�6 ��e�Hk2n)}�/+���6",�R�6��,(M�ٗ̐������(����U�
� ����;6�v]�j��"ІA��2�[��C��E�~�)Z�A#���N}��A�vC}�-�Mݏ+��%�J�}+��Q2�@k�("9P��2?�M��/�_j�o��j�τ
��xC���}�4 ?��9?����7_�+YW	�Q�eF��xSض�;��K�6�J"��3����@�y��}�a̙��γ���(��5�-���v�����/n�4�?J�:�Q܌9�g[`��Ď���;-1�F%���o[� �UGeH���s���F�S\�������7��Hl?b�"�~��Q@�Ͻ�kA�H����g�D�����O?��or��k4�}��P{Ղ!�&n�KH0�;t�]�J �=��r�v>��}�����2�w��Δ����:���*���]��h3
C������+�V_�e�1/�������t�*͘@`vt�U�R��(�dڠ�����x�<z�� ��yL���������3亸R�8&�^�c[� �E��!�|��M�W^�Ϻ𤋮Y,H�������A��YB�i���JKO�~�ww\C`�{%�U�@)X�\���;ǟ�4F��E�,6��$�>�k>A�$K, �L�V���S��[�*�;T�&���X\6Ls4�9���}�b5$c.�nt���4� �@h�H� %G�*+�%mHr�%�o�R�cQ�� ($$;]���e�Jx �4`��X��e��$�iZ)��`���#�S�X��G�#sE�D>B�1���4��s���y@vn���W����	�1��Hc����X-��9=A���.t)1�)9�-�<�¾\����eò��W4���A�x�Gk�S$s�^�q	����F>��S�R��xG��4��p�}�H4�'ڰ��F{Ҋo!O�`��?r��Q]@ �c)��/p�eVH��쨇�E�����3n5`��˲�1�J�j���0�|�G�t�,�O��;u���\��w�I�~Z����+�z��o�;��6��r�̃Q�G�Dtͱ7�\XEKV#G��7��g��=�
�.®*�NT<���_��`_<��V[���.�^�L��˚�v~�YC ��u�b��"��B|눫���\�{uŰK�I�%��$��i5��g���]�����{`���2�u]+�`2��U��\e=�G�g׼������aj�( ����N�チ��MO���ג��f%���S�}��~�w���L��O���Ѹ0�Io�vK�SF��NA���n�̊������lG 	\�	��p��9(�&Q�Nr
�ɷu�(��ެ(���3Of��T,\"Hr�@��h��h�5�80��̓Ϡ���F�2G�ĈU��MF���oy%�3L�˶�Ps8�3,x�
�z��_��­�.B�BW&�)�ϫ�.>�*B��YP��?��!���m}A���Hw����Ƃ�e,�y��eH�Q!�sF�<��w�Mҳ^qvE%��Fe�����:D-%�_=��lH����[Ȫ�w6��ΝѰf��������kk]
}��	26hI�?(K �k���\�7�� �Y�T�[�>�#�)c:��&֍��'���|H޿m�k�v�!���7�R�0����1)X��l�ت�.x�|������s��+��E�KD't�~T���~���������j�����FPq��~(im����@����y��:dl��[7� �(S��Y��-����lv�P@�ɍi�J<h@�3�(�?��Ђ͟�@�%�|W}W��/��InDK�w;�{�):�|�BO3��7�g5#"��R���0՞�'��w��?��eil@���$Jb����/���3U�q�R�~ژ��Bz+��/�˻z[��
7���K���،2Ɋۀ�+�ŀ?�ŜQo�*�>��b�膞�x=]�T&ވ�����`�3�(��+I��6���h5��.��$���iB��үq��J���*n]��Ri�k��-��>KͳX�[G��n���@p�iTj�%;O�焼.n�����S>��f��'�,�p��Rn���[��W��4E��6�����w�%�֚;y�p��w������'�$8�('�����qm�z\�f��#eN�F�[ ��8�E8ס��K�z~�v:��\H�
m���/��jy4\N�
TV���0��|+���8)�'%��?s�T�^ ��Dt9�t\76��Y�N>��]���������Է���@Z���ۡ�j��� �칹�.7m���|B��J�U{t�? yT>��8HKK=~��c"�pFf�2{.͘t�39����J��K����Ie�ȇ|�cm�S$�T�W��d}�0W�a��Y%������r����v��TL��s�N�>���T�g�.`�0B*�HLN�?W$v)(��\8u����/s�'x���J�	˓_O�Ku����� ~/SQ7��m��B��k� �ֶ���)�X��@;�R�:U�Zy���$=1����|6��#z�@7(q 3}T��L�5�0�*a�_�@xȩ�Bi.71�7�=z�>z+�O�E�@1�(��'=���up"ϟI8�E�WY�����B�B��~]��$~_ڷZ�Ɉ7:�g)���|2���\a��j���ú'O܉	�ܡ�R�"s�X�h��$��fR�����Ƨ3���H��\������B:�-�n�p#L"�WH�4�����P1�����Q�ا�c�9"fo/�0�}r͓d]9D��
�^,�I�bl���u��T��%��A����o��#��p����W$��N�5�د~��%�j�=N��*?<b��RH�> @%}�_%=����`$T�ǋ!�0���Iv�D0�#�i"9RЎ�h'qk
�ie�]��D<=�y�#{�]�����|��L�|Zv�?�N9s�7�$�!r�y; �z��n��|�W�vBf�ͮ��S7>��)Lх�efG�W��X�z��r�Θ�8�{��
r�Ω� �KP�Q4���5#�G��;D����l1��:Ă?{�c������}k3˂�ZU����ᒨ�^[*�?}fy0��']��,&+� mz�ͺ{��l�C����Ow69=��X++HOȤѷ!�������m�Dr��9�|��E�gҮ��u���mfu�B�v�g�ĀPK?J8�dM�jj�i��8�i�nΝ`�	3�Ɯ5��׉��zպ�G�B����7��
ӕ�tSw�T��\�5(D���lY2��y�@�}�	�k{�Uh�c�1�_/���S/���O8K��i{���6Y�tV �Ҵ�s�տYV���A��@��Aͣ�\���^9��_�S9�:���Yޕ��ƪ`%n>g�Gl�a9�����$>���h�ڑy��g�Ae���ρ�e���r�V ����1�d<�8�$�V�S�W�����ݽſZ�o������h�A o���]������v��$����᷊qMى,�.1�S	jP���朾��m���Iu�o��o��V��ւ���Ԑ�e���a�n3CX���W8�c_"_{��[�����O��*V^V�p��Z�2�7��qU0y�D��f�(%�_]-�t�j��*��s1�{���}��O]�l���Q��X0��y�=�ڟ.���\8�^Oaߑ&�*�"5u�m`�#2Q�:������_�7��o�x�xo��^P�B��Q�B�Q��ԣ���|ĵN|a���*4���9��1>-3*Nt�����Q�i�(������a���i~�"��t�������|�����v�~��u��7��� �\0�ǣ
�5i~_ ���:'$�W@ݐ(�����U\�A���0�9j�bʓ| X3�I���~ձ���}��R�K��Dx��A���>�j����� �
��Z�t����A����=��+�eg����?E���l�T��~�p0�d�֩��n�K�G�_�z<�P6놁)gB������_��B�@�%��v��.���!CŻG�eĠg�}�+P���_�|�?���a	D�Ni�R󛡵��M-����G��x:~�'e)�+M��+�Ϫ����D��O�3=�Vx�j��V_�*o����gq�u��)W\��#O�ڻ{쾥2E��&��z������e%�<��it䗆ӑ�z��IA�-@<˕J��2�@��ݘHd�߮�5��Ԯe�cwjD�l�O�G����U��b���X��4��KHx�s����~?���s3�^&2'��G( 'T�W�ܦKw�oa�Q��q�h�>;`�۲��� ���}j�{�N(�W�
Y��P1��{'�BJ`ק2Q?���`߭$�b�{K������	8$K��<�
��~_FU��xt�NնH
�Q�dm]b�\!`�@?%�K�����6����#���?�U�>��Fj�Y���qk���@�X�Vg����m�酒�|����­�4\�+���&\,���זt��e�ղ4��X f���t
ĜP$���yk��-b|�0��B$S_rh��jt�NP��p����F�T>��h�w�M5��!����ᕰ�T,�+Sݡ#�6�[�H��D���=
��gm�EF3���m�He�Zܯnѭ��qb�+�]�Q�i�����0m?pŴ4��V������8=����5�rl碓J��/ڽ��7Nj��;��*�S������Q�\`?��K�,�
��0od&��?�*��V(��|�W��vv�ul��P����H�ڭ�澧r�(��ϫ�'����V'��T7��|�3`/��U�E�+�������e�t#�o� �S�tn�IT���|�2��۩wz�2��rlǮ���2��5{+C��Z��a�g��^+uD����'tc�7�;29�V�?���v�fttr�����W<���cq��ÇI�
��*��\��_@"
s��?���b$6�(����Z�g���ȩ����4���K�va�?aы���C��q(�zv`�{&̍J���̭ta� 1�'`x�	��*	�x�����K�e��+$��5� �u����7Ύ��L���+=q�T�+k�c�,i� �,������`�hr ��^ht"�D]�����b����Ѻ�	%i����o�g��<D��S��U����#��/`��f`umխ�����Òt�����w@�����3 b��8I	骁��;�M�@��}"�Ւ�ǜC�j߽Ժ;���Qٺ���Wn���I��f�Sqg�O@�Y*̛�y{G,t��G�2�2��K:�4�(}<E�}��l�C]T��ڃ�!OȬӓ�Fd��˓#��o��"������E�F��2��t��8�~
#G�bQ���!�k_*敁�?��E롯nM'�њUYڷbQ����+f�������s�S��?�TЫJ#�&�9�S��]v�i�0���zaL�Õ^@��~ND�	�eܫ�a�}b�� |
>lvm�e��e�Y/��J�M�x�;���K�,�e��@̋H ���f�e��p �]I<���~:O��a7vm6�l�NvLRf�[��Oܰ��ү��O���ҸF��-�61�$�ߧ�%E�l]������2��:
�-���׍�]\�I�����dN����n���Ե{�B%Gj͵Z����ȓ��ٷ�A����H�Ub��_+:�~:T��/ı��h޵����o�D���<|�*�Sjh=Q'=b�(�(e��
,�mڗ	��B��{v���`W�wK�_ɀۥ���u��9uؐn�c�V���z18�*cd��!�V�F)���&8B��;,�rx��wvbt�bL�!ZjM�WF���)� b�nT�P\��� DUn����D�K���]��ߵ��Z�U��J Q��~�N�R���=:�QY���/�2�Ţ��eޓ�O��Ȣ����\н�;�$�"�[���@��������1�Z���#����գUn�7�	xU�,,J$wv%�>�?ǵǟ����eQW�p� nَ�#g����İ�L�T�u�|b?�������Ғ��>���Z��C �� +���g��[U��`aebnO�鼌�c���V�YwR��Q�m"g/kÐ������W>..�m�>��3}@{�Z�R�����N�8���D-�"�N�� �������3�ߋE���6��������G���_���`[YI���G��[oJ�ö��W��UFp,�D���d�>(>�)k����]J�ȃ�+����}�(g�B@<��F:8�y�r��y�E$�EM9�֞+E��3~���|��ىD)c�DIO%m�|ie�lU[�7t�����W
�á�#3eAR�1Rh��X49==�e�/����+�"T�)f���{r��գÏ�L��,`X��L
O��`k\�4V��5Hm�q f�q�b�X���U����7�+"������%���;�a�$1'q1�0D�'��ch�}� n��FG��ܐ��N��%�Q՝�:bv���t �8���g�Z��غ����@�@0�[h�+��r�E��������[b��lW �c̔�NT��z��*��K����r��B��x������L��)Le�l�r�+u��0�j�O��D���նjp�~�i�iJ����
dޏ�^3���ݟ�+�T3$S1�@��d��z΁�Bi��x��Lz�)�`�(|����wW���[N��������C�ʬ|fJϯ	��q:��W� �����%���{"A�<���- g+޽�t���K�!|� ��懪�?�h��T�9�_X������ޘ�f�@��8����uC��B��7�ׂ��4Ъ��D�~R���-���[�� �j�Ya�ܙ����U+���".�kO�0E�$����R���E�([<���}�̙p
î1Wo����0�������W��y�\���-'�������� 6�t�$6�/sglg�[+���`�b��-һF�h�NOP*)4n�`�W�Kkiw)�C(�T��0�A��&R�:v�²�kN-�P�x/"0�w#����	ɹ�_VnP�5�֤~�
���&*
��/��l���>���{W�XsK�/���}�H��ۥ�
ZRB~-��K��z�`yٚQ�Mh�ݶ�9���?���4�Xy=6�z� �$>]YG�k���n�� 3����ծ�08��WS�������9Ӕ�)��g�b�Sk
'/���<��	�P�򙭛�
J\zeɁ���.v�� ��Y�o�����ϯ���y��]|�Z3�.��6��#�&��L��=3FQ`���!���E*�|g?�񏩺��Mrk��Щ*o��U��T�?J���j��#��T1D	���m�<�~�:��-����qc]��ϊ�oz����Z%$����8;��qfL{�b6�_���-t��Y\L��
(F���u�|�>?s�q����I&-B8e�&��U����fgo��I�`��ˏ�zr+������z��p6��.UK������`k56�m�sF��(KZZ���f����_���Z�=	ߕu�6܎7��˞|&dp��V�<� �諩@���t�=v[x�/�p�^���Ȝ��7�y�+�Z�ޤ�m>�tT���c�;k�"���H�޴;w�a��WM8'����^X�a�/��x ���5���n\c�'�"��4��8`��OQ��ʪ�M������뎇���	�R�%���JQ�(��y��eg��J�K�d%+e��8��G�8��q��~��~��C}���k<�����<[��>QxdY�����S���%9zƂ=�tV�ĝ��w�8�� @�����G��K�%3]6�f���I�Ŝ4ܩ��Z�x�{�?�8a���9洮�� �2�2l�-��M�M�8��"�m��K 1�J����>+�%vd�ş�_�-�h�Z���q�=���. �����	�k=�}(��L�J*����n��3�	h��Ӳk���;A��Ο?�ټF�V~��}��d�͙E����W7���h)�^��L�����Aty|�����Φ�?��
7%��Ka-�p܁�tϳ61��fƭ�R�Џ:���J��gi�Ď�M狡N�i٠1�GĐ�<���U+|nS���6Աv:*��`W��r�Ku�o�v�]L}�@����8G��ͅ&�~`'��q	�ێmk��O�]��f�����U�8}�������-�wc��P��x��e�?飬tP��w"�l}x_dDAn�~�hcQR��<wus����K�g������KO�3ݽ�x���ivG=��Kt'[�u.t��}ȿKW�����o��o>�M|�y}���sQ�����_�;ބȤS�˔:�%��;w0w�ơ�֔ݙ���?hz33���'g�Lְ``'m�R$�)
�x������w��X:Ή��t����s*?1C�w��~�d͢�dM]�A�
.L�s�!����ާ�4�w����`c�ֶ˻&��LxN�ǃ���H�H|z��G&x	���2v�"�VUzgS^�N7VA��0��~�Or�B��ʕ<�Ա��R�`F����F��kI;������T��ޤd�^n�����#X�w�����G[�XS6�LTIT����g�&��I5���C��4���;�q�U��R�ؤ�za�k��Kv����ƻ���ʭHN.�v�^�겮�U�R��>��2����٘y�5T��+D��Y�VJT5Z��?+GP�L�i ��mq�N�)o�g!�Ea`)]��q<1���>)�"�z8���y���(O�j,P��m����=�{L��b&ѿ�B��7S�ex���B���gɟ��?K���W{/��3��J�OCm)ˋ���}?����O|������
���P���z|*
L�ͣ����g��Dᳺsv��4��j��C��q�#R�&7�c�.��y��kB����D9�z���}	�(P�8�<q�����3\N������F�(��)��E�L���D��&�8竕�{���8<�n7��|�/���)$�-�l�#�B̊�_�s�c���s �iIe
�Lm���PN�L"���/]�*���5�hb�N���=OI	�IAbB�vl��T/�{YVo��ߘ������rT��G�iNx@����0+A �z�C�q�^���i�	�QeC���r����M~�aM�Y�ɳ�2�t�2>B��1��\o@ڶ�6[��sO)�Pk!�^z�g���~���}^2}[�/�ō��\r	��)������Ǟ䎤z��Z�G�uV聻�#j�Ms��$^�+�7E9�+ϲ����Ā�r������	b�Hb���[�AIM��}P�γ����`��Q��R��S��8~��t����K`M���ݲ�]�:�Ko�m����;kp#�t�R!�5ڈ�nA��SKl�G+*�y��ͅc]�+D�&[jꛅwύ��0����Wr�J-���ޅ���� ���z�o@��l�K`� �b?�ib��qPRf�������O�� =~�3�Á�����bs��Gxpٍ>�h�ϭ�l��p幎g�9q<� d�sVym��r��f4��y��}'3Y�z���i�B�D��.I��JJs��L�Q�r�	`�|ZO@�SOKc�Ix̞�zC���lZ*�r����Q�%ƴ�����̄��dFr1��	z\�έ2(vq÷W2�hh��"GB�"��s���ѿ3�l~�;v����Hn氁�:�Ї�4������Zu*��;���& �n��R,�i��D��a����(c��6��߹n���|���?,z�˻(W�
^�&��;��nu"��Y�>��GKZ�c�j뵡c6����3����f�N�\M�InW��%F�.DUj� ����T�V��)s�(�
cӤhu��\�,-A�ã�V�E����G(�9U������	>#��v��1Il)���|�4?��:1X*�9R�T?b��>c�?�� ��%P\A.R��1���f4��.DA�ї߯�Mw��H����T�W�2R�/�1 ���q����K�e*%�?�`����%%Tw6������b"=�+X҆�x�sE5ʞ���&;�������%R�x�U)�)�6� �D�#�z`��?T�AM5����t*����GPx���<mrk�x�j>D���v0jP��AF��7L����Y��)^)<�h�v��Tl��.��2�syn'���R���O$,�v������QڥMT�۩��P=�EI�����R3G`�&VW���n���̛�<���2#�2�j�$�l�ɦ{�0u�I	�*�aq�9�e�_��&b��H	 �?��������(ޡ��-��$w���L�rc���D�<�R�/<���IS�,o�7��d7Oa�%��M��xR��^�18�5N��s��C���{XS��Ɇ��W����C�w�v��dQ\S7{�!w ����k0��2ond���
�gޚH�s�-au��D���LqRL�B��2���u�4��O�/w_���8z�
������L�m�aMa�Wt.�9(���C���+�jżbuB�#8S_�γ`��RDO��\�΁(I�����6��dI�q��Y�C������dY� �u��o���ţc�&BL{E s���=>�I�II�N'��VT�(��;�ʃ�5���]��J�dD������� #v����b�ԃ�@�hEi��k��#k�Q�z�o�Q��H5pj�W�SƟ��ḱ�lځ�]Œ�F;��;	�&�1�,�Uq����?�]}��fU��n��;ƛ�L/	s�Ể���v���.f8d�����>OF�G��C�s"��I	�Y�7A�Jb3�.��s�=y�?�ֆ�J��g���^!��I�T��vi�ʅ��p��΂�Co����4!��b��i<���%Qê���}�{�d�p����PR@�.dRq��Cn�����\Q�u�z;o��%6w��0'=��^����&�JX���]�{�����q�٣��F��OC��+ tt*@�}�3
f}�B��]�;7�}��$���/�A@��b��xBF�G��zPad�n|�,�lS<t(��}4nj���a��=g��rR&���������7ki#�>��l ����~	گ�������+JlJIf����$c(������0]b;>���B放=�s���~��f �c���(�#V*�L��J��޴ n���w!�s�a|Z�U`9B�C�? o�HL�)�AXӦ�QL�o$� �_���`u�%��8���B��(s�o4QȵR�$�"��(ZYo\�q�$�v�Y�ְ�N,y.�7~�P{��%��zU;q�3���v2yﳧ��%�'��O B��	�7�ʷ���2���v���#�g�d�Л.��/;{��G0\b9���O|s���/>�Nz���}\e�û��鏶�5F�ߥ��+0�'�b���XD��L���0d����PB���Ni?���g����E���$��g�2�t��� ���8Y_��?h�QUkv�h�0���J�IF�?I��+ n]�����p�ᓱ[Q�� B���.�&ӕ6PV�PRluW�-�K
Θ�����*���%���S�v[�d3Q)-�l}����7 d� 1]jՒg��	S3�����ΗC%�,b&Gv&u�:߬� �vRÆ�!ZV�r�U���C
C��|�5�~�y"�ix�J����r�C�
�Ƨ��C��SY�[B��Ԥ�s�J���~����Q��%vo�	�(b�+���0��`~��7Y+9kp��� k�D�5�����5,8�iz+�ǳ@�����(�m�>]l�q�^�C<��ܐ_�����5�N�B��&
�!H�p�J��a���\v_��5��7�a���,3�R�Dp)�ؽ�Hݮkۨ,=��ݫ��Op��2N^õ��[��Z�f��9w�U��ì��<;����P%=��G~h�2��9�W|cp�b���X�Rߟ�x�)C�b�w99\�#[�S@�Z��E���j\9I��`�NP�U T�~�CΎ���䁼T�e��L0^;�L
�E�Ќ�5}f�G���/�*%�D3� 潣�����9�F%�q��e��vm$ �f
'��s�Wh���Q�n ��i]syvB@H��O�E���%*	���I
���D���@���!F%]37�EW9����Ln���'��6���i���^(BQ5�omI����E��4�U�{��%)]�/���RջM�hh�4�8?o�o���UMJ\�R��Nn�S1�����aF-2�D���	 	p^�ը�'7l�4��cU!�w<�U�� �����Z��/WD�T/�&����#ضHY��_�﹒��rAk��Ko�����	y��m2�^Ǉ�].�$�yu���}��X�#�/TН�g����,������qc' �^KW=7�LxƯvǂ�p�|�kvP~Oz.�Ĉϖ��l���_��B�r0"�`�2��g����1�-iCo��ּLzҩF�>��k$��W~��./ �q��(Ix�D��� � S�\^�ˋ��>�n�/v���I$��JY$�١8��rU�&�p�G!�/l9���[��6����sJ�nc  ��ڃ	YD,������gH	�tHb��\,�h[��i��?�>��0�
%�
evO=o�Y���J�>(�̴����y&�/���sq֓/lL
e]r�.��§�ܤ�$��I>!��ۂR�Y(�������j:�)�v0M&	�t'��A@Jt�<�˝5�c�f"��w�.R��<5���Q�����D�ՠc܈�؃B��Y�k�JX�����E �"ו�y+<9uĶ� ���|_�@�T�|_�߭s`�gwf�N�9�6��/*�"ׄV�� 0w��=�F�p1O�䋑cD�7C�?KQ�@^��KJ�)����.�9��-`��5xU$
|�ڇ��,&?����٨l�"�*�p�OVdO��ǃ��|>	�m�ߕ!�����Ɉ��W��rƬI3Ԕ�r��lR�͘x�Z����A36l�F[�cko��Q�����YgC�:8�&Hh͎Iwi��@�"�]0Ʒj�L���ȋ�����z�L�|$�#޻%����$����,j�yW�`*(W�S���_��|ڄ{�$��׼`����z�:�0_�x�,`�J�6�^�N����C���E����:��"+��^����삉�]���F��G�߬\�	%2;b ޥnA����l��8Q{�A��5�jp��zS؆�q}��;,���4�B�X�$�ycT�f䃞�3c,����F�:��yT@z�~AjnU�j�ǩ���ĩ��	���=\��ԣ$���f��2$�<pA(x3����ǯ,.�a��$��HFRu��X�l��<��mL�@�X�XyO�I�>l��������w�
�_]���틦�V5�{�CA�y��<c�����#29����c*�����@I����T�\�0k��_}�Z�l���/ض��8
'��f;5��^+P:��@�ܺi�#�ؠ�י�B���B�M�+�i �k���+m���.΅��.9���o�;:6E����N�����-�y�-�S|������("+�7n:�X3�7�4�a[���*Ԧ��k�T�1������w$�f�) c��t��>��h�|�&6ȐpAЋk�\��j�2�r�����7Ecu{��%�^�\��}֚��0�Z��)H�.�5�6RP�n,�B`&�>�z������븙��@�ר�u�	���D�ұG���{�D)��<�t(���k�p��CѨ������Ǫ�e�_��#l�ZƼ!�c~r`?C&��vfPNޒ\��@Y�C���;/��w3V9�K�4���7�Z�}̿�[���r~�J��
�i� n�ڗ�JB����5�1S�K�Z�;�@����"�F����|iQh'�go�I���8�����[�]4��a��%�J�+#Zf"<���+�Y�G�W�gQ+�W����|E���\��R�.�%��N���S�cl��;a����������|t�#�!o3F	���*(
��rg��PmG��w����؁Yډ(Φ�yZ��Y5��*���əa�nW����^���������c@�����ڪZ,�;�CQ�M0��A�=�}4���e��ϛ+��7r1
L]6>�㾣��W���O�@Њa������E�C�LꈣHp$�в�z=U�Z�л8�Z~���vF��]�Uz(S�����<8nU��_�tp��wE,����>=�V��7 ���-I������V��]�&�� ��e��+��O�B�@� A�q�L��,Ơ_�!Q���2JvՑ(�
���Ǡ��QW���|��ª�y�r��h~y���S��6TN1�t�\a��\��#F,M��Ҙ>X���w�r���B"*nSu��[�bw{9��@��>���1�؞�z�>�� o����������gS�&��� �+�
Q%��ڱQ�D,/Uz� j�w����*��n[��&Grj����n��@F?.:��u��� ݣ�V$a�L=9�;2Ħ�o� ���JktT�p��e8��6s_��=Ey�I�ѩQƑVe�}��iW9'�`P���T��f�� IX	6��^��j�����F)V��u�o��	\��!iq(��)���9qb�>���
���d}s"�����Z�Pr,����w��o����8���:��Z��R����_I<��o��u�c8������Cr7D�_>�����[6��ozK|��B����X��0�,���H#���E�c���u����N����J[�8�GۚW��A��L�Y� ���M	�.7-���zk����z�)�L�.T?:�bNۛI��q�H8ued�h1^������)b43�u���v�/���2����������J;��U�.'~��XfӦT0g0��#Q��g$�-�t�N�#�D�&�֕9�7�@��֮� N�=�ɂ]] ��H}�3\H$�V�iӕ��5~����m>����>K�w����
F`ym�q�V��& O�W����,�G'�W"�,���w����_Pz|@��s%�=��\���:z�X�j=�tB�����f��*�RrԢQU���wz��q>�q�ޘ��>���/�W��|3��mp�ܟ� }R���{>9�S-��*�8���V;��M��)�옂�pw>���b�$��Q�0���bX�J�Y���u�s�������{��e�u�%3w�,4��Vح׊���k��3m���A��p;�2i;���E֧b�j���^�ͬ7�?O�`b&�#V!"Q���zf2�#I�dQ�+��#���Vjvt��N���^��qs���׺��:�[���Ɖ�[S�r�D���60��s���X�n�"DЃ���A�6�Q�w�I�)&��y1&Kz��� uPKW�Rʚ�ފ]�GzO̲J|�q֛�l�lJCޞ���5��u�#>���}Kw�ǦPzO ����߿��p,^��~k��$��'-2,n�:���B3;�Eٯ4ֈ��[�䖘��U�3.�r���� <���O�r�jdI<o+�f���gn����
��T���J7Ǉ��7F!(@
f���o����Q���+)A�W�%�<~*��L
js�_)����%H�t�O��n]/o�j�B�p��U�j-b(�U*j0��:3���.�|�5�Z�y���r�Xſ=)�ծ_�h}�{E���ה-���BM��0�����1�d�o(�-�p �͆�������-1��� c!�l��ɴ$�_�J�z���z�yM��L�ZWчգD�%��Y�CO#Ws�\/����m*��G�f5����.K$�/��Cޭ�����_�3YJ��t�q8�~u|�w��J���ɈQ������nw<�x=5Z��\��ǣ������� �cd�l
�n�i��d�/� S�w<A��+�E�+�e�ï8���[��o�A[qMP�ެQ�
�d�ƹg@;cV�������߂>��h���WnJ��G����1����'ݢ��������c���m=U�`#b��,`>/�� �����,��sDu�-���c|(���PpE<�sT�Ho)�mˍ�h�d[�{�%����'3�&�B/����;��Ɖ�@�)%�Ds<��[��P���.N��}VJ�@)q��B�|K�V�-as_������h��*0�#�#�l��m��Y��7H��g��T���Ǆ��A��;�L����`�:�ӷg"�������h;u[U�����H+�g*�JZ�s��56,A	yJÊ�ۅ��!��ks�����Au<u�:u�ey��a}�a����o��x~�������:z�����&E��6�~( ���ޔx�.��X~����1�_�+h�)�E�J���?T���c͇�YΟŽ��1_�1�yu�@����B�g&h��Nq(1>!���-l4�$!$�-�`�|^�.���� ��e<l�$T�s3�}�_��[Q��Ѩ8z�+�D�7w6��G*��<M!V˦�L� @���[̇^!��-��b=�֚h�/�h`�lf#���p��4e�[5�r�#��-jjh��������ޚCU,�8��!F�M��]�K�w�F!���U
�KD&��o�Sl�n�%��KƼ����z�Հn$��Y�cTx�aW��=��^�zc��79��?9Ie!<t9�T�$�����h<��U�h:��'�ʣv<�A�8�����[�m]n�)E�Ʉ�3��,lB,�؎Kl�F"R�ǌ��g3N�#�/���ǡ����!|��/P'ίj����M^?�D>2~	�;@Fs�	7W΃�bP�@�?x5�zd���)�+�b�2���翃ct{�6�F�������Lz���AvJ�,[�r'���~W�u�qi#8�0m>���!����xA*LD$����$H@����4���y��ϕP��
��mz@Us2D��ݔ��P�\���W)j�߳�/�ݰ�,��ƃ^����D+0r��1�i	�iC�6.�>+A�=��T�uU�TF\�J���B�+��@��doQ��a=0���l�,R��Z��������D�{�U��$�m���H�fi����A5�jh�4�:�VtE�@
����b�6�Sgm������jXDtVj��/	`5�����f�Ώ�����~���4�p)�p�㐋���b?+�%���#����AO5��NV��ZQ�M�^�̏�;^N*�@��Sz(7��V3�Wv�mq,s�I	x�R�B� �p֡]�ܷ���E&���>���� ��8�\�KǼS2�Q��0��.�1U�fɵ���1��kbɭ_~�:9�����ru�A+	!Q����>D_�w���&�/*�daˡ�n�Oq�~0�|�S�p���7��w�3�S6����v�.�y\+4��rd��,�/�Lם�3}�f�xn�%���?	� � ��_��!FX"	m��o/�������H"���P���+��Љ=�ח�˻N�sG�'Wwَ�kΘ�VݮTfR�������+���X��S�Y�N�^���Z|���cr�1 �F�!����-j�._����th�{�P��`�e}��u�{4�0��hq>��ّ��P�Il*�|eP#����c�����g����+�;�'c3E�(�mo�=sړ�$�v�T�3�&�,1�]8٫E�X+c��������g��ַn��g�U�}�TF���B �,��*$�����K�~� �3_~G>��m>��~�U��O��?�@P�vFM��1oy&�ew����8�M�N�~�-@�1Q���D�S�$�3�}��.g��Q�{R�4�ʡ��ޢ��K>��\��Ӏ�]a;
m��X�M}i�|T+u�]��6�%��uX0?!/S��~NI�g��c�W}+����o&󘗀��Q�Q��x�I_>�.�0��y�����X_ %x�h��}�(D���ؙ�<f�g�q�j���h�`"#�����K��g9�TN� �N<`�o������_1�{>���P�ٕnu4�؏�Pù,����RG�}�fH��%�r��/J�� V�@X*g�qOL��~�IIs>��'���W�#�Yf07�T�s�W��t󉞯�u���	�?�Agkl���D`ƼZ�])��P�JP�n i���S��)?�L��W�\ñpYMS,fz�^�%v>�)�D1�C��ѫ3�p�|Q���x���-��^J�؏%{P��B@	��j�l���t���+�b	�S�J�N鸋����R��D��5��J�o+��۩@ػ�� �>�t���e�8-�mWV�qZh	�;=��W>~�z�hs�`��9P�t[5��̜`�A��2浊f��W ,d��`����%��tQ5r?u3ai);�
�Q�Z�5�>F+�EJ�H��L{G�3�[فU9�-�.�_l^B|�n�$��g��g{d@���l��=h�mڜJ)���mAWrcK�sur+w���3�bLߡ;3s(b��-��fy_>1���4�֒ H#n��r2I���H��H�U"���e��!S�
%K��S�EK	|�B5�d����<�\���Q�2��?��/�v/ZI��=u��� lD1ɝ��H���l��dz3��^�-DCY[����ΔE�z �׽�]��nqHfz�;��qF���5�Q�fOj��t�(P��;>j���L<x�ɡ���\GX[r����ں3F�3����f��it��O4yR����q7A�+���������X�0��*m��v����]4�F(�Ouƃ�t������/YEf������3�_:�_ �>�"���fÆG�Gi����Sx��>��UQ�}�(Ԯ]�,Q�C����`�`���J9�F�p��b%��#�cUӤ��͍(��cW��T3R����F$�!A��#��$�s\R`�6$�J0�9��:��?�SG"*�ri�����ۡn�	*���GBES�#���E�Z�7m%��d��ww9���z|JQ��MR��q<�J9����N�H�]���4ۚ����kW���P�O=c��̓[�$�F�;��oT���ծ�Տk ��Ȥ�r)�A毋�Xg%^@�Y\�n�y�"e/~�ZL�����B11���B�@�X�e��/�� ��m�?�FQk�
%�%#�3q�'�TL�������0�[�|�m�g_�LF�>�[y���|$�����jjOW� ��x���p�k���V�`�x�5�q�E��r�4���£����`�v�j��Z�d�YL�]�3�h��dxx]bʰ���x�����C�9:���ʓt��o�d����O677�C�!9�6��f'�3z�}�*r��eu�o�NPu�O�>"���x�-;���IjS)��%����K�u�-Ws5xɦp�����K��,�	H�9��xH�	�Rb�`-�"��g���y�
��a����L]�m�*X�oǝ�w>^����V�U?���ܮW��
��[�A�V
DPԷ��B¿Е���*	L-=
@`���F2�h��B��:O�v�\��!��RS�f45�X���ņ�Z�ϰ-�4T�(�\y�GAG��6
橠�T,.$$�^У��g�Q�Z�&� jM��v"kLr��|EL%���As�5��'� ���˺:�3�Ayx�ҧ� �p�d�>81͋%�/�B�<	6l�4�ζb�U?-N��=>98����Q��{O��$u�RȽ,��ym�&;�.w�k��{YM��1y��� ����ޠ΍��J�[ �6�������6�p�����#��+�Ʋ�'͑~�4��ћ	Q�$#i�ŖT����Q��)��u.���#�In���\ots�����M+���h���|�(���2wi<|���`�D�Y=�P_BBT�]p�Y��B�q�k�lKm�d>�n��������}��l���!�Ov>�����9;Z��|�K��O�	�����(�e����@�l)�ڣ;�  �%��Jg�b;k1E����c@I; v &:]t�r�/�R���Df4v#<c��Yd���`��5��h;WJY��kB���'�I��o�$?�ޢ�]G�Õ:����m34�G�q#Z�:��V����*Ny��?l�讗�Õ#�����r=�!*B�0�)%F��������6���>m�W��&|�Q�h�܂�W<��*b����"�9��%�z@@I���8F0���,z%k��)��Zmь��� �[~"g�n���(IB�F�5��l��B`��Ǒ�Q}�-'���������\���5�� O{�}�.�c۰R�T����3��}0�ݔi�¦�΁�qx�A�ٜ]n)�A��h)N_��z��������K������w��`>ހ��ϝ��[���sriNY�m.1��j'�lי�+8�c�L�D� Km�v�~��G��&bQ��Z�ϰ�Jv��.�m'[1uڸK�$�f>x6�D(t��4����z�����R�+�/~�Dd����X��Q�g.�����C��̓����
yە�a��/���L���7�>�g"�4f��FX�F(��{�IC��(�{dj��XlL���)�YO=F)@��`��4x>�u�ʛ���=��$mMD�^sQE+��⯝u��N�)�V�d�"�;S�Ŗ��>y���+�δ��;X�ŉ�GQ�P�r�p\�J���v́���:�N9���xw�fXYw�MȠ��2�L��l8'mҗ�~��$�^Z:�XN�ߔR��L�ơE4b3^�)�N⎉����]/����)��^%ʜ[�źw�koⲇUV~l׍Z�w�d6~q��]֤�Q�r,��f+7;\]V�z�w��Y�޾,�Ai�_�� �{B�8��A�������G\�|���i;
C�ṩ#n>�b�>�P/h�ͣ�Kw�ք���}|��ۢx؈������S\��m΃��A��-�},fne�ag"O"q�H��B����X�lmd�N$���r���wwq���!�����Nmp�l󇦹[��d�r��"��dv
2+2�P�8�S\���%ϩo;5�[9E#�%`���UC�ǜ�*V�����4U��"�Z��H	*��;�]K��O_ �v���^�Ki���/���*���̥�o�Ɖ���bf�b2�5JU��˰��W f(g��������/Z�h��j�._�i��?f�}���ؖ6°�ϩ7D�Ⱥ*��5��(�_jf~A�SL���)|�Wj'���΄�M_`�{X�4���@�_�:��͜Oʤ��qQ��s�!��]l(��J@��O<���9-��sVk?{�hN���d}�%x_#�@0/�+���؋�����Z@J��W���ҍݏ�^�>O�ǔ�M���J�-�J[Z)˼Q�1��s�=��f�O���v1A�N<7d��.��.j��=p�Ƅ+���A��I^��ģ{��}���
9G����~����# f�����]�W�Nˊda��i=SC�N�ؾt9����z�7�l%����Z�e��8�t
�ӼR즗�n��!X$h[��f�<�Ii0=� ���NtgV�[��$��ě�C���:�����	k*����$������+,	k(�B�ӻ�$������i��\�k~&���N�0[����̋��k\Eb1�[T��S�=�n��ҏ�av�����A�P�5f�W����TI��d��zy��WR��f{�ϟp��G�}�ًK�ѡ]%�M�y�˲�)��ب }r�����5�Us��FT���J�3S���Re�O���Gc��m�\0����Ǫ�_����s9<�$�]�?}Y��}^ ���m��C���q�#����;�]ь��k�N|������Fi�˾n��\�=7���8#H�(�ԄB2�b����Fox�N���PnҢwݲ��� ����ې��B=�b�r�H)zp@�y����4u0�Ga�f;�/д��<���b]����н�Ǩ$���1"~�����S���@��6�M�;Bd� *?�����3�m��Vd�'-T>i�D��BA�����-��Ea׫�,��L����PC�]�f�f��x�E9�=�H ����S��ω3�At����d	�t7��v�1��sR���#(�l�^��ir	�����E���AᎴ[�'+���&�s!�����[oO�,��̙i.:��o0bu: �^�p
��~s� ��7D�ŦK�9��\�����y�p�Q^�{�9�- �>� �2�Q�rt(��c�vI�le�ȑJ��-7>���*vh���X J�Y�'(�e�n�	u�d����.����NoJ��-Ż���FҌR8nV �<��Z��'8g/-F�UrE99�!��d��ő�����s��`�s�{��1��U��+�rSݰ��R�ؘr�r�/A�^ݽq��R,҄���i-F�)^�
��\��-]�L/@��eD�S�AI�212Nr1�L�H<0����� ��~�Ju7D���wUK⩃��n��q6�k���᫉+ۦ\'�N.='x������%���k��b"�2�ư�B#+12�[���)������%k���\�ə�-#����ޯ6��Y�d����k�����y'��7���K��}69� �9���D�����%+�����	n��]�'45q����|fГ�{�D;-��B6�"CUj/�Ɩ�� Op"洐�Ӝ��p�H�2�1S��y����/�7A����[%�b"��`���k���C��}$�hր��1W�:�~ˣ(�ِz�v�S����D1�1�)���y�PQ���
�s�k�������N;��SX���2�FX��n�$p���Tj}�5��"H��⇴=|�)2F��"I0�
�����+Hzy {iX�0��W�zt:���%��tݙ�1t\r��ee}����7��DJ�i~EN�������S
�>��?T]��$�9�q�th nW3�k<�(�ɝ�۷�;g�B}�s'�<�,��"U�]bЊ�&��o�5{BV��5ͅ�\_�����;]&�(׿d0z�'=�l�T�l������6h��r�)�^A=f�[�f.=H�����M�a���~!:�w!��s<�1�m�<,,��i@�Ȕ+�Sa�
O�Z�>+獮d}&r�v�;�@p��)���q;	0QZ�3+R���^���=C�ʖ?�,P*Ѹ��tk�u+�gk���(�����+�bt�@y9I���
��[B`\��H�ޛ�ӈ]��%�4v����ͦ�$��BܮX��X-�-�gۿ�6����ʋ��������%��ʡJ�9��m�5������o�B��A�?�����heK��Me:,=L)����K�c7^��TX�R;�;�x|v�q�Eށ�R��FIK.�H���Q�l��=�q��Y�CBE�Zx-cmn
��!�l�J%�"�q��M��4PQD��������hM�x�F����ƺS��j�J��虣RA�1U���>4�0���p��7E�m�&��zG�E|pSl��:\���<��d/�n��t�������M,(<.�����tH}�g�\l�c���q��7c�:]�I!����Lʜ���ob�f�@a� 8�B�;��:�%a���	�4�+�U��A���?14:��ɦ����Lt�v�	�^9��i��4 J���ze����D)�6k1�{��=N�F9��, �|�魾�Τ2"*�	�Fg�j�z� ����z�$��W�nFC5��L���1��� �-���
�Q
)�ֽlI+��y� ��*����!־�����p(^0
�/L���m<8�V&4%:���ti�l����jV�8���5��4���%''|�A̤p�פO�B�Ǩ+��P��{4*ǔ���O,��0�ԫ��qsS��\�J�so�]'��KH����0RJ{�񔢇R�[Y|2t�^�QMQ l��o�ˀ�Xc��)������یҼ�^���1�k�]W4p^��`G��)!Ő[n9�,�zC�v�[��aY��q�3�o���o�R�j n���M|i����U�|��~B��p}�Z�*3-��������淖��R"�q
�?�Swn� T#���sg�f�;p����	y�W�&n��?~��^$+�e�������j�eH���`]V �>ᕹ[�����|?4I��$���Y,d~���D�y���l�1JQ=_.у�h3<��r�<\IH�hކ#��c]�)�*���y,��+�Ǫl�6'�>��Tcx�n��1H?�IŰ:��&����;JngR��KW�"џ�9!n��zOs�ױ���x,<��#�p4�ܕ��{�X���sʛ�����yH��Ff�ek薴��쿟��'�kc1���&h\r�?^i�.��D�>FD�����(�{��ǀ���XX��VíJig��3�m���:%zvM�-ߊP�`\�~G�k[�<V��)���o�T���s	�ܴ�_�=��L�=�7'�j�ލ%T������ڽf90c���_u�'6ԥ�{�����w�(����$|wG;=3O�q�,�j^Z�+^���Ǖl�� |��:���5�8I	���s@~GJ�GRZ���u�E�|�Yhl���hԼ��R5�5n��.D(�P�|�O�ws��\�q���f�ݢ��W�I��*6������S�{] �������v�ߖV����w�?)�-�$=��bpmK��FG�%Jw���u�Õ~�k��n$�HHv#"���%EH�DM�D�:�`��J�`�`	c�ݨѢ�2F�1�э�we#�����=��������+�nXFM�{�/��������}�o�������C�yA%��GE����cw"��v侱d݄8�h�P�������j� ���U	��md0/YRm��{N��)��X��}�3�a���F�|
�El�#��X�7%}D�q��|1�g�h����h&΍f8e��M��Y��l��Gi�����Mux���(��Tg�ldFa<]fֆMfG
S���qVU��n��������ڭ�HHeN2���^���. �j�g�����5|���뗣/%]�W�TXfL��Kxkk�Ȣ�.���'{���ax�:�"l����U���}Va%�'���?R�ֶj�����]���y�zBkM~����oxj1Io�����������]U�p������19�Z�4��#\���K���:��-��xT��+yN��$*�[J�`��	�7܏��v��<��_��y��j\����-ZI0���>d��M[v��q����g6��`<#�p�y����-
<��8�&�b{��j�:�&�^�B�aG�B�|v]�Kk��6�'r~����c��B��q���	��J�/���'Yy������nޏ���~׬��U��#���v]<��a�7V�Ic���Z@n�=����M��ٺQ����_���}��Qb���O��>����`p{�l�L�>��!dDbϪ��Oq��,ny辅a�1ξ"����N���e���⁃��H���:+�H���m����� *Mp9~�d�1�[L��l����A��ܷ!/�0?M��EÉ^��X��7Ğ���=�$h�������<Vۑ{S`(��f<��SmhOE�UGm
���B���ޑ�E�}תǃ9�@(��W�k�ϓĹ�k�!�zÎ\s~�J=��i!'A��^�śs������U���H7�:Dʧ���;��_�z`m�F�#����F|B��w�,�|,��������/��@�ÐW���n������߼8zݫ��@��6�"U��L֚#�W�gX�L"����9F�0��4��Uބ�U����8q9���'"u�X=F;����6ܿC�]��=rZ�Ao�|��G��Q���nU�@����'�D:q��؂��J�v���eCb̃�K�K��a.�P���;\���63Sf9#�����&��ƶe�9r?��q������	�0��ߧs{v߯~R���*�:�5���LE��K�>k���K/\~ED���l,�.��֛
��>p^]�"KM�
����&`V��p��N�$�Z;����Ǧ4�SI ��<.�3��RK����~2�,g������K�ǛP�����u|��������T��CL��s�t�ov�)9�n�L=�2���w���������@��/��?�k�0�ײ���C_^��#"�g�C!�J�XF�I8�CY?Ս�k9����>v�k����ddT��U�IRW�_;*�l"[	
��]5;�uo�vg�S������Eƌ�a��[?N�_Xy���cKrսȦoaKYCl��TO⾠"M����$���8xD�_w͍@��݄���&o��׵�e�Ҕ��=�ڪ�4%x Um�q��c��1@LcYKXY,��)����r�h�7�u&��v����W-�lM��i�`�#k|��5�3?�=S�ЈwĎs����V,e�� u/G��So"g��1��8�Y}Ǖ���|3*<0;��7��/R~M/�}�B�li�Q6\���x�FY	L�B���צL/� ��xk
��<���g�[溫���<�^��RF���%3��g�6ƫ��B5�ii�w���'!Xz+�q��v�ɶ����F��*��y����Dk���َ4�V:r�&�Z���x�C���vDv��h:��:	�ّ_�A��
>;yo�S����&5�Wڵ���zK=��h��י�Ё
x����&cNk5��?��P�� Q��ml("��Gv9L�:1-R��e� �ox~�S��4�՝zDoGt�n,}���ُ8<��<!�w4�*�����LNO�ֻ�5����f�d�%�N0�֤�IJ�(��S�刴�H�v���q6�Z���p6�92u��5Zu���Y|�o��}�=9g޿�}�ŋT�o,��?Eo��!�*�:�P�y����
]7�9���:��K�l���8�1����yaWF�òǨ^���`i���=�6���WC�=B/����\|��%e��Ry�k��	��B�fd��V������`w�Mu0���$�/�>J͵L�/��Ȉ�z�����Rԩ�	
�w��r�*�9$=3���sv�S�4XxqO'�^/	��Y������0;(�X)�A��T�j�D��߿�!����������R��@���b&�k$3I&7]K�J�A;����ʝW�E��S������(�k��b�GE����P�OS�1uKfJ��V�j� \3���5ͣ5}�\�	�='��3�:xsY��Y��A�a��^k�{�x�&~䎽�mɅ���Ye�_xj&�Ii]���c�G5�^b1�|��R	HW��� ��=o��?� ߬��жk��;�ܱ�D��zaնnb��u��i��8/c#'xnq�t@-[�0�[+f�Y��/���t��7����{���C���+�f�f�W�{��h�UsUi2]�Z�KҖS�X�����u�^�jȊV�0��xT,WⵁQ:ު۵"�q�M/�����q�"E���Z~�I�O�cuܟ;#m��="�|e���#�����V�e3�е�}�-?��č�|w��|�+�@7�gd'+��jΟe��A�~)�{��Z~b�\�|�`$?!��+����釟R�F���Z�ܵ�&��9pĀ.���HY�J�Ʀ�k%�D���)F#�LY�׬�+��xpj8=���?�fzUL���]����!�[�v�z�l��l
gj��k�R�m�K��7T�1����>��ݽU����vUt�:�h��N�Ĺ��N��{���N���ȩd�i?@�gIf��m-����.�j���K�T��H�9n������R�`k7�}\c1�)�E���*MڎP\�%Q�U��K?;�u�b��_L|�>�U'.�UO$��n��٦/�q�3|�=̧#VsDU3�7l{�8:�ؿ+\�"�����K�+�Ⱥ�'��%,��v��_w�Vl��#���_?ց��+D�⎆�w�tʯ�_.�-ߒK�i�{ /X�W�����!E�7w��V-��;P�*[Lt���n��7S�cC��� ø��J3gj�����"�����Ŗ9���e��.H�Oi������5�n���by�ӧ��N���v8�����1���MF@�m�"8W�[#'����.(>l��Z�y�����ܹ��P�@e9��-���_H� ��Or�4�g	S�J��L]_�6#ۇo4���f��p�e�LlqR�7N��ܫ��]ܪ�(4Pl/4@)LQ�N7��(��LRUو��o�l�화Mpl�x~d'�|����[���c4��ʮV��	����)�r���`\���h	.(g�E��D�2à�!%�m��:�*�	M�3������� X6�W�7V� ���E}	����˥��L�9De�2��P~�|�iX���Z�f/�uu0�&����n��n�'4��-�~�`���WYEb��s�j���㕠䟦}��҃����_:#k�r'h,� X{�]%HeJ���׊,����
�a���Bq��Q�� ��ٲ��3���9t�џo��1�[���R.�������5��J�5A`����a���H���g�T՗-ɥ��VQc�%�qw	��Eg��G��h`��W�7���+�����,K�������P)*�ՠs�����H����dpk$t�1����+,*��3��ݜpM�)I�:��/�`�pA��:�~ä��5�`T����̣�a��ոx<�w��V���A���1ǲ���:8Ҋz�p���f^Zg~'��ze�Q~������{��O��
!%�Y-xK���TT�+����48���2�n֩u�]O�3��Y;�lo���dg���];M�h#�fG�J�uX�����.<8�������r�zxS�d�!��͉\�wm����2Q}��!���#m�U�g�?�H�#߄��1Eȡ �to)F���`���.��XX�[�����x����6��j�����9���V%�}��0z�`���^�;�T�ϼ[�d���})���5��V��Z'3M'�j��G׺I��]UYN0��!�QS4�Y��i9�5J����J�[؊�[��?t�����쀞�x������A`B�<K>!*K0��,
�J��B�_E݌|��Vi��s�^E/W}��t�����zE?���>�SoG�1�F�q�u���� RN���֬,䦍��ܧ������0���B��\N�L-�����/��E9�`.#���_.�Q��0�rԝ�F?j��!fw����2"��p�K�\v����f�uR��k�yz�9��0u��ꤲu����5M)N³�~7pF�,�T�O��_1t��������H����"�+R�kC�;QxzY�6K�JG��B&�����7�jb���~	��hw=L��0�������HC�<�^s���Hz���9�B�<b(`��@O���]w��M/
	�eO����g�!J��wͽ9Y�PA��r�a^֟ld���Љ�/��_�2,[ZZ�G�fe�bn~�A�G����WeM��z��ˉ��f��C�)?����Z�H�8xF��DF�������Ԃ�����~�������
*�1�z�?K|�G�<v�Jw�^�.|��)>2VRRY��Ur�L�4�Ws��ve@��'cZ.��u���uM�#a��u���������\��-�ܟ��u&kE%��}���e)ƥ˵�
�c�r���Nin������S�t19�����%����̹]��\�GS��&�K���>9���*�+L|<L{m���^Vm��hq�����)�.i�\��YH7�^r�ni�����`�03�n�Cj$&���2_J�<z|�)I[7'.9�4�T���P
������g�=Ԣ�ov6i�g�w�]z����{s��l��<#{|8��eޮ8�zA�#�n�|r|�|���J���Q1���_�W�+,���U:���X7Z�V�ʭ_��=���`*�e?�u��0 ��XZӈ���&�-k����Ѧ0�6��5C)`��g�KL��a{��H!㟵�^fwv����+�?�����t�zr7%�ȩw�:fd�e�;ZM�DP��G�g���J���I�M�O4S]���Ԋ�6F��C��V��nA�a���ъ���KB����� �Q�>qw6b����E1�?4GvA�n��%�(|O�]�ģ���<\�o��������ώ[RoB�$�[���O{,�ā��5]�$���X���n����0��7�+HY����֛ Ɗ��!E{��1��nZ8�7.zc��xc�j�C=�����o���kȓ.7�A�l%�O\+�4`~��x�b���Q�m2�ܧOc���8yFm��4V&�����dȧKC�K]��[�L1U+Nh�:m�G��5�����(�O�3�L%m����Yn��F�k��y�Nˑ'�B�c6:�K��@f>�5�ԋC�(�fȟ�윽�㠈#0d���_�ũ���Vs,B]�����{[=)!V�R�=��?#�� z�F�u@�梈eFY��T!�Jxa�
��?�_c{0.h��X�%}��zۍ�H��H��cz�����Ig��Vd}}�f>�Q�� �[��6~�r�$0C��L�Pc��:%\�[�t=�'�%=�C�OQ�ȇ�[O�~=TO"t3�t2�z����md�K�$�l3ss�����1Z,���w~[�I\de"l�9�~v�k��sh9u�9�}dQ�S�,���������vM���s�u:��No"=����d� ��zR��M���Yr�W�rn8�]�n�DE��2c�#c}^E�N/5��2��P����ѳ����-8 ʺ�J��<k�����LA�J�܌�-�	\�Z�⦱f��X����y{�;��]��Y��ф��ɬ�4�l�L-m=]�T:qq?>% ��h!&M����[��ƕ��,VPƮc�K,���6�p����]�����~�������I����,I^�^=8��R���h�ڋ���pDR	:CBt���1����:l��O��u F�P��g���)/G
P9Gڏ_L�
G�
h�$�$�$w��I�!�5������/�����Ab�Z~��gޙ�9�*��k��ݟ��lϝuQ͋T���Y���#��LUo�X~�u/��6�0DoW6�����2�V���0�ԁϷ�y�m�KS�ő�1�A=�}�iu�%4<���&�B.�(�J}�)_�E��#����fu�O�w��\^-l��Z�s׷��S��e0�=�mc��Wa�Xy�$А;�ɶ-2�����2�t9&��WI�;�EýL��RǙ�cɀ���D0���tb�4�X)WCE�׵k��eK��
��1F��l,/4���Dx�d�w0?˝;zrЉ��e��;o�Y�8���b�y���y��nNo�7PN��r]�,��Ʀr�c)E1R�}}p5銔4��/��|���4H��i��@�C��od- 1�j�����ɉ��K���S���i�����3"��������
Z�1��WĄ!c0�8?s�:%�E&�����y�g�891f���m����|4��z���{z�L��o.�����ګo|8,�z�Xa��X<e?�n�����2�H�-ڒ��m21ϻ ��F��n�&�)��vmƈ�Oy����I�q��20���D��r����q��C�����ȃ����on�*�8i��nt�
�.7Ʋξ�|Ӕ����z�i\�}�=g��X�m�� ��Э01�0�y���.�g�@j����?m������G��Ob���t�Z�ٔ�k��*���L<'6��N�5�R�R�� &=�����;��W?�>�W�ȥ��Z=<�x�'��V\��F+��/cHi����.�zC�]P���ts��b�=��h���v�{���>.�cUY�`S��)���𵦈l��U��:��չ��m�.�>Z�ϗ���`�D��B$��Ӌ8Io�U�>܈��S(0�?��Ǆ�C�{�n�������O�ќB�@R�QM�q�_��ӝ�����,q+4wV� ���ɷ��s���+bq�5+�;��>�K�j��<�Ai�<k����U^0'�Bz��T6���Z&�	����Ő����Nz�&\�#�\Lxq���>+I�G�J*a��&�����9�+m��#�=���Co���}<�IX�;��,p�@=r?��,�i8S�:�ؚj�=���P���y���׌�7b sH(�=��w�/l�Sj��t��
����-�8l2�.K�ه1/#�~�;L�C-�u��!bOo��S�[|�ƫ��~��6�m̮�[\e$#��?�ʝݩ?�)��
.IP*�󛷪���w��~�#�=��d���YdX���+�߀�zu�5����ZO���f6�������K!����#3ْ�i�%�䘳~u8�Q�x�0���i�3F#rt�o����Y����w�w�Xo�"��=�:���i��K%�&j��j\��Z\��<�Ll���R*�^�rAf�s@P�LY�.ZI?bⵧzH���y��pzh�s�`CO��3t�����̐����^����Tk��	����J�;�Nr��D�u)��+�)M5�?Kԋ���J���br���:YQmG1�qӨ��
ZP��� �ġ�q�C$9��l��B 1J)�^���<>`�]a`h1��v��$ϖ�;�+,���t-�wx4�eጤ_[��z��R�\H_B����~����OD|��̻h�wݏ������n%ُ罡�l���#�-Y�Ҿ���6�y����@%X#׮�umW�AGz��5��� ��,���:Drqg~w�����j(�=�ɤV��s���FTr������M���%_+L����Z�.�����=��[dt�%[�2���-�uc�_�vڳ]���~rևT0P|wɹ����Q>c�rH����"*8˦�8���������V�/����K6��Ee��DnbQ�sȡZ��f��>�"�>�W�SXٽ�(lb�E�����	�<D�nO�H�o�|��y�,=އ�r�>4�����?F�|j7��}ӧ�(e���T���TPZ��Z�2���c�t ���Xx��;�f�Z��x!'pj�����U��푾ƽNN~'%s�id۰R�?��������x%�^c�� 5?~#�ܒ���\�\�+檦�f���F�A6��+��YWɯ��p�UI�&wD�����Я����O���
+<�����}��lp�w��'�m)�/���G�]f��W�{o�\�;9[�M��8R�ٜ�L��8�<��qʖJΧ���1�7�������
�ၢA��QV��"�E���(�0�{���47�fL|��V�M��36g'K��J[=���}R�2ݜj�Z�x�A �)n���]",��9�+�Z�'e&�N�a+&��Rd�WY[$p��\Q<���ܙ�D��9�X֥�z.���_�d�!���F\k�����T.�a���|M������"'��1��M�W�v��0���ĄѺ��Θ<��"ٟ��ԑ�����W0��ƛQ��	��ˇ�\
f������ ,�rV��{o�8]ױV��a�%��v4د��
WVV#�͹* R��)�+�������1�XP�W[c��Y���S����H��p��JQ�\�Ut۶3���+L�k��<u��YwO�b���<�IƇ������b*nr�X�%���SV�{�[��]3��܏��>(�$$,�V��F읝Wj�����wu'_0��:ڏ��>8�����t�;cV5[jT
��V�'K[��D��Z!$����B�3�N��Y���R���7�ݙ�`ܟe��fW�IŰ�v2�+ht��C�zQ�Pi�T[n/b97��������q~��i�Y�5ԃC��aҙ3g��Gh���륝���CyҾ�����7�33ī��C���������ㅓ�[^f�3_�JH�]�ؐ�XE��X�RZ���\�+��<S��r���Q�����	3��N��ݞ�z_���"�FD���-b�@��$Z�6]�^�:���?!H�ڹ��s:�SO��[�}_.�!]�hG�C�~�c�Z�(�S{C2�H�6��=]}X�嚆�G�	%�,�^�X�jо������ A��(2�z�Z�Ҙmh��C�D(Űj�aL�|#E��#z��Ip;�o�S��|��r��8�-[F�G�X6���A�rZ�e�߮�����z>|��^��H�߿��O�)���3-�0�?`�Vkye&�%M\���6��
�6��k�į���x�=v�����p__���9��*�������j��:H��SF/��.On�����Pk�V[cK1����#�����#�ž*9�K=���t�/jy;��A���O��vSM��5�&.M�I���	 �2��Μ=�ԣm�ʆ;_[���~J�/���D?�d��v�Î�"�c���2�sv�6��ۅM�T+!�8�|64(^Ǚ>�_G톬�94W���b&��Rg*-J��r���L��eѓ�x<c)s�^Z � u/C�JN��s�*IC$��T9-"`�EO}g�e�����]`p���7E�J/~}�B
�G��ɝ�Û���Ǎ�V07�=�p��u�=O��u$�է�(i7���a_��N��^&�
pz7����ΌP�W{�[teJ�aapn�뇫����4�����Io10���b˘�c���H�����{K��j�z��<[��A�/�{р����L�-���B�H	N�d}Y �춑����kf�_OBX��Ȟ�[�̊Ǟl���!��=��B��kɩY�jq�^{U�Q��ѳ
�[�CH2�\�1pVBC`ᅅ�a��OM<֜���B�AѾ:j���û:��ߥ���K�#튶�h,M�ݐ󅣑�T�V~��������}~�owV�1������s�J�u�|��G;rC̉�,��5�y�{C�=�������ʛe(�me墬�|��[�&�-��0���
rD���y��G��~*�.��p~���T����S�����=1Ы��!���bO�<B�"�N�ˠ�c��S�V�9C ���,�6.�\��p�Z���g����Q]5b4�����`�c�7�):չ'����gQ�%���O2���W��$���0m'�܃(TQ���B�6W8�����Fh>Ըc�z/}{ �%����A�lvɎmB�[p��uU�7�g%bt+�_�b¾�t�uY�>4Ì��LX���-]���I��K��^���7��W��u���K:�����h�(AY�94��񊼺���djLl"�{�tfsVV�~?6�?f�3*U�{O)(���x$���bO��#����k��������X�GtvV��P�B��yGk�D�~߲|�B������ }���_����sQjF�`&Kπ3�-��^�8�����FphE��h��/�J����S{�,��%D�ܤ���kB��Ƀ���
SW;9ֻ�;��寴9TT��I�o��_�tYqm:T.�h5Z���fFi�"&?J�e�p��-T�#Ӂ���.!��eO�g�@��du�RT��R�lx�2pg9��~�	{9�w�@�m��(Y4�)�@x��	>b���kj�<�4�ؑ��fӀ_���N��aSٳ�zy�qc~#o��Ot�{���9Cw�=Qu�����I���so�	���B�XXX����b�kv���/z�w�F �V�Z&�f.�N�Cm�����D�p���������t�C��S�b���F�R�L���&�lK<SӪu#P7%�({�K��{���հQ#q���G�DK���Q�'K����cem��0y�Ψ���T9+�7w��G���!���.����k8թh�/�0.ðbN�����=�d���N8״�n�If�U���hD�������UU[�;ݝynN˕�y#�YY� ��MEC¸5)A�����GιN��#d�����&���ӝ*��8W�\PNuG�ҭ� "��9z���S@�RN�]�C�Ug��~X�J�*J(�@EOMT�LE⚧���%H���d�����
ۆ=HZ�1E�]�]�0C��Q�۶���{�{����]�Fj��s�O��Op�FL����.<z"���(CQ����M������	�<y��z���eG�V&������U����3���9�Fl ���Z��2�F����n˴��b�&g�Y[Ŷt�KЌ��,5QXb��RX�*/��o�����B����Hlq�Ő+��b3���Ӕ"���S�/�<���8��j)﹝ �F�i���"�=�J��Od��-_�qr��Bj�+�'�֛m��=�
_*��FÅ#�r�UI�uF�0�e�cy��y{�%���z���2+UNx�C�0���"��ď|}x��`u4Uu�K��E������o=�Jrg�>�
�Db��z�j�F�Gi�*(�W����~��C)
��f!]��Ӟ��N�y���)5U�h�,CL)5(�l����el��~�t��7��iA�r�+r\�c���c%�S�]IW���(齂���'�92�I��b��*q̹ᬠ{�x�E`?�kv8���5���X�(�Қ=;�6�Ϧv�`���l%��ڇ���$myףR51!m����������嚢������G�[�҇��Uy��GU��W�]��t<���i�\w�`�gQ�nN0������'?Q��ykd�:q0�h�)*SO&@��M
s�����Qy�E���72����$�<�I�?GZ�e���!9� ĽŖʩ����)��3M�S����j-�n;�]�����N�?Jڮv�Xʹl���S����7��'sAO<ܗ���m?)jt��̝$êJ�b�X���Js����9�:甕�� ��.V�ƛ� �.ͦ<w���z�F�wsc��*��}�,/,�Yֈ�W��>+��Gi��
ڂ���R��6��[��_E�	��*�.��h�Ӣ���S]H�.u�$aKm�ɩڍ��$*K_�^�e-o���TNB���--��S���	3}���5�o6'YT-���^?k\Po���O�v�K�=o��kr�%�����P���ڵ8BbR��nQ/��7����;$��n�Kp�z4G�O�05��u��6.���PbS��l$�N��e����:�h�O�u���ɶ�a訉���ׯh���7S����ϛpȸ���;�B���3D!-���>�.�2��PE+os.�%+�k���^"�����
-[2�o�� 6��yOy ��/�Qfg�L�m�bNt��"���(>z�ra��ϤGk0�ىDo�5� C��Q{���D�|`���,�Ս�i�ٖ���LG�託���E�ԭN�v~�cٖg�$�4�6�3r��Y���n��~^�3��/1�W��Z�m��AN�X�=�v]��'���C0�m}����*���C�����ٌ0�W�yf�c�]�Ț
�j�Z�wj��l�5�.J�R�}J:��6vrp�U��j��m��x�/��!$Υ����x�"�K�����
=u�P6DG�{mx�1*6}{��<�AڼR�'��t<�<�K �c;���
9�;S�n��k�)��O,*Ӎ����
b�^R��F*S�ǩg)̏�甀�b���czy"�y�`�$ur�i?�gy/l��+ÚuK�~J��}��(z��+S$�=�O��y��PHal~�U>�V(�,R�Z���:|�s���?�$ۯ��jٝ1��1�\��n��;qC�:�����j2�Ү�VBrH5Dמ2B�z��⧲�w#d��M%]FJ�DN�Mj����y`"ῆ`*-^0�!$؉�/f��UPݬ�f烐:���}��#k%�rΣ�l��R75��W���Q#Ó"���Y��;�%]^z���2��pCQ/ѧ x��)3\��A�3����e�ۦ��4���Cʲ�qv_�|1�&SsS��0��b�,��×�q���arb"�/����4Xɫ���y��5:jt/N䎝���)���� ��jT���b��c���-Y���௬S*"A�Ҙ���z�`���vY�rg� �Y���,�@lA��v]˚� ��ܐ��Bʺ�O�I����o�������n��\H�+y[	-�"���`��\�X�Y����K��hA����SY��ڶ�a�hh��:~\㥝�����u&K����=��h���Cq����XF��f�:�"Лd�]�;��wN��PY��`)���yR@D�M(l�)����e�WzO���`S12�TubF�4����Z�����C�5/�>����n��%�T=|�J=_} ���q-�*3�\�cS���ȏL�!��37YձJ�8h*���@��{������r�pBj�=�0�dy�
䑂�5^ױJ.W�$�Q¿�.�՜���c|���ʭ1#YU��g�V{A�Ȥ�R�G����Q����4���㙜o�����8��m�����J��]�`�SYU[x���Yth�<��"5UU�ȃ��|sNf��0Iv�E��{!6�~,�vC�ٕ���3�){:aV���U']E]��jN!��X0��rl5&$x)Ŧ^�W5�0��.zǦ�Bk$�{Ȋ����a�����7�/'sf˪ւ
:�mx�gKx�mKf_F���Vb'.��uy�~_�:�ş�� ?s�qI]~�����h�7�z��S�Áf#�A�}E�O�yF"�c҅g�O榺���Ӧ�\�G+@�����&m6�ϊD³j�M���qv�*�+5�������à:=�xl噳U�dS�����3�p���s	������x��P8�ѝt]!��������,�țt�pzP�V�+�S�����T�X�dQ}�����)u����<�D�>���Nq�=k�Қ�Zh5�t)B�srȞ5Ġ�{��jh����}q=�!v�w���#Po�0�DD���$ dp�󼨌�U-i�ht^�c�g�]X�	�<j���:wo�F�O?�����V`�fEF�.G�� �:�����y�E���{6.��X��H��F���gS�R��,�� ]�����g�j���Ǡ޼�?ꙩx��Ti%�K-��X/+������;3��#�?�4ݫ����$]���dm�U�/�ɑ������Y4�Y-=�t�w��hu��u��=ò�{���_6L�X`�ff'�r�t0zv�=B�:�2]�>{�`Z��ٳ&�,��f��ׯkUs�Fvʿ��o��u�w���R�"�|&��ɍ�]��w��s����N*�|G|�$���f&9ի!)*�L
�yO�����f����@��L@�jb"��G��Ɍ��9�/��\�ь����6����5?��6�80����⍟�(��i�w�Hy��>ײ$�H�MB�cy��Pur��?ù��A2EA�#��4.I�\ú7 $p?6�Z=��bvQ�%�h�<F{x���LLؚtoܵ����)�6A�p#Ij.��D��R��踚����ޢ��-��D/J=�}P���������չy^�Rr]�mZ?o'����j����p�~k�w�W\s͈>[V;���AA�Ip
\q�'\����8�	�@]��K�w=�g��V�m1HJkl�������ld+�b��AK�z�����5*�YԸ���QmA1�C ��������yr�H��5)��b�K���%!#��ԉA\Z��G���F��b
��Q�ex�1g�X��&8�����*��;Ǳ�Lѧ#y��2��<����@��Y�m�X���;�U���u>�2�'��=�Y �JW�b���j5-��3%�_�������ݤ��=������y��_�+���GG+1�/���8����l�w��T��\=�u��������.�H:�Cb������k&E�+*�2��ѽ�Ij������;��:�]���D��6����vo���� d���7v�[d��A����z�C �(Rg����d���.�b��Ϡ�^��^��0�W�g��(o6)����a�g�m7A0'{�N��7Fn51���і��<1�il7�{aY_�F����F�H��U�ς9��{��*�y'��a�L�,.��M��bQ���ԙ�5VZi;A�y�CXnk��E�8��^r+��t��2�B��9�����g�۰�#8��^JDpHʵ�����G�=�A|ſ���u�~��T�jM�^�
��i'�j/�FM���&���r2��;���qΕ��ƹ�6�����Sx�4��̽K�+��þ�8\��fԈ�,��$(�}���z/e��bz����{�ǣ�÷BÕ(k��.5t�Qn�&vO���˥��l�� 19~��^�Is�!���d�L/���G$čD(3Yuf�:Q�q�{{x�hH�{�C�� V���M�,ng,�Y�����@��4������`A��m:Ij�o�O���4lA�p1I׭ᘏBO��{������=�1$.+4��,/��x"H���8r�-z�=4j�V�(su�u9
�k�s_@�<+þH�>J\o��\=9��n�"����@�wܙko��>�����0�$U.XN{�}���Y�r��:5p_9�T"�B�xd�F贇a���_?��|{:d!��v���gx[��&��¬� o�ǅr�R��K_	#�Zs���cG�}��VI^q�r5U],�.���~O�V�M�v��8�<�RҚ�,��U>"E�j2W��/�����ž��=0��^y��]����O^j�C?LW���J�ܓ4v?�׼n\y��;F�˗��f5���e�v�DzIk)+C}7u)0��B��<�(��DMp1�7l1u!H���P�R�T�Qm��J���x��m�Q.���eV�a.v�|?��Yu���_�K��Gg#y�(�1�� 6]5�ۢ<�"f�փ�� �Z���E�b��=�O�%��O�dz��pɎ%�(ǮS'��9/f��sp���h��W�l����G! ���@�V����PD�rZ���,�ܭEk��Ζ)g�����ԣ�[�mE��b�(��DãuC?� 2k!2xd�HSt.=��&�,0_XX_��;;�'o^��ѩ�H��m�x�0<k52h�[\g���]$��D�9�J����-��ï��0����A���7��,D1�A�0uQ��lz=�b������o|�O�3BىZ1�}��������S|�f������'XY��K���l�13Gd�͎�b����:�CL�>]0�;H0c"y����o ����0�3	U����|�\݈�hX�b�Ɖqǩ���v���<�%Kvu��7�e8 1)}}���N3����L4@G�x�)f�x�.���&��Lx'?���O��v%���v���n���j.sa��8��%9^0��i���̷��)s2D�M����K�6��Av	q?��?03�HUc���N����
�8q�_�4�p��+WtԸ�#i@n�G��R�tT��_B�ۈZ;Xg��cl�M�UC2���e��ze ���#��fށ�L
x+�ű�-�"v�W�L ���ң�U��`zz��0���v�s�=6�Г���/bKhn�7�y���7��1>������|�߼��������(,n����*�ՓG��(n��+��`�c����Z�O�0�TIJ��2Ug�d:4��OS�[������G�`=�c�9V��E�98������b������B�=�M��gh��?���j�9�����O�{4�u��òʳ+�F]Ai��,�����* �tE��+� zW(]����J�!�� ���f����?�#�3�����s'x���6"�T^�hTf�3s�� �Dǥ��D�7�"a��ʊ����>�ܴ�@?����n#�'M���ʑ�
>&���8�q��>�g�X�U�xLt&On,���~�"�3��1?��:��JY�H���o���w���{��8�+0. �����'��y'XŇM�+F*���(jX��y/�t �K{^z����b��9���E[�	��m#�Ή7�F�\>�9=�g�N�dD�9�J73��VO�Y(��*<��a��<軾E��6����.��p,�t/�4��$�kci���֞[T*e!����dn�\HBFG��Q�Ag�~ǹ��n��q�0��ck�|��GS�w�(��t��]����	�$+�<�ԋ0x���G}<���acU1H� 0NX8�ȼ�/�/��~3�"#C"���'���%�c���W+�u������|�<'lm@^lwL�q�o_�xav��h�X� �İH}�����U���!���Y8�O��E�grV5ñl�6{����Y��x�7�ݻw/�âI�O|H�O=Ji�<�F[�����Ia �<�X��ߟJ���m�"e|E��?ɯ���B�(�"`�NX�
�=e ԀAo��Ei���b�����Y��P�\Z��rh3#Ω��SgU��t��v�K���0�D�d9�~R��s@&�\�5ģ��e�A������h��1� �����i��Ma2�x�R�Y�����j�������ꤵ�ENP�mDhn�x>��k#f�20	��ŀ�T�a��f�1�O��r���� �	#���"��!iFҢ�p��s��]��,�'���`�Ʋ}@b��� �ϹŬ0:U��1~⦞�1[���n�c�rV��le���s��}g'�8]z�<�ωV�zx�?����w�
�k��������Vz�!a孹;�e_}q��Іk]���o�#g��ߡsFѩ���o@�����mF�29J_#�����m_��c<'RoF^�3��S�A�����
�������13�s��?!no�s}m�J��B'8�]����
lU?/�GUL����Ua�]�E��~��nu��C�԰�1@)��gTñh���j�3�}�ƕj�Y���1�
�������/_6��V�X�J_ϗ��H̥+7�S���T �\�t�G6�v���j|~G�낽��ޛ�����.7���=��>z|�>;z"8O�>r�q����ĸ�)Rh'��8�qk��02_��P59I!!�j]�;�̳ɔ'ڠ�Dsl��O	i:��->��ڶ̋3�vV�mi�r����U8�0��"K�3�N�5k��*�{��s��P��N����� �PBM����>H���Sכ�- �a�j��|�Jw�:Dg�ͳ������������wP���މ��b����q��Kac�����@a\�~ �@�W>�0W��[J{������F6���Å蝪��Z�u^_C�<o�$�¡b������0J��mf3��Wx���s�F=XR�qcAװ��
�\�f[�_�g�A^Ѿ:�8CC!�1�!)϶�A��{�o<�+��w�Jp߰�6_��f��=.�Y^������̿)��w�Jq������@:�E^�m�����[��\��^"ް��Ҳr�y�X`l�v��=p�&�_��k����k�!|3~��]�Kl
�����y���\�]o~���wިWA�3f
ȗh��@û�����!��L��h�"n�m]o�K�\z�D'��EAx�"�A��3ޝ�h�0j���`�%���t�ِ_��!�-~\1�r��-^�5Fų��BĄ�t���Z�[�:������٣��Wm�p��&o��8ֿ%}�)Ɯq� _DK'2_i�#YX!�|I�dU���Y��^��F��lM�5����`al��t?`}�sZ9H	}F�h�ϗϏ�h���)Bbs��6���
r�P6X�)��ƪ�#���`�>;`���Q���-v��X|?�F��_�$�rgi��1��*�h32�L-��m�;J���`��([��֢���<�xWr� �r]Lky�ă|��Bz4��Eo9`Fǥ����;x{7VN�|>�|%��������tc��Ʃ�]0�-4F4� M�}�a�T��vC�+���������[�&w��6A��9�Α\���g�7)I� W�;"�������9�k��)<K~��^Y�I�BJ���8t���IׄG�6yd�!b>��������v阿�y����Da�ܿH�n�RQ�P��2�K3�4�[� �+��<#Xe�@'8�^�x� ��~��^4��gZ�y�#�	[�OuK���߁u�=�[j����CÌ�����ܖ����Hr�r�V�fg#
��'.I_|�2é3�'D�e�����%��";d�\k�(R�ɧ��D��r9��>�ͣ0܅�v�^x�]z�(��ԛgl��V�
��,@d���+IJ���a+�+2[C� )�8OϮ�S�]X����sR�������n�:+s��s�џ=��7��e�-	��7ӊ_�0��3GY�QS���d�_M"�޸�����Ir<��R9�[���6�`&��/F��D�˗���ԧ��!D��ؾ���ʫ��Q��S�� �J��Z�t�鳘�s�L�l?NW�R���8�am�Z��R�.p �^��4�$��"+'61�?RD� S���2q��d��08�Ӡ����s��&�jA��0$�6��T����B�'�z�ouci�R��fD0����c־(r"Z+�p �����<)P78�%§z�"2kh���w�g�-��kG�^��O�Q6esmP��	���4��75)��RYݡ���[�/Ƒ�X�� 
�9ݛy���:O^�@�ɍ�>#�,�g>-cZ�+I���N��B�nL4#X+ �$�x�'	p۵m8H���D�no��IM�NjaaaŒ�w`��n
�$̓��.SƤ�Zt��i�s���BxԭLQ�\�
$�}�R��R�&�q�"ß��Fo�U�i�T�Q�[@qps[Yr������-��:��&�^�|ui,����a����As�B $���+�[��(�g<)�H]��x�3"w����Vy �.��=�-��VB��g�N$����D���U�N���.nj���iE�aS|�+H�+P-qC�۫?� ��~¸��d�.���i�8O��&(z�k�-��z�_�~=�3��F&ۜ�d��V��˂�I�ede�.=y�*���ۧ�ʧ�C�2�{��	�	Ԑ'�ߖ[W���
hƾզ�hz�O��ny��pYob��w�E$�9�6�Au����U�:.�"�qżM?�pEĨ���a�:	ܟ���U9��")��X��&gT�X#ȓ�����"����]���̢)4<7?�#����^��ᳯ�_��������j`Vyb��q�0Nd<�m�n/#�;���'~
�wi�LWA]��d�W�ݜ�9_�w�j����+��^���׼��?�W�A�s��븯N'\�фn�+�3( ۢ�����{g�\��<{R�g�1��Kz����ne�k�S�'�<Q����n�J�]������g΄�Y�A��'��v��Ea��w�Z)�%n#4��G���
�M�<a`�Ww��_�!4>i�?yz0�eob���� L� ����<`��(�NAw} �d�|PЖ�`�Q�g��"����y^0��ΰS���=̃�f�߻��α�vs��@�՝����4��sM}R��*WS�]�d℺F�wR�\�8^DP"�6b�!M'��*�}	M��B�Y\����e�PBQ����$7"eX���y��:�e�����`6���]=��ez��_)9?���Z6��:8��w��W����BB�L���ـ�b�U�*�!02�u�#/K��AHg��^�C��8渨�0`��6�z�T�x_�r	����d�"����-_��*���|�������]��� �U�8I�H�������w�(d��ㆰۇA*J��;� A�WSO��:S;���}����{����{,2{�V߱�p��g�"vN+�O<צo1���B����&oэ��&��H�����/��.^�84�[�3"Xn���-�ʫ� F��hߓu��$����v	*�^K�_T1�$�"�%ϧ�=�����?��HLk����6��_,���ڹ[�"��0��y����b���������t��z�h��<h�8!˔��O�g`��O�(^Y�������r�-f�nP�n_�,����#����DEo��aD�Mdk��ܝ�hf�9VV*-�����GQɿ�f䘇B���+]����4�w��}Nз�Z3��K��wC��G;�)�k������6�uW��X�ZO�!UP�L��}z��g�1#��O��hKa/���9n�,r�
��!ʤiť���.TjQl��,��@�ԭ���^S$9�dj]�N����9�o��w.���EA@�"�@k��|�Ҹ��2��l>"n �_C�w'\|�=�Î��H�/���G�X7]�R��뜊ե�Em�\��v�;c����J��ƒ�գyV�9�~�$�kq">�1w��݇��"ߪ����ߎտ�pj�H2d��VP�}�JHq{�[�,�x��g�@���@mK2R&���M61���k|f�)�~��O�r��mI������:Fx��x����V��g]<&ݦ���g�: �#*.�e'(���Ȓ�j��2lig7v>j�|���:���䨽3��m��,��X5T:^x����, ���� }L7 e`�.����Υ"�Z�W@��Vc���-~�(�wr���<ـ��ͪ6��]�M�|�OITe��^i'��_����.��J��l����֧�#�;	��@(����x���y���9$�RոiB��~47�9��T	�B�M�!R��v��������~�����-�]��-��lA�]�� �+ Fr��)N+G5��% 0b�é�ׯ�΢�r�-�f�e�H3�>Vm�~�L�����i�B�xG��E)��X]^� \�Ʌ�~��)_?�)�6���ʻx�H�ym<�1�2�ɬ�$z��?Vx�	`޽{)J�:u?�	�%D�F��W�)ѱ����q��҉�����ʿ�Q_^z�Z���յ���#���O�<��a�	��9��P�a:�O'�û�����r�5k4u|�c=�ͭ1w|HPA�=]�I���+;����$���{ʪwiB0�>&��(t�ʑ���Z��.�S�(��m�_|`����_�+,{�7��J��=x� [ܠ��+U$R:��&(�9��h&h��QI�?:�u	��&&&�9�de�e��a%%(AH����f΍0?l>�����K���S5j0��n�˪~�Ř�ݯ�A��+�����D��1�I�s![[��a%w��_K-�Gl�KO�/��ބ��'-�n$ǳ�F'@��	mb̅��X޸��u8���g�c�p�k2q�fy^D+����,�߹�Uq���䋠d
�%��Q��B���7o޴)��h=<)�^.����|�ↀ|!kNͨJ:($�ɯ@�Yxr-5����~���KY�C3)�۠~�c�):'+;��(���}��w`���O���~*���H���CV���7��8�bl(�894X���f֜���QF@�vEt��[����4�O%��^ ��^�.e��z�X��✑��y0�zӃm,]j���G���a}�7��?U�l?py.#Mg�<�*��q�fQ?P�6W"�Ɓ�P`����vʝ��C�TK���Y�V�C),R���u��1od�>v���vt&8qwy�t��nq�R�օ=��sv�2��1/�[�?��~��K$t���Y�i��,l<D�T`�� � ��]��䉬V!U�	0�v$�-o���mS���c�\�ʾ����6���ӓ;�V<�g~���l��^P#�}X�g$�*��`�7?Ō@s����Ą���n��)r�c��$L��9����S �&�1��!���c"�����m
�뉔�d�Ý��J���l��� �E���f`5�2��-���gE�����l����.lStidy2X߮ &��j���`��=j �H��(���=M��qO�5^�PրF�����1���0J���Ř.��si:|� ��!�S�� �W��w��Oj�'�
�`%��Q+��A����>��Ӂ�ɔ:�yB�h��V�F�]/�̇�gQuo��B��ԕ���"�l�I,�q�,�Е�M��������SM�l���,�G�+H��t����v�^d�{��K��Q4��9L�o�N�툁�l ���
<E��*�����;3��PԿǖ��~ڪm b m/8��%�Kɏ��X���|�#MC͸�MLY�y�C5�9t��|�G�B��5���#�����C�%gؗh�����dlf�>�&�����spL�'MJ����q�>���<oc����a�=��L���:8��6£E?:4��:҄�;8�c�dۮ;U,�i����s�99��X������M���[?�����T�ݻ��b�<������r�?�%�6��l?Y����An
�?ȡ�[������m8萭l�|���+��P��|����)R��-�j��m
���C��|��= �;
qar4��~#�q,����:_.$�.����kn�����v�?�\�H�����w�tjv���{{��Xw,�+k~2邫���,P�P�b bcU����+��m Э2X ��(J���\���em����5J��uP��6��i�aCN ��p�7�p��܎F܀[>伷\5� !`#��n?E����Q�}}�:�a#A�۷�x@ߎ&�s���������m�Av���	���t��QE�S��JX���8��J� �9~pf������q�:7!Z�誌��	�*,�>��A��	Y7(�G����:V����q(γ�Q��XQ��5C%ֻ�S�Ql'���{cgg�0�E�f��
���m�����rq�|_�dX��#��Vw	�r�=0P��E���	�~9s�j)� ��o�l}{q:,p�?I�P^�;xM%	F��n��'�=+W���u�S5��.��y�5G�$C8spr�7�6}��m~l&zS�5� �jNx���]8R5���ثVk]�i,D�SYλ�_ݚ��	�q�unE��l��4����}_��$z'���6���G�pzv�f�-�{�z�����/Qs8P��ͣJ�E4+|a��UR����X�2ȅ$ߍ8h���E���ǲDӪo%�^OSxa�
��薞m���/�L�b�c5	l��uWg���"3��W�a�������j��tO���\â�kfl{��g]duҠ��s�Au
@���Ӌ3CF>��r���L�H��t���IR�mO�+{��gn�ǎ��D�h�].�O06I� H�{ny�݉5�'�>����b@�x���q�4���?m1hma+Q�!�`}���ʏ�\�����XS���; u�����t�d�1�>gq"�MLJ�]�U��{\ǛN���k#XW1���T�ւad�]ZZ����t�Yd��DeC����`�4I�l����M��_9�'�v�쑈����>�!0Y�c@4=�DQ���ّ���!v���^�'��"��al3�޹��̓�SM�sX��H���e�)�dHFr�k�����E@��6��]���M��\vGz�Z�+ؠ�E��?:ǡ;��?����Zښ���YP�Z��ْ^f����Qp ��I�c!{�x�	'��o�S����cM��z7O^d L�-lp����1�a���k�:35����!ODV��-~��0z�Z^��l7�����iu�|�
h�)�}-w� Ӌu8z��*��yB���eU�K/!���!t�)�ӿ��iR��1w�l\h`��qε�,6��T׳�滜T���I��pw���C������������B
��d�P�#~��3N����Q'=��Ώ�t�,������[�`dv��T��W�_�KX8�v�W�Țu�3G�s*_T�A�p�UM|�,L�����V�Iͪ$�+�L����9K!�[�4��>P�A��o1Ӓ����A���Zm�r� �aJ+����3���͡,��r��g�&�Ã�#��0�ڮ���D�.���AN-|<�c������b)Y���#�WL�O/��&�@��e��w��P�f��9��I��S�(��u�h�*<�*�@�C��I�w����9%$$��.!���_49�I&�/cu�A��M�����Rh�n/s7�	���W�-�i/����9,`v�����N�DAH��v���#�Q\��#�V�5�^��ս!����r�8c5���5��� ��#�ӱ���u�" d�����)Lɢ$�Q�9YQ��0�������WͭV/����M�݌rO]���[�x�Uy��7��(�,�6l	��/X���\s���5�,̅����&����:��W��]QA���s?<�� ����X��,V���І�	,�#��q�`�
���k,�{�Ɓ�)�lʹ�DR˛�+[+��>�s3����3Z�=��_��㫷U�k�;�Kw���O��c�'�R(�m)�o �
�?'d�����E�s;�-ï��=��K�/�5=����Fq���w�}a�8�g�.��K?��c<��5����}�XI�yT�z�]$]�R�2����!R�$��w_,�i���BCM�-��������(3�m�K���H����?��i� �m�e y���r�7�g,�� �:k%�c�>>$!a��sz��wm���Og������E��C�=�+�?\����$&�Ϻ��\"?����?d�q6�u�K�d���d"�.M�h(�B��n�Rlu����LC����Tw�T�K��y�Ti|:��W�'�G�"�����6�[��h���LO��57��	���k���F�}5(���ͷ%�Y�Ç���n?���L���f4QN�546���r�#�5��H�c]b}�>p 2�>ʯu5�6�6Y�[�	���D��rf�OI�C��Ue�0�T��Cr�hI�N����K��2�Xt�P�T&^���l�c!��}k��B���x?#({8�H,]�ٌ��/�Y��&%�9�7-�u�mLy@�Mf�
7�D�g���`+MOL-7�_���p5:����|���KH�_��L��~!4��[]���vA���փ0'��'��@cd������7�⢉F�Kr�*K�ڐ�]\t�% U|%��g���QXι�������I]��Q	jQ�*�vNu�z=_�<}��rx�>ځEW����m
H~�ŝ��t��r���=D��lٓ�˨�e��D�kF��uh�䥅��\tykN�O��{���aA����WS� �d��=��bስPQ��oHrfz:P	���Gy�
�K������j+Y�����8f�=n�4�B�~����d�~N�����R�(by���ϝh������?��u�[��S�ຫ7Ȓ�������*&x�@u2W]z��-�d�Y��J��E�p��i-�����@!]��M�A�����7�d�?)���.!������Ay&)c�鈔YbI~�,��Ղ
	d�d^����f�3v�df�Y]9�TF�+,/�3�RnAs��;_pƢ���ۻ�i/^c��:��o������:�Û����o����}���p��8Dj���d��;�n(x��� *Ȱx������]�ROTHdP���5VF� #{�h�Spq��$ګ+u��V`������֥4�?h��76��)���D�f��,ǧ7�u��ЏXﮕQe9��Xe,w |�s��br�}����s�z`��r��+`?qv��@���T��7� o}M �n��6o�����:� ����aF7ܻ�s�;G���f�3���]I��J�����R��������?�̜��(x�̵L!'�SU]��)��U���j�<�~��c�3�V�u�H\�~�!�3#(�nq2��A�����o���ڜ���Xh��$�ɿ�ҋ�
�����2v�䜹M�
S�i������-)��L�����"�ͷu�j,�OP�k��a��To9vo=�2�S�&�
'#	˱�� �vi���d7s �%�+tZiEY$o�-+-�[n	#6��3��͜����<ɘ�í�Cy%�s�{�����-���x(2��~��L�˩�����x3�{��.|�D�^�d�f�xv�h�/��U ����oƪy�7���`�e�D'%j`�y!$""��*�YE�xܩ���\����^QG�1Шy���Ht�!�mB�Vdd$�A~��J�C�16 ��uĳ_z!�ǅ���	a�B����
���ޏT�Y�3�����y��6�,��?w��9%�� SM�ʑC�;h��\�cyR�<�7��M�0�[�92.a���Ӊ����`u�\�A�ϱf5����7wcq05�#���ĵ�m{��#�r�Y�gvx�X߂��$��Il��#,v���wD����2��Q��^�F���N'L	���|5�����-���<�P����E�k��i�
�/�.��6ċ�BYrò�Ǆ����@�&#�<��?��$�vAO/0��h��*�^@��'�v�{%�2��9�	�����6�qF�J����}���!�����?f����� /���^�E��՞yI�T��k�ǏW$@����=��$��`�N_�/�N�Q-��Qu����#�L��O�C�'.��`i#��g�r� |�}����S�2#��Q���8^Ia��߿n�
��@� ������]���g�k�A)�R�E;��  .�ρ�|�^h�C�Nq%����n���*��kF)ޓ��D\����="Ќ�t}/��p��K_C��Ƈ=��������U_�F��{�U�Txb��j��)^	���Ru{��S���hb�I������rb��*�Jr	 �U0_D���kNB�T�z��*Y�{KW��sH"'P,�]�OK(1��O%�
��J����Vs2�=2�������-2 A`H���-&.��
��
�dv�B�wJ�=��H|�71/^|�Z�GH� �܉+h�X���Y�a<��H�{b��\@[����5���00$��k���O���K3��:��^�L���%ڷ��h������l��r~��p�E��ز)���W� ����!��k���%�c�3��A�Z�bEd/��6��2"��̣��`�&).�Io}����1�r��H�bK'���\0sl����_��� @di*��ҙ���hF�^@����;�S5����['^�>�bemڅ�;��H�o<��[�O �C,�?����dVߑq��pAn'.�����c3�P8�GAԭ*�h�~Ya|��B�%!�����%{��~��m��0�Һ300�W��:j���J�/ �8�·�Y�D7	s�Dۄ��dx�vh����[�r�a��z4"kaت�1�&s��p�묅��ܝ���͚��K\��B&�������+Ag��s>k���P��8V(��T>塊�� ��і�>Ja�j������֍�I��
r-ښ���)��g�x����X��DA�	E�0�}W���oޮ��%s7���E�&8�4~�g;.
BW����Mf7�WU��?_����3��N�	�U^Q:K����=~3����M\ q@W��(��_s�G@+�o�a
�?�_�p�ä>�Z�k��~�a~��=4��؃{X*� �u<�ګ����kq߀d�"#
�����;pa%���]�7�ᛖ���"��"����Mޔ�cԵ߈2� ��<������`u�)p��']	�T���9�r�ݙM���u	��`c_;jP�9���Tz̊�œ)
�qΨ�]�uzd���0���q�7�� ����ᣀfbq� ֜Ob}T�@^��N����
�."'�555W7N���)#n�Fq��YbL�b���J��h��������0e�v��2=�"���p�~O���V=!�f�ͷ����*H�q)_`2����cs�f�e7�D2�7�����<�K��Ձ]?/����`o��H�J�M�_UA\a�w�7 ڪ-cs����� M�>4��FXI)�|������ভS�8���a��.6tj�_^�1�M��$&T�4{�T���E�X��f����Ԍ�j)%�g�Q� מ���oY�����/����I9�����W�8��.�.@E^|)�O�
�
,	#���
=,6��̞}�����ua�6_����S�	S/&9�#4GOu,3��Q�Ja8}<#��n �b�7�����Vw(#M���Uйbc�\��>W��Ξ'/����q2��k���I���
`�k��������eD ��"�:Y6���Z
����d,3�[e�S}��W�p'\
�����l�QP��XWu=v]u�:�~�/H���_р���z�A���?{�����-���j$�v�
�>�^��� WTi�uR�r�@QZx�4\�)��\Y%a�;_0'��~�R<gxܟ�A+�\s�/7�9�qKA�b8��2eh0>�o�{͹�{���iT�lF�ww�AlHi2���+��x$
�0eT���3*�x�ֽ�}<�RzL?��X��w��dȩ���=`�>�x/<w��>��:���Eo[�Q�o�PE�Gv"����>�&����l�5��'$�����AP�}�3�
����;
_��W�'?�*�H@Nd
��-�`�4��H��#泮R��0�n�d����|xAT���I��9� �o����I�^�bAh�F����)�����Ƿ�r�v���y3���Ũ+�$����p0��1)� �� Ľ9x�D�ٸoC�8Öc|����#��f=
tMͭ�%�$����C�p�y
�R2��]5�I���� qa]}SC"n��Z��4��>�Q'�U-A��Iƚy�
��Q�¨�[����;�'.�b��$�n������Q�8ލ|=ǫ�*g�;��=k3{$$d?�W�~�U�������
�A����GXl>�B���n2���HgNz:|:[�T�J���r�3�Ѿ˜��7+zx��� ��\��KJ��.��l\�H�������kcmY"ܽ_U��}��a!E���l���#����}�XKa]��з�RB��3s�� $y ���Gnb�<�\>��-���ç�p�<��`����|�Ǚ�Q�G,�7.�� x4�`|l%�{@�*��p��ƺ1Q�T�>M��/י��G����kQfW>ɔ���'��_��CaVa��$�6�O}]��(��l���7}5Fx�`u"�Ue��r-�D:�of�)��8���]7ȔH��*Ϊ7��%�����B��fsZ��-�33�dD�%�����646��a�t;~�J��O��c ��[;�ßS*v�T��5��'��]��6����44$e���țo����7�-8����ȵ������͇J��%��9�N���t��$��+����@��oCFS��kn�oٲEV�&j�D����5�����u,�P��	n��:��o�s"C�~ʢ�C��p~v��8醭�/����Z��j�+�A#�T�U�X��_�i'*ź�r���j:V<���������\�KO�q�f]cGɖT�Y����ϣ�6�ѷ��C� ���t"Z�-��ip�g,�F8-^`�ȋh��7�x*$��ړ��c[4t�PJ�yaOQʛ���$�tWF����D=�~`R�x�А�e!@�+�w��d~H�P��S�i^ g�L��s��7U�S� �&H����R�|����
R�
�Jḅ47KI���h�+!������
-Ji�J��wFb�W��ZK1�� =�����CI��je�돽��(���2�p�D֍J�5F��Pn-ρ6~���Y?���n�7"t�#�#B,>D�/Ř�x���Q�Ř�&y�7Mc�4
�@Mu�R ������%� �7�M�)�e Im&xyA��n\��8P�rk��B
a���YCjxwn~��#�ե��(���.5*,��(�C�Xg�VC�}��.L$�� ��l���S�
��퓼�%�$����7XCDǁ'`o��/�c���OovR�!���H�tfy�q���T�`��'?�c;��w�Q����J�{h�ln���f���~f�������K�3�< "i�}F�F��0��B���۸,���TUTU+Ρ�ky��F����B� �ROj�l�8�Km���<U��G��.h�b���Gq74l��א`�3�r�CQ������W>���X�?��G���	:CuX~�7�Ot��ϰz���@�@����2Ȫ��K���l��s����#:i�1e��)����2�s�WV�\�d(��A���k�PU��	��9hE��~}C{��g�R�IyASh%i��a�C���?-~�D����˙G�$J�k�q�-K7�g�ā	����r���h�S�����f��#✌j��3p[)w+��-���w\���(����fD��Y�VM��Z<7PS�\���0��ku�5qF ;�g?������ئ
���Pϰ�t���:�WHc2i������B��b��H�k��ȝ��������8h���-JoP+�.>7�}�,5�x���7�2�a�>qb}�,�����P����z����q����|�Mv!>�>� *�uϬ��	�n��i�4�CRO7?w��^P���&�s�zN!����Mq"e � ��NR!^�"�mA�H��݋d� �Ђ����,w0����c=`�AEO����Υ��J�O�k�[,ަ�.?�Lߧ�e�"(:�֕��&FO���]wso�!˫�-W�5���X����,�J-���7:���ha���^)��ŗ����bm��6���$�kL`�ƽ5�[�E3Ǯ�92��_CC>��邤�Y��'�@���r� �j��Z�����x|}8�g���TS�o��=����q�����u��rB���(`Xp�Yx��Q*��'1puQ��+���κ�9��[I_C�)v��'{��Aoc�:��	�?�kDc�0���/��R*��������j�@Ӵ�����/�D�'�M�5��r�_�U�Ӟ!,<�j�~/޾OGi��'ɵ`���(=�=�३5u�9R�/�Ԙ��8__5vdDUn��[�vtt�d���Z&�*S�z�����H忀U���MදV�XJy��k�.��8N��V��Ф�+Q~�_3�e�	0�ȝ������j��*��-|\Z�Ibg���f�.@e���%�aT��
|t�Hz;�p�:�+.��ʷ���N�$�744�	�xa�c������HQc}}ٟ����i�o�ZZY��,: ��	7=˲����+:#��؅�L�%~F�ze�\�nWM�j�b���8��*�_��ȳn��P��R�>��!�謹�2~�Ⴆ��xC	�S�PNs��MY��s��0a�%&nz�%�����ŞC�z(}}} �|�ɋ�Р�-�����K�JT�}\�E]?ɫV ~��=jS�&E�7O�#̰´;�c���d�p)����?�A��W �i��w>�	��b@@$==6������=kӄ��,A���� �b~.����;	�h�4����Ă:�߂�P|�[P�?xc�U_�b��e�i�p�6ڼ���!<��͂EC�')��|�a/,�����8#�%9[�O��s$��hw�)t��kP�'@;i������,l����z�
�T{�M �<';��B�S_2���Llܩ;R��x�(_ȴ Xh�1� �� ����l	����,딭T��	���ŗ��>k9�@Y�.N��!������o,W�Da*$
=��Rm�ϢT�B\@E���Ó�	3��u�t��զ��Qx�������� ܛo˪��B�"�_�&׃��x���.����:(�_\����4�+;h��_�� iS`��̭f�� ��$ʕ��䓤���mco��\�tĝU��XW>vp���	�i���`����X3��H�J �������w�L
˟�ռК���=P�:�u��Tw�j`���x��F�h�C���P ��D��#^
�N�r�sΛU]�
������}�<�!��D#����;[BHJ�@ٹb �$;����n��yGK�Ӗ�6�?`SP��\�{E�.�����H/iƥk=�(�X�~r�.�=�GGX�yƦ�e�R��"�3��!�R�!�v���m:�.oW���{�����6v�m�e�Rm�o 3�SK���n�#�S�&#PE��,(���Q���*or��鄅��F� ����ս�^�\y�s x+W�Љ4��0��ӭ�����x!��-?t�(P{ɀ�T>�x?"�����(��3�O������
[ %-#V��ˊ���S��(�$A\d�����
	\�E�l���R���A�z#��^OᲠ�;x�ދ�W��[F��yQ����AXx#�.�uY�rQ��Z7U�t�5��'�a�j�p�BH�1СD�k$a3}!EU����20��n/`��N�x��{"<�@%=��U}��M:d�⮳�h'�މ��؉��gi2p��A������T��������v���^�i�(w��sHg(3`FdV�����0��bW�q�mb���D�Uq�R�[<�D��+Dxu�H����Eu` _悝��y#�Kl������v.o�+Ԗu�\�Qc�@�m$z~q'e�[�_��-'%4�A��f}��}F�4�t�
��{�� �A�G@�J$�YS�xr8���.���X��k� �ݘ���
��in�6綃�Y_�P�=�܍��Iw_'m抡!IU�n�s�p�h��ē�y彉�>D�$~�� ��Q�[o��r��.�uK9P7��p�u��+��s���YP_��WWלzy���\��ˈ����V{򕼼�
�g�ڊ�=vU�a��5t\�=��Lc�@<5��o���p�G��gL�����r�԰�l9��v�R�p����xC{���8kB�� rj�������w������0�r�q�"�7	E�p����$_�s
Ϟk���wi���)�a��̜�m�>����������J��.�5~@���\�{��yI=�M\��I���4�sY��'�&�W>�$YK�-�6ns��7���)��?�]'җLU�͊�D�ղ��4�?ͧ��%M'Ɉ�
_�l��嗀�ڷ�
)�7���(>���Oz���K���t?�ϴ�8x�K=��~ō�&�	P�j���Z��<`�V���7"E"rνm/W�J�4v}[�� ]����ڵ����a;ZBנ�IL�K������)�m�Q�e��r�O�&�m�b�"��a%td+7U�e�_T�;
֤7�i����Ei�"�3�����So�d&\Ϣ\N��,�A���2��Aň� ��cu�}�P��Y��Ih�����ݺ��R*�R��-t���q�?ޘV�Y\����D�A�/�_/��_���,�t�8(��#��~ߘ-\���,��r�_V�oy|'�=K��Ȩ�:��M]�k����T
�������F��n�zt������UzA���`w"^YQs�h��hK��ϩ�*��ʿ ��]��C �[j���x��Xj�Mf����?����]�Q�ZJ�{k� �����!�&Z
RK�J�ӓ�BG������= N���>*��b@��]���"�a��
�bر��}��A~��"!������&mb-�7�B�����Q ��0�޼w�Q�}h��f����ڬ����N^��7��0PWKss�>^i�ݖ�=�8��%%KdB�����F����&�%����_������Y2rk����GM�Q�-�_��E�����9�	�2ڮ�<6���N���e����e
���IL�񮢞��4]�0B4蛦�b}���)�zM��-J���y������;�[�� Y��I�����E&�&m��s����&������o�=�#���@ii��Ԓ�d�\>sH�2��W��X�������l�>�̞$���e���[���;p-�ʕ^x�?����ڮ!.+��g�i�y���$��w	�Pv~���^=�x�sWQR��k ֏����-/n�=�~�������B�͸�D���O�6sG�Od�����~����D��I�䇍D��9,!��tC:x�h@~~��1<V�脩�*�g�C5h��׳��R>�D3˪F9h�(� 6�k5čv&��dH�u{��j�C�4ůy+	�J��������;;�Ia��9;�q�>4���tk��Օ4���pǻ
m�z룖i�i3v$͵��d����;�_}<j2��+��g��%T@�N�U�z��Έv��z�]���jI���e��CG�e�CCN�� ?s��Lp���۰���
!u�|�?�;�R)c	C��l�3����H�d)�Ό���L�h�*�v�խ�i�qX����a��6����-B���		����'c�O��eɪ��̯e��5%��	��L>���1��P���S�j?I;���;�کDQd�6�+��v���r#�ڶL�Ԛ�:v�D�FD)Tj���\�����|������>�O^����<���}�1���o�6�2�*����qQ�jK0:�Uӗ��QX�:�y�r�yH�?�:�ӑ��眼������l���n��\��d��!3x�X�ጫк!Z��3m�̆i۫�<¤��Ɗ/�a����g��� k��y���T�K�ȅ�H$�%zc8���	��g  �r��۲u}Ǟ�O���E��UxDo�����d'��`�<EZ���Wkz�/��y��툪7&KFoG*��_���*k�,�$��l����:Ƅ��ir_�Hz��֪}VYt}]ς�tz�s���������U�))����4Iϯ����*M�l[rVi,�wdk���ћ���+��:��a$8�2iJ2c�u�^89x�v�.�(uy��d���5J�+VW�Y3Z���[�[���P�u~U�~�6�3��zZ�a��ik������#�4����?h�3P�#JZUʨ�ojP���S�'xG\��Z�DƆ���_Ά@|�[�c�DOĄ�k=��
�rԴ��f��5x	��o���y7F+�\�C�d渫	�����+��B�8�Ac��t�p��X�[�E��g뚚l]�5��"��e;F��e���҄��c6r���T[ޒa��ݳr�Qz���0�*����hoo�qQ�6K].�U��B��V��F�moS��7c?�
�w�	��3
�6����]X�����|��Aff{��n( �t}ާ2}�G��f2r~�
�|l�è�dɥ��Yw��?9�������̐Y�ݻw��ęv1���t�ޛl�������ks����t2�w>lly��Sc]��&�G=��N*�L+�0�c���X%��%���z�D�S��ڮ��z�?����,[U���l�����U �a�x[��PNG�*��.�
�x@�{�����P9o/X��{6���YoK�A�.X�5*R�~r#$��4,��{�r��3��|1_i6eƳ���!4���oI8�+	��1�D)�u�H�.ƴA�Y�#�+������u�5����^Du�p͗G)����L�@��#zv<^�42=�ly������ٸ?|�J�}���Dʖ.�F��:)�p�z$|O߹$x~��u��n��ٺ,qger�ܝ���_������Qzy���?|�W1�#���Z���怱���3�켦��K>Y��g_�d�'�?�CЈ��Y�<�'���Д���W�rf\��9�RN����f��Nn����ˏYˣ��E�=0n��3z�����/k���>�J�W�Pne��1&�����{�4C�ɜ'3�d�n	����݌���v��0ߧRr��*�2MF�+�eo|��g�^�Z��_���$Y�ϣC�?������8�����?��b�1(�|֭�ͺ6����#Uf�� �ʇ�(0����u}��oK�?q���P5���k�ࠁ�DO���ōC�+LOkY��D�v[���?z�h����]�n�r��D���Aڦ�[�Z�H�S��Rt�_�M�����2C��pT0Zʈ&�_���Z�ڔު��Y}/��4�k���j<��w�\s��++�n�z�]��nݺ��rm��^��/�-M����.�^�	[Me�-��ؤ��T�=��T�����GH���>媙�l�d�Q)ڲ+��Ő�§��i����/]�LH �:k���7��cizZh)�X���"p7�w $d����O�=�p��u�|g����={
ft�g�>�$tC2C�`��ӵ~�>U6�y]��2��,з2�6��n=,1糼�ub��.A�Fk�h�jժ������8�b�J���^ٺd�[V=׍=�*nr�����<w ���p/�h�	��V���C��wP�{��������ޭ�'�S&�R�p	��h��\x�@�\���!7���bX��{A7��h}8�6z��͡���S��s'�����!S��#�Qc���|����*���17Wׇj���h��[��Y�;5l1O���"!y[tYk:E�7����fY���=q���:6�-�(�m̛Ce���3�N�W�xW�#[�W �Z�,]qx��^+���I}z��^���&�I�Q!����cj}13��k��R���g�yx�yN�F��q��?���{�	��PF����l�Џn�b�o�b���|���^�N���/����-kS��Tq4��Z�3�r�B�z���lK��f�#�Ӂ:���D7�ȦH���=7o���k`�
�1��#�AY/)>:�W�{�l�hf��Zv�	�c��������������7\(�uj�W �N��l��{���$��苋u���>9۔�$������#���T���2 y|Z�@gw�^O��`�M[W�MX��f���S*;m�Iz�'>�h�5�8�8���&�=��E8����U���āU]A�|\�l�$D�T�`���:��={6�H�I9J��g������r����Ѧ˯�}PEȁJ�%�d��XQ�eYI?%o��rq��իW߹hi�����xN�:d;}*�5� -��t�c�<mYzubl(����6�	�#1d�K�%���"m���HJz��-սLt	5g�J��X_Yo�s��
^�ؠ�k�2�& ތiw���왽���:���BQm�\�����^�����G��ܶ���)�g� �X�o�~����1P���T�Q�1�c�����'��+�Tq�6<_��.]����BV3���[ �k����������j{� mn��[^�%�F����瘌��t�?^;�7m��T�䌥�H�9]N��������6� $}�w���h���F
��+��TqI�.���f�W�ac� �#����ma�m�zZ��%�2TM���ɗޟ���ڧ~(U�ƞ}`���<x����cW�i���4�U+;1ў���@7K���B�&�Ա`���۱e�{������p��Ak' �=~�5�5ǰ�o�1�� �Z�?P��d#�����2H��[7��t�dqS+ �?��+�M؟�5�Ũ(�12�c�*=u��Ƙ��x�IT�剪�&~ݜ	�g�<�8/�x��̶X����'���Ş����Dp�l�uӋ���<�'����ܽ�_�qyJ�鷭X�v��_�j;��,;[���g��,vVm��O~d��	�i.ޣ	R�}/^�P��� �^v˕��]|���h���p�=zw�ԻCk����^���b
llV����U���-���:���F���͒��(}�$4���b��x�ET��[j�;�1���$�hPV�i�d�Y�{K4��ݍ-��1�1�v��yg��)Wa����H�� GE*��j�Mq7�Y�f�-'�q��y����ؓ��<-�q\1svpu�u��a�����͋&��j@��U�1��A�|�Uا~��Ñ�8{>� �O\�p��([����	���f����
���V;�237D�B�W���Rl���]�@�C�M�8RƀgqY�eu�7�
xC�*�(�E�������K��v�o(����&�O�|���p7O��˭��1/(��o�ÝW"�}��A�D���A$Y����$�H�D �A*�w2Nvd�pt#�'2#׸H����5���%�K2즋���	J��<gK��:�2C�jm�\���ŤB���&���:�dh��AAA߁zd�ܚ��TőGM���?����z4p�W!����H�/�RU\�8(.��ďo�r��m���s���v��8�߾}���Y�l�E���d0���1aZ�D�T�RY�0`-�ڠ v�:��+ǝ�ך=u���������ц[";���(_���k.�	��Zz$$&N���d�z�����5��זSJɔ���lv�x�38��/ၦ�2��Ǧ��*RԶ1�vT0�ֈ0c_�Y(��$-|:6gA�J���9�@�5��Eͷ�V�Ҵ|y/�K�������(����;���{�c�����'��?ЛN�6�s2&�*"f�i��: @ȸ8� ��ĵ_�%�cM�c���2Z��I�'xtTe��<yv�qY_Ֆ�%�*�1TW�r�����0Z���E��_�U��k�;3��ȋ�)ψ��t	�Qp��p�.�T]xe�:��{�'��7`�K[�6����K��tjr���f�Q�	>���/^�x��0�V�4������ŷ@
G8�S$o�!�{r����M�܏��XkC�IF󈃬�Ԫ�����)�S������q(C��S�9��S�]�C�%��>��S`.&����\��;+�-�/*�hx�`0��3Zn��!85���uP�o��w'ϫ\"�:T���?d�"�8���g�Q~R�����U���)���j�L��M���v��VDJsʯ�@�d�R�G�۬R��&�Z 1aV��S>E�֍0`��~����U�g��7�]��Ѵ�����۷ӷI5��Ac��{n��0�}Rm� ��3� ��<`Mu�HП��rW���Q+,�.(|Y�����h���5�I-; D�S>��ܲT�x�vf�O����"a��>|���2$����L_?�$���\,g@=A5t�2~y�)n�z#y<��������-6ɟ��S%�q��ѝ�����t�2E�Q�F��@�8��O���Ą�����v�{���T�P�?\r}p�s�_��%J~6�S��f��g�Wgս�d��[ϛ7��ۊMظ����:M]& "��0����36�)��h�+���O84��  �)�a*�����@jA�2~�A&��}���ц/�P�܁�۾��ϗ�;@.�����1�Ucl�����L�'�H؅.��_Ng!�U�:c9u�{%R��UN7���j8$��'-�{aL8�q�Y�r�2x��g�^l�ߍ�0@-�۬�"�beg�Xv�(��3)w����yI�%���/2�O�� ^�8E�i���JX�b�޻�9��.��s>�Hm������c쵗~����;+�D؍0�]T��h)Eyx̼��Wh&��͓�ͤ�����=�|ˌ�����>���HO%\�:��;<x���+e�x���L(������pH����j�"��Ծ��s�dH�vE�o��y�Q����Ⴏ�m�
��yvر<��B�CZ��_AgM�w����ן}w�6�pM���h4���x&����/_�� �N���o(��� ���!U�w~	�5,�u�\��a)��������%�NTpn�
��׉L4�A��Y����俪���SGO��g|�>Ud��@�尊ᅢ�o�S��7���h ��׎�����N,r��~}�����9ƅ{g��}�����=3����Q�p���H�O#m�ѩr���K�_(��t�%�����9����Z|7pEe}�/~�]ӝ���is�p2t;v���祟�L:��H9��O<u�� >_]����R��l�����v@�K�F�C��&LC)�����wVϾ���Yii�-K��z��&�F.����R@^]��'鬃*2~�)��{��ŵ�D����4�+��?�J?�"틽}*�7[�Th�?�K�H����;�O��Fv[$���䩥y��a�2(�6RI�_^7�_NY;�&A?0A�I\!βt������H���p�J���,MF(��K)�zH��̶6��� ����0V�3�(��,�Q�?6���N)���<7.�2��"����`���$Cg�%6�'��)G�[r�h�Y�/����Gzr�jz:m��ֺ���$u��A��_�:ceY�Ju�|�k���jeٺ���gp�X����E�	=�M��E�t�^Ш�!믞Bq�Z���M2쁄Ze�T�\��u����P�"���$�������iԊԓ�F��A����?G)�ڔD:���H���50iŝUu��h�,�8�{C����7o�$Ng��"����X"a�ݻw�~	��ă��l���@�>��e��?Y�m��x���-���{�yr3{)�E�����'O��n2?�1�s{�*�<�Cv*���A�{�p�����)��h��_����k|˜�^o�oBķ�l�i����g��2_������#'�w���t��<ٺ�+�v��H;Wx�k��Y��i�|�iSF�}�,ܹ� n�wt4�i2���F��
��*L�x��.���"^�o��2b�[z��¡ӼK�N�hmg��<����b��p# �g,�8އ�'��P]�)/l^O׭�6�eɐʺ7������H w�B��w��Ԫ��$��2�O�㋸{ͷ�#)l10h�Ӑ��й2~I�橶TO��=w��.yP��>I�E*�ee�1J3�@kd�-��'-]r���3ɾ�p$�7�@��������P����+�K�d���ʬ����
�m�K��/�/�/���L��|�:���GIw맔[6RȪ�x����-l=ұ����k ��l������1������qS��ޙ����q0l����ӔSs�m�@Er�vW�w[������?�D�
]� ��j�|s�ȩԲ8�S!�u�<�s�o(}� ��'��`��tЕ���5$RD<t�$`W���$(�ڬ����XV.s����ᖠ�Hr�~���8Ƕ3�>��0����?��=�d�b��^�,��ϋ ��R�=cY�5C�>ɕ#7Ik�;�N	i�*�S&ُ�i�_�S7�3�`i�2��l]�HF�ȍ������'L<�e3I��VX�e���'�eF
�S��ݑ=��N���1���be0���s�mfzz�4G-/:�7�E�חnh�I�<�/�,���\�k�&qky~�YV������P�0�0y�t�&S����#-���C�1��$i�6aF���aA�����KM)���+"x��qGPYʊ�EvS����x��t�u(���V�"�Ӌ]U؜f�D��"rMl�Ϊ�����2��e)C�i�W��M����5N�l�dk��Yh�������b}�7�Cc%�-�f���M6��CՔ�7�0�Qm�';�u ]�����{�/���bYֽ��lmJ��7��﷭�ʌ$;�{T J����x,��̀�wZ�ԛq�lzߘ�S}�u�'Ə�l.Bҏx�V�'a��W�榆u�NIx�BF�w!{�ۅ�����v��l6�#Zq���7z�HrH�JEo�zDփ���`Ҹ����9xm:����8Kv�oq�X�#�����Y�`g2��ۅ]��m�])9�k�+��i��h�Oɒ�խ��T8��k��W}�0\%��,�����Tbs�I�1�ɠ	()�eraW�hN��|3<��*q���7��ߵ�L�k�O�vKă����;���8X�7״��.���P�1���av��/wJ��V�7\����2R>Ov�n�ݽR�������9*�W�]������O^���×M�ct;oU��Vm��o�v��u��Yg�zf���x��w�ï�ύ`�0�����>۫���Dx�:v
n8�L�U���[�;#�c~���z����X� ф,���a��s�D")/��,�w����>JN(�d�]G��
��jC��p+���W+�oXv��鞬���`l{�ΏNLB@�b�*lκ�ƢbZ생�(F�~�5��jpl"k��м�^ ,N�Es�݊����/E2J����~<��,��m�k�;T���M�E�q����k��ߙm�o3�cU�JG��E�>��
+D��®!�Ҙ������'%=��m.�������x�+
kG�
�*e�0PST٩��L.���t��7|pHy:b(�m.A}�c��N���r:p�TG��
�Y�ͼ s�)���u1��>F�D��O��P�a��Kxr;"Ư�!w�$]�a��ŋ�t��D�ʦg��63O�y���۷#�lH�,�"=�4�U���͗��省*�F]CÐC��F�Y���]��-3o�v��B)���V!����A�У�Y�z�mbp�5&L(S�5JiQP�V���999y�x���#N����MfQ!iz���&��6�v����~�OwV����i<���J���~�K[ۼ��*T�t*U("PBc�l|)�m�įܹ�Z �e���Q
zJ�ɭ�t��P3Ed�'W��e��E��������;�j��p��W��ӃRk�sz~��?D���e"�&����4��\E�J�1$�%?�0��6~G��D2��\�21��IWG��|L׃�o���BzՖ"G<�Ƌ����0�F��L���#�c8]��݇>��x��ͪ��F I���۠��q��T{Uî�6Nb���=�}C��J3kd�~d ���L%x@$�T1��F�(.Q�[��N�Z�kj3�|�#k�QX��f
RRS�#�h��&�19e�l�n���� ���>L��g�ʃi w�74<���x6i6��>��;�	,�1�Re&9��{��7p���\ض=Mr����W�0�dh�*"�{m�tY���r�19�,�0�B����Eb�<vjU�>cr+�3w���Ȉ"�6܀����?�q/]�l�#ct&�Uw��!M��@<�Ѩ[�h�4ة��.��m4���r���՝�t3���;���ީ�6f�yHS�(¥���#胓���l�qK����'�>�@O����y��'C������g�D�nc�7z�#��kW6�5��a]$���"�4:}`�_2�B�	S{K�+Q~�/�Z!�f\.VRC�{�iD�q�Da�\)A���ͭg��u�y�?]�UVq�O|C�3|΋̞���3.�O�5��wE���`�!�u�5�h��Mֶ�Χ�LE]`�HW���X���=�ʞO�2{ 3�ǭ���:cbb��f�Vȅy94ɭ��[����i������q��%�X�BC��U�k�L�q�F̓���ʬrugʚ,~c��b
Z�`��3d���Pl# '��Mr����g��y�U��V��T���ek;�G�&�e�2QV����m���o;}�Ew��O< W�?Qxd)�C��>��*u��G�j3��QО�����^ZH��+����g3�xH,�ZAu�.������U��s��OH�ѓ};v�P�.��@���~�A6Ο��v�i�]���1�_�X�%a���s��>|�p�e�ֿ�I��4d+xI�&��V"�R�
8"���T�uG4{?���*������`�^������u�&��3�"�����,���i7��/�����oE�~\͏8x�<-���"I�q� ����$�R�t1Z\��/͓�ʴ����5�)�W� ���"�zZ �;�{��!3Q�r�ҽ����T.�wH(�7��D"���L��La)_�_�BI�;�+!U#4���f����t���4�	�����b5��mP+���ӓD	��TP�`�1`���z��e�LM^�o3Z20
bL�r��\������t���Nk�f*9��qn�|w�m��q8�d�0c*��D����{wb{�Z���c��Ϡ�J3����2�����Nz�����������`�ߴ��򳳇����svoڙ�܆U�r*a���$LI	��0�5��X���l�)�՟��/X~��q��e�?�P<��/�8Q%(��9�X/�z I��[.���'c��cb�fL��7���y��R:������ʄ��7�z��!��w�&9���W��e�Wmj>���#oA�p�t[��t��s�a���Ǐ� �^!�P�Pl��H�����.��Ii�ع3#[��iD�!R큙݃���Z��*o���ea�ABiԼ�S��/�nTh�!�d�L��0V�K�݊�<�R��pT��!��23�;��f%v<u��:�}s�+<������q!m��GP�v9��$�^�n�7��L����+�����$��`_��]��t��H[����H��.��۝���[��J������&��0'���CUH����z���Q�]����Y��6�7a
ȭ�_�>/�VL9(&K���-S� �J��96�=E�AY�	��2@�p��R�'� �P	���� x`ͫ�#�X%��7[P&-AM�=���/�O,�ͼ��f���C�wtrJx��lH(�0Z��l�)p�ؗ�
�#]&t���uga�<��f���I3�0���w����& ,~kV�>��5kx��g8�D�C��׼j<uS�8�WC�&�Jڹ�z�X���ٺ��e+���������=;\|u�TA�_sCd��;�l���
l��N��à+I��O�.�L�+}B���V��)0���{h,�����^�kܾ���8]��]�~�2)���z��d�!�s����Rk
`_�A��__�~���?��y�����+ʸ͖v&�OCA��z��G���.Zl)j�{�DKl���mC펈��h�ec]��n���4�-�.�Ķ�C���"�NS�I�~-O��'�[���)�f��n�m�y��G����/���2�M�ry�����O����^�#B�7g�,��dp�ˮ�.B�G�nY�M���(���_�]�0��֬FI��Z�=������[�*�u�����!_q��V�E�H��Uf�(x�vz?9�$��E�
�	�>C�	�h�N|�6�dLK.+?��Q}�y�?���P��k�3i��x��T$���>άV�"���z.7�m�U����͞G��e�f������re*8L� �!��t��*��.��0 ���f^֕�S�ںu�&p�I"�r�a�ЦÞ�-���`�������I��H�
`��"�<׫]��T�<zqWWW�h'"e����"�W!!ܹ�����MT��\"���_QQѐ���Ps�Ifіo����Ca�L-��?MF����K��Xk���#I��Cd�㜮0���`�0����4�T2g������r |R)๼�;�l��}L��,螋Ǚ
�>X;8�$R%���$���G7��l�W�Ֆ_�L��|�I����ζ�_�� >�C|�����Ј65����KO����N����;���aM ��t��Yw�،w��l#NM��#-0�,��5-"'���#�q�~gd^c�^G8���T݋'�=,M�La���g�artF�����ଞܹi��_�5"��l䗋�R���[IM��G7��D�\�F�F�Pi���ǻ3�i�SY#x�\�IV�Em��u^I�YY��C|��*2~ў�6�f ��?����%�|D���߱���E�����3G��rL3���/�_va�\i~�6x�4ߋg�_�7iMXVj�C6�Le�okkjz`�a���~i�Ta�9RWJ�x~��,�^�= >��"�`ŗ���h9�m&�=h��
]�����{�h�r�l�k��ξE�����N��7Ev�%���l=UJ�3�4Q�o���ƛyQJ3���f���4aVm�F^�v� s���E�nkk+a]��7/Hf�<34�|�H�ōe: $��L��W5Σ��6o8ρ�� 0� g�m�Q�CH0� �̦���7�K�O��V���ߩHsX�-�����ᴍ�(�rw��,�	���'��ѡ�����9&�v��!Aܹ�J�JIuHC������h�I�zY��������Y8�����XL�y�X�/�
א�� }v���Y�<�ahlN�j��ٽ� �hk���+S�#u�e�"k�qj�/��r�8��;K���b�~7-�s�t�j�:&�ފ�����"�wt>҂��{c�j��O^���7o^�R�py�2�D�#bЖ����A֓x$dj�����	ji����0�5��kN�~A���cs��ƨvy�ڏϱ�0�_ ���ǏW8�Ӯ?+;�&��r���7�{�Ŀ}�w��	£�6r�f��TByu5�	[�\� ٺ��7}C���F6��xu	��/~n@V�2*"���/�I��<�X= y��d7����?U������؈ن��3}�d�ݮ��} y���S=!�*e��i��-E�������Z(��J3#6��5�Xo��-}
��6m��,�H�������%��4#��C���F��K�f ���(O�����B=!%ޡ۬\f�9�M�����<-�U�Ma
��2T ����=x�Ν�;�G&�~�'�Gk��a�Y3�9�����w�����?����Q`U�;w�94��!*���NB���c��lU�mΚS�!tg6�o�TBưٵ�����nC��GB\\N�[�"yd-��<�B[[[=����{+n�O|�L�����ܱt�019o�л|c��<�_����@�~��v
��K��f�g���
{���̇G�������j�G�_I kWf޻��H�¸�)���xA���е�5G��I���W��x��du�f���t����,�O�͡���?P�	^�����Q�h�_C�gL�)@�&��tPRa9��*�v;+�I��S8E�jniiiܟEk�+U/��Y&�'�檆hib���j�j)���$
E7��E��u�v}"���l�aI���[��u�ZЃt/Xh/�S��pF3�;VȖ��`ĕ=�	�[#�Y(�E�榥��od�I�����[N1[}�T8�n)j\p�n=�r�l�-���G�I�̶Nҍ��
�,���?����:���F��o��Cׯi�n 
ȝ�U�i�\�ϡ�^0�m��g+�/R�4�{�����NK�ݐ6S�!/��Js3a�5oM5�fCU�&�y�f�$af���8����8�Wv�Y����=5N�P9���bg>�6O�Lj�N_��+-�ˡ���ʹ�Ш�[6`��t~8y&I�&��M��i8�����n9]P6�[m�05՞N!~q|+��DeɞW�>	�䎵U�γJ,�>ҏ�n��$�@Pi0�p����:^�T��S�K�E�>��G��+ G:���%������Ѯ�o�YRi9��c� f:�w�ˎ4�?~�b�b�k��8U�{������D�>-ʷn�b���h��V
ƃ���n��AS�H?lɪ�8�l���_����ŝ>DZ=�.m�Z\�W~��E0�
d�P���#���r+��c���Η�9�Nt���ޢ�Wj�A���ڲ0��=:01ĚRώN]m6[)�_%������>���H�c�s?t�S]���kE��c�%b�8��8�`�b��bi�����2{vѐqQ2f��@�8�k#����q�#��A�*����kN�s=���0�Ư��,p/N&�4�jժH
L�Xś����9��56 �k��	��$��(4��h̘�kyA:Pѳ��,j+�$Gv���5=�����[�n���R��xA�[��`36~Go��(ӈH�ۊ/c�,e�,pX�/��x�U[va�+���G�r�G˟hi��t�T�	��o1�Q��/O�8�Sǻ�����:�$��-k3�9]xJ]��t-�K9�vqP�k���<B�w��Wf��J�k⛱��S�a��������\nF�!�']��;�I�+��6��v���!��w���)��3B5}��+�Wj���4��&���}C�U��:��U
�Df�u��@)�f��o7�a���������p�K�2�K�	��8��V��1J1O�H��Y,��($Ni�g:|�5�����xw�4�9sfu����G���42�]�0��A=V{@=�I��72������WV���b}uK�
�"������/_3竦?���-D����m���,�7��as�[�"my*$�n&T�]`�N(�ŒW�^5����e4�V{ą^6�Ma@��k����#}�3na��:�:��f�AGۯ�k�ju�J��3d�Ν@(�FDZ���Ɨ��&��t�=�����̓?����!�춶fR����V�"���6�qT�y�I��o�)��5�DŞ����d�!Ae�M�q��O7~�����7�3�����gk�K��W���(��3ߖ�ʠ��%����9�^	��;Ry<<��r�K�ܚ�H����p��-7�����n��vܕ�~*V��Y� h���1��u��R!��J��z�S�D�T��zU�ܺ���(�����GCdZ���l���Z���&��Η���� �\�t����d������o���B��<IK�p�x��W��������i� +5���5�Ҷ[�y�`k�:՘6Ing(²w�L�'Y1ș��t�t��c��>,S��_�=X˅�E``����=����(��%����@�\O߾};BY���i�E�+X69�43-|�dU׀��������ַR���:�o�۠. �w�K���+�=� wy��4�I��4�՛�o���nd�l��cÝ#6�PHz��,�DEz=.�߭���IU���%���jg�e�i�{
���5���,��*L���y��3���{�]�sC�Q���h� �Ў��ʛn��R6�l�=�*Ќ;Kl�d+U˪�t���(H��TN���\1�����>�h����_���U�X{���Q�Fl�Iq��(��ԾV&�5 O�.�XX�|��O��u�$`�4R4l��?Q�+�����`�%��2�uG�<�~�x%��,Aa�Ϳ�Uy([5�3+ߛz0$Zw���n��4I��y|͏�%u�a���(z� q��چ�!Ե�i;?y��Q5�T�����G7P��SP�oKIph�.j�f��iM!�G�����5���JI�J9��������YF.^���H_@���4�=9K{5�47��`�������ё�׍U�v�i^O@��P���
���W���E]���d��h���h������J?�u�0![��,��}'�� T�*#�G��"I�+�C���&���`i"<�q�����w�6�o��I�z�
��Q�nv/m��@@�d�&Yɑ�L� ڑ��L���{sy�rd�Ty�<�4��ʷ���mץ7i`�Ƒ�5��m���P��g��_��գ�XE�6��De���p�-n0�"������S��as�?C*��*�!1a��M�R�F�Nf�Y��x�?}�I���r|�2�o���$��q��dQjt>�%�}?4�q�g�p�U�0�)��bzֲ�
mծ��,ɠ��m�������̐���T$y�q��W�8t'������Ý�-qn"E��$"�ee<i๻1ǯ�R��l��L<+	C���� ��S�V.w��g0��[��ܜ��J34Je�f��@�:mef��4aYGT���.b�D�+|���G,�f�~�vD������W��L�Ba�
��"�x��rI�.� OW�������j:R�)�c?y��LX���p�W�[�e���s�U�����a.�%պ,��o���@|�_����x�y��p��O��m)ڂ�g�>�:0py�:���;�-�W6���i�>�JY�.:�������!8����S�7�aw��&��E~`Ǜ���2񮮮�,��V�+��+��cf:����+�u�%�����ʑ~�kˢ�{3W
�0�Zw?�,�nh�s�z;j̶��w��qd��C���kI�z#x��0����?����Q����g��+uu`�+嚯����G�R%4�+:�]r��`6���l��/�T�����I���tA
�G����<�������Z��|n)Z�4$D�@]z��T�Y?�	3�Q�/*���#�u-rP�$���0�7���1��X4��(JXLL��-E%�.��M�~&�u�����G*�g�r�R�jQ�UY����*���������[���v��Xs����88��wҦE��g5}���N}K'���?���?�����;�k(�f��C��Z���Ǝ[����u��]����<�g<�M�s�j�_޿�b����J��ͅ��(�.����4�%�q[�n��2=����[� ��4�fz�ۄ��@�hr�����/�����١x�#mn|V����J�F�_�V�e������Y�Aƀ��R�ꭿ!��[��.A	����8�j����7�{4g��`�|Q�2�1���V��ލwfJ��s����S�B@G/C��)��SO NZ҈���I�S�������¿�Ɵ�R��l��햴�頵Z]=d+��䄴}�Xr 4�4�j39���f8�|l.l�H�?++KF�E������a�lƶ�����&|˔��S����c��X������D-���;-n�5o��>��kէ(���ۿ�Wv�wə���������y��ۯ�,[�v�̻�?�-�>7kn��WD��O�q�w�{sz!��o��cc���v!c�۳ɓ��f�s�׃6��1!����������3�O纪��3T�{`�5�686�� [�tΆ[s��/�6��x�{�Sl� ��#9Z�㒎�(��Nޝ���AF��2���oi<�A�fL����<f�ƭ��@<�?�f�#ġ��:d�G���p��
ܳ��23N���N�X���Hҡ�[x�_��g��:���Bzp~��p`
K��}������;]��L�+���ErQrO�*���$�>��<Tnz���>u~�ߋ���	�9���3	�R'z�KO�\�5�Rm�+��Am�F���vf�����}�ǳ�+֗T6~wj:�BS15�zVjM <9��$��I�	���[�c,�2_u�4�4A���"Ao$D�|��A������a*_��@��Y��c�95~�6��S�VdW�y�1�ݻwG��)ޟ3�Y��U��Be�8�÷�n��6)C� 0i��@%���5��o�{��<�d}��URם)���H9.>>h9`�X�%��1��b��A̼�Ɠӥ��`�@=��A�bL����i�b����Cz[��E��%*�;�W�oR�Ȉ6��[�c�Q�2yDK!�ã1o���#P����M�,� k�NZ h~����)�b��DrmO�ORФ���"��<�;164��R�>�oUW}<~�B�FLR����U��D�V�?�z6} ���zw?<޲��ĩ�xh���jgc3����������H<��TZY
`�*I��R5�y�stL&�kI�@o�;-��$n�4��0p�߇ې?��ŏ]d���?<Y \O�����^(�R?��~GB<U�������.+�a#8�F8�?j�ꍊ�nW���_:��٥�� ��l�LN�t �ރ`���{^ �>�Jx;��X�zٲ�f�@ ��9W*;����TF<�h�tH.�T��~P']-���]޵{���?m�V�'���|�׈��DK���|*զ� ��-��d*�\�x���Κ'^E��v0����;�@U<��$�ba����i�<���p;"w;(��[:9�����=��`�IC��}ܑW8�]�[ekH�����y��cA��%�7��c�	�IW�צȰbU����siQ�y��'p���ì�jK	�a*�n�����*	�����>��}W1��8��f����3�>cWV�ؠ>��S/��~���:qa�Mϴ̼u�W�e��5���S!w�:�!�����J bM@ij����N�:P����YX:B���*�L�.����O_�O��_����0�!�Y�ϗ�3�T �0*"�V��U2��vk������E,XB2�z�'i�����pPY�|�(��4����w�bzIr;���
�m�e��Ȃ����o���v1۪0q�y+�?�w�Pl�/�
�Bc�@�tТ�k�<�3*��U���7*�=�9��E��e���/+p��a�!S1��!葳����'űG�Ӂ|��&u��=�q�x�m���h!Y���׊�y��4v����q��/Qm�k��M�%*���ȧ��,�?�^sB\�'�IC�h(�
?���Ug�n<L]\��v	uP���3�>gF�i��2s(?TgL���e�R���N�ŅP/�9:9�xЊC����ݠ�+KϢ�lڪ���v�G�)�����1	G��%y+yH!e��y~���{�Qah��F�2��i<�/x,U�Aax��C<8���T~�>�:;�jf�0�,KS�j�<6��H������I_r�]�#��r��,��
ߜ��'gi�c�����W1Z��-��CV�l��5���ב9��?Sk|>=Ĕ��m����'�QZ�s�W�N���D�V�c��'
y��Ɲ�C�Z���a��y���ઉ@���U��4�kщ��{��1�ˉJ��eh�У־��6�6�H�����z�6xGz�wLڲ���n���<z��q�qBn���?��_�ߊ\����M�#^���y��*�7-t������?u#]�Y(W�wE��m�Ч�q��\#py���!��ٿ7k��ƅ�|iKٍ~^plN�9H��h���.��2�X�٭��*�8ܸ�[(&̾'�4�VTG����sL�ɨ��.nN~�4QT�!�����.AܤyA����D,�pB�5�� �>���G�Ci���U�g:Q!��gW\�9̄0�?HB��75����>�N��Gc4xgdd$����%��{�,n�p%��ݮY�O?�M�R���/:}�5!֪Z�ڬ����v)��D��4yQ��;>h%N��&L��ͱ��iU�# ���	��YG��G-��sȐ������R�'�.PC����@02�j=d���1�_ l��(������4�
_ t,�Xb�Bz$�8Gi�G���p��p ��3���[�V��~�f����ZS%�%� ���-�i\�E1n�,���% >�r�Io��߽|��Wf�=�ߜ�&���"	ٜIү����/� ��!���3mՖB\o����8�Q�ￌ5�����j�Xc!�%
D�}C��g�Z=,�ۡ��9�0Ʌ�8+��fDk��a%��-.�����Zf�S�	��V����D&���yA�;,1��F[��	�]�j�<>�O=���yYA.^��Fi*�f�)�O�/N���B�0��$� �>��/t<�(3N�N����Y�s6yVU�t�(�lʢ3��2O�I�b���^dRls���`���

����q�<^w`��si{* 鍹H���B(q�����K�ֆ�]Ğ��7�<�ZI<e[�&H�h4;��ɂ�G
���B4�@@��Ķ�N���i�s�r�� �����C��l��y���R�?��!�^���x��j�~cjT
�u|�v�z_���E��N�4lI/H���cQ��� �7�^�t�"
��oD�!�{�w�U-�J��߃��.l�����\hR=S�������Z�CY��L��`7i�ݐ$�yNT���lvȸ�)~~󚠖�+R�h4��=\�Mq�@���
1+}���g
/�WGۥ�yKy��_���#�u�t����3���k�g�z/��R�K�gG�ڳjy}�
��K�$�����faq��8�K�9�h�3���0���DˬR]0�Ec���*��̧�D�퉉����@�F�	P���N�k����Ձ�������\�-��IO�0L�aL��Ϲi�S�_W_He��.�Jtۘ�5�Ih�(k�TTJC�#n�%Z��d�ME�%K�6.*7[��Y�V!�$ي�l���<����74u���^^����y.�<lk�H��XTPX8��E�c�g��J���%�`>!��lr�Ft^��;�����06�Mo_�3�É<�2.#����]쁊_��2�X����u�۶��*�Uz��޴Ƌ{~�-YK�����0яi����q[h�e�i_�˄� �ճ��#!?B-���=���ܖ"�g��^���Xp|����*����,�y�xs�[���ʚp�M�7��gcp	�/*,48�����@尧�n#��Y�~];������H�)���-@��N­�<s.���ӫ�a����2�����ʇ�@�KPW����PZn�l4MK�r������	��L!���m5��k~�~�
��rS:�y����k#�=���&f�u=��>e���)�Nˣ�|�{Q
(��e=t�ԉN鞅�@��>�Z�o?�^�9�*���T���0+{�e|t�OۓҲz6>D^>�E ̻���.3���y޻6~�1��¶��|y�	�j��l���/�z�b�E�Y�j�� �c��ƹ$�Ҟ�#�^Y�H�!����^]	՘*T<���M����KpTjR4������KrܾZ�Q͕�j�t�1a�ifQ+��!W¹�z�_�	�R4 1��ȟ����P�����=��Pot̴06T�aq6�UG��6`�:�e�gL,h���h�B�ql`ƫ�ɂP[ѹA�����ȋ�L�.f�՛ō�{"!R�#|/��v�6.Z��{N� aK��`�@��&�pN�Cbf}���X�Ӧs���I���T�/$���K���0�R��F0�/��@l��E�A&���	�4��x��B�0M���*�5��4E��ϸ��<��Q��x���R�?=V'l��\y.������v�"[�����9ek4��[3����ω�[`h8�o(z���0@AĿ�_:��U���Y��R��?����ӡ������Ń>�/�x�4Jҝ(j��ɑ�trpw�����s���\����r.}�]y�6#*�(�Af���:f3QT����w���`�C��6�LS�ZA�1T�y��[��*��YE5i������)\YS���D%�e��ۺ�P��uP:�ATZVؼ�N�v��Ox́e������� �;B�Ȅt��l`�0���Q_{^2'N����r�f#�?��!M�E��?�;g�gf}>�ڻ�ZS�Y���qD� k���;E�|��Y�0(zx6�B�j]pd�aAUʣ�R�.��u�Dx�"o,��	y�2�(N��<Wϩ1iii٧�1�����@�Yxv�J[E�#H�w�25���(L�u��\q���y{N��*F����t�S�2T��/H�o�`�"�O���h���bm�)�V�유�#���k�az766����8��E�<�R��|��7w����c3�ǤD��1e��=�����x��ó@v?��4�'��w�,Z(�bF���C��Eҷ
����@��K�>��Wb��T$�'��@R���Z��k��A�K�r�O��?�J��x5��/E�G���������e�|��>���'EϘ�'���5ϲm<xz-��+"D+���jyuX7�̨�Pm�����^���n�g��L�F0�h񱆧���]�&����9���ÿeH�g�[1�$۝��e[� >�aQ��2����Ξ��U������n"�8�m��ԙ�&r�u�_�D6�Јe����e�Y�,4>�{�#!`�	s^���/:�R�ڒ�h<6�?�����>+\{͠lQ>6��]��B;q{?��Y3��oĚ��IG�Z�kDF�D�n��Y�:xz��:��=W�}Wh��Ȧ
���Hw��`?d!��>�P2F}�/M��5�������^���������q�@��LU��Y���{;�U Z��-���ϸ.ۤ1o^�X���n��b�s�Tt�'��z�������lll�f��HU| B��O_#< �-����J����r|Θ8�Pn/�����.k��-H�~��$uN�LJE�q�N��׎"Spu��o%���l&�{����H_����������#�����Y��ȏ��o2��$q�#�i[p������duG��yK�l1�K�Q(sB-�Z$�����m��	�g��o�����d�p�Ź�3��p�<�ڜ�18h�f�V\~%�Β������|�{��p�v��E�2��ϼ S� ����By�~~mI<X��E���QFd�b�T0'���8����Z��y%�ګ��_�JG#��
��.�/��o�;w�oh5�ҡ��v%6ݩUh�B!s��eއ�
$�:l����EP� �Zs��%��24ϵ�s{F��=�T�J6�z��-ڊ�,3����ƛa��71��c ���/'�ߕ��F8셥���H��Qm��#˿���-N��IPg��N��b���ps
�x Q)���;A�-q"�)T�7�c� M���� �5���.�`a[��@|�)>'h�nB��<����l�Q�'m�{i`��I>�b>c���h:�2�1�42Z�ck)\	 {y�-W�Ù�����C�č��u��$�����A�Z"�!�W���.��?��v���X���
i�:���#���ɾp�9xB����m���)?�+���2�.���"���q���O��ρ��@�j�QQ �w���w^f�F�1��%�Z���1}9�r(�*�6�SsU��j��&��32D�5�O������նB\TN�t{f���������H�幝� ټ��^�o��@�Tn�rMp7����!-�|Po87���1o�0�ʹ�����i�h��zL�$�������U�5���>��r��_E��0���뀹S����p,�@[�8��`�F�k������u?;�1^9��$���,�rn#0ׂ+��[���~_L>����RR:�e|��r'o������&�w�3��"祑Ac����6�2"-��E�rJ��^�dmy���6�	�q�4#.��0g��T��w�T��DmF�Φ萊m��N� �2-]�gN"��3�s�en��\1��GW�ɶ!p۵���#'�K1^�,�c56�dD��?1��&&�,����'�jj�~�}�i�N6iT?nC�Z�Ŗs�3@V�P���G��`�{��FS�v���^�0+�p��z)w�<t����}�˔ҾwB�ʖ�;��M�e1���_Y�{�R��ޞZ�ϩ�����U�ډp�Ox�Q��ʭ���.@�}s�98�8�������g���L�L��cC]�à��k4�h��g�V���Z7#�%���&�,K���[��r�2��Ŝ(�Iac1������m���d��kF?7�{)��e掌~���u#�w����9:��yی�;�'�J ̗y/)����P�"���%�E�@�n��]�p��<�a����7�f����⥷o߮4S�0���F ���� ��cQ�`wg�
}���&A����Ɍ�hj9؍IfT���n8zp�*�J� ��N���٨�}��e�i۱k��ك�+}�y(m�2�q�rb���,���C���]�=�ntZ|P���y4�lfrk�2I�rl�lC�H�tk�7�����3�����Ns��������'Aw�^H��"V ��0׳�d�"��Arr�.�>�p%��e��\���@���W�
�O(�k��Z2�ցxl��7�� D�T��������{�&&/��N"l$+&� �wx��P�(厅�x"�:�14)�V���R�X !�*�ޫУ:9��կ���*�@w�7N���DG%����j�-�\�g�z�I1~F��,�h�&����s�F�n3;�od���}/�A�Ý����ѥ�>~\g�s|I�A��އ454���{�����Iw���� ��|(Cޘ~���jF;��Tĝ�&p�Z,~3�F�����]&ׇ>�����ɵ���A�Ѷ�5û �`i����2o��>zh�&<���.Y�)@��Q�H�Z�5~�4DiO����~��/�Ʈ�%�
�$���.y�7�<����}=;�
0�?������c��C[��S
�qOW��'��M�H�����O�A�@-S��������~�1E����&N���/��郕�u���>�9�����Cӕ��	dv�T���bOUgc!c�4�#u�+�Y�����>�gT�O����
��hL��~�D��B`� $��L���{{�a{&���C��ں�������;��Y��� �8�q"�bC���{��Ӊu��1��cb'��E���U1�����,�k��~A�*��V>�1��]�.�V�������,Y4���R1VVV���U�̉�b���x��n���_�Hr~��FZC�ت6�%Sg��Y����4X�|U��{|æ�;�bmh���A�_�C~wȯ`�Z�DM�(����
��$�"���eA��\&�0t���En����X�)BM͖���O�#�����{�P}af�.��d�lJ�1�k�733�`bi�,di'F�� wHbj� �1�Ȉ[^gg�$�"]s�"c�AW�pO̞��3�/�B�g�ָ��v3��౥V~G8��6ُfc����%�v���� ��$���UL"��i�I��sil(�9�}?D��Y����6�ĩH`6T$�����.�G�-ѐߊ���Ƹ�y�>l;�f)�¼��������`|�nE�fy����[���ݘ<s{��,�vK3{�S�Wf��s|]]a�����3H�&�Ճ @hxs/X�I�n>�d�dx{�OF���G�ռ��70]�1g�occm�rk����Y1�Ƹ��_y�X^b"5͠v^Ù��m�2'M�59q��q�dV��1�ŕ+ޫ
2���Fg�7]���#W"�;������dD3� �X�m ZӕUPP�
��:�$�_�����в�Nּ�q�Y��:4��Gׅ�&*���{��e�6Jʁǻo��unb+|��	�>��|��滎V��h��m�9��!�$H���i|5��?�Lp��Ŕ���oX�,I�0ҝ�|�u4�u��3{<
��y�x�&_K�D���g���53T�}�� !ڇ����v�OA&,�(���ڌLX�􄙩%:"�2�PQ�=5�\��t�
J�Μ9Sq9�C��q�'Y��Qm�>�O��o�^?56٭�v]���30���ߺ��d���H�ښ�
G�+�I\g�����m�8�����'�O"kr��M�V�Uܾ&��22k-du?6���.!�N]�[z��z	p�5��+|)r=�����$Ȍ��c�j�%8���%�̇ �Ug�4�ϙ�d�T����{�z�=Q��� �� �u�<�(�_�e���_+���k�X�D�a�W����p�zS�� G�k�I�V�ЯM[M��t��=;a�!�a����[*`���.�<9��e�ߊd�6œ����J��`�����o��Nx��{�i� �Ƒ�S�����>PzE�����@����Z:;X����y�Mh�cC�3�<IU%s��\[�ܫ0S��ǆZD���:���d��>��n��H��uN�d�x�S\!�^I�9����N��'�"���@��I���p��[�S�&
��̹���㔦�(�9���4�}�b��dY���nUTzHxK��!I�Xz�Y�(o=�d�G�bC� 5�k�pW��ᡞ�G���h�K��M��R�L�K-��)�3%]`�*��5%Z�CD��|}e��y�  �n±��F�O�g��|ힿ����*Ycl<���mU?'6Ey�B���>�&�CR6-}2����O#�++ܬRq1j%k�F��+P�;�I1S��c
�ptf�aV���#����y��R5�3�am
�����N��6�H
�4VcB-��43���E��[Vd�K�w�:���g���mJ4���T��w"V�9$��J�|S5��F��%�>�-�e��Bm��h|��O���s[0@Wr7VMF��Y�_�0{ݕD��b �w���׵ �v�Z}�n��� ��Ԅ���?��	o������$?ɷ��
�:��<���;�g�=�2V�����RI�{	�T����e�� bH���(���^��|����_i'�q0�; �?�/��:��m��\��;0��{���$�����p���$�7{I��'�yr�W�:\�j�����E�p���!���VvS$E�<��/���~Ho�!�B��x��oZ���bB����=8���'��*J�w���J��i�G��/DJ�9��'U@|�<@nw���:�y�kT���'ڃ�*߼�r�rg���KTkZ��){�b�z�@�<�������V�q� V�i��7���\}[4�� (���I�/�ī�*�LՔ5q�ːgs�D�T�-��k�aο<�����i�^��_8Ġ_�3	�{��D�?M�Q=W�������vz"��*{2�B���{�ĢPs�����Ţ���׸�f0Ku����1y�� z�����SЖ�w�<@����Y@�����éTKvx��$�0(F�GP"K�c��-48O���Wb�#CfŔ��ٺR������h�g�����M8�W#���GV�����gr!E�QIT!����fa>�05� ��<V�%!Ë��1U���6��ʾ�︫�?����?�%*�2O�ؕf���0>�>����j�Zr�k��;09��P�4)�)�㻡�s�I��Z�P���� Z�,�����͇n�v��>���:n�zS&�ۏ��bm�y��d��T���т���ڜ�u����=A*�C��VRU�t3�O������OkH�b���$�^>+1�/	���g�g�kGn0"��U]�o߾�S��gЄI�^�k{���7�_�%�ۍ�^�QwJ{F�~��
Ӕ�L��
z��c�0��W��-Ga}�:P�_ȉ��X��9S�)JA��Q�=Gđ���^�/�܊�+�":L��ߓ$�=�5=ˑU;�E;K�ӌ>gB�8SQrO��Y�܊ �!������EF��eD�8�@i��!ĺ=,#f�X���0���� ���Ao�8�KcD���X��Jp�1�̻�������@(˥I�^�/�َ��ѕ
'�1��ؽg�n�K���GD���:�B�ǻ_N>����:r���N �<���i��� �i�H9�r.�Zңw�t�n[��M@��8��JVY���%�6d��W�,9_���Xb�_3��{~�k���LW*����st;��F⅚���k4b]Ma�"ޙ�%>�ņ
��S�$��� $RkP���K�m|�ګ�638��RP�2 .1B�ї'e��f��&���))}��z?%2?� fQ��jH�1h��M��?�'n�;ۥI�/Ò�y8�E����|/�Gx�<t�B���&�"����j~�����7���X��8�Z�8�h�Z�/��6���gN� 櫋�1\�-�F�{9��Y��|P\y�4Ni%(KL%�a��z�߿�S嚾�C9�7(�OA�Џ����&�r'�#RM��eYܦ�����b���+���E���-�����d����	���q������p�����Hx�=G��]����M���R�W��j
�v�;<�����/�&�ܶ�8!z�w����}����ܖ{��Ls�{�:P���������v?�R���,k)��2Å��T��g�u_�t��",������"kM�����|��YI�t�dPm����C:�c�&�L��/���jTg9PL��K;�� ���Ã�Haq:u�:�:9Aw
Z�V��>�m���ȵ�w�
���(���������������Z�ݓ�V��t�C�:ekk��Ə}���=� �F�`uģ���,@6��R���s�3�@��|�Ze\_�Ѹ��9�2�(.$|���H�>.�Yz�]�r>�\�̖~(2�{�l�����n���@�ť'<������w�"���[-Y�e�����'KA��Mv��F��9��K�����l��s��{,-�2r!i��%˫o�X��0M��{4fTD�S��"�_�8űJ�?�K�h?=�k_�y(�;��ŷI�'��V:,#N}�)�h�<�Q�MbF�"�>|zu}����+g�O	���'ƴ�򗁮��a�Ѧ����|���!�Zc>���߁�L��Pufd�6�r��w��";~���ل����	#Y��y��/s�GLC5�)9Lb~Agp���c��6����;������w��j�=*�>�d���Y���Wn�O����VY��՟��j9����2��NMP0U�ҚrОi�h� �4Z��tF0|����uU1�����L��{((�yr�3��G�?��4#6�����`�Xk�b�⍙֢��g���DIr��G�'	��b	x�{�����=���MO8� �)���r�p��R�C��_o~tѰ�-%G�_���U1��U�����_�ۙ<kD�r���">����-X�ꘙ����0#
�q} �I��$�Ee�s�"���l��&fE�.X���b��4���񧃥�˵E���u��@)�E!���C�����ڪm��������������V�̞���}Oɶvѿ"&-H�l�U*��o���)\H�פ���mM"d|��0R�ׇ�C����`�����J�4��V-�=��p6K9>	i S��B Y�7�B�.�H}�t�ݗ�hʂ���4 �����6���
e=���ڪX�H��}oIǬF��dҨg�)��4&��F�q�׻���)�+`k<!͋I�L����ϖxws���B��ST��8\���w��w��"o%e�*�j@d8Toh�5]�b�'��E'�~4s$�[#i|���*���f$K5g�c�%����2��^i\�s��>3���O���A�&��)�	�G�X6O�}Q6kl�S�������",���J)����%
�vW��ʀ\F�{0P8�Xl����uHȍ��׽�7R#�h����`x��,@��B
P.;!��&��Sj��4����u��0�'����L�2H=铇*C�� �ar��4u��@n��'�H���Mxh�^U��ta�wsų�0��L�Z���vJ�������j�be�̴�ͯ'0]�7gQ�_�=	��^�%�b�ԩ>(��V��T[���8+���{�`�3�Gə�n�"D`@$��ɪ�#Q9�tΓ걤!����� �\ȷH� W�*F~�΂`L�M";�}ж/��m�^hs*��:OTUM�$�I��_�U���^�D3�a���p��j��1B�fK��\uF�'��]��@����D����R����+	�5+�3t����.�� �s�Z����(1n�sbK�瘂�&�`�A]k������Bs|{�}{6�5j�A���W�f�^Pk>a�&m?�S�C��Y�Q��9��}��d�A��o�_�b�.��k�fKuY��d�+n�D�,u�Aj7!Q 	���)�����T����z�8&����J�m�]�4������ '#��jϟLg����NQ�M�D�f�8"��r�9Ԛ�]����Ey:*=���������j�Q�gj������/.� ow�� �`�&���/7>.�Wu��IjQ�g�=��x�U�c#Fǔ�k'�(���ꯗ�2����10�6���H�*�gV�v(U�,98��br����������Ak�]	��.�j��>B�z%%甿���$�ȑE�P�C��bӲTlz\�6I�Q�?`���ŋ"~'^��:�4�ne.㳁qy���c���݈����@Wel�;:�cz����1��٢������;��?A3�y�����3����?����?b:��%D�Z��	�`��7�E�d�� �U17ZTjg�RT#�\��5�b�vm_z&L��z����u�H	����Q&�kK�xͤ�ƨ��$�#�	R�J�M"����.4���i �bK��9P9�4�?⩖�&�~����}�d�~|^���T+�:���P J}y��Z��]�r�C^ʰP�ː�o�c6yq�b7���-��,�ӴÏO�pl^���Va2�-.�bp����=����H��-��Q�l�&�^�d{8&t?-W�  �S��P*@��"ʓQ�Ǯ4� Ғ�FWYʝ���y)�G�_�t@r	Y�s
߼@ok\T���HT����*
��4�쨽��1�qANᆭ��$��S��A���,xq�'8�\)����ϐ�����`,]�̠��M�Ao3���7 �猱��XsA���;���T�5},�1����!��q���Df�2���o_��0�~�h#�w4\�q��J6F�Y5�n�煦)�8ʝ%ZL~�$*��{ [�?\Z>��4ŷzeud�{̤��f�v4�vU�fc<��]{�ؘ^bϳ��N#r��t�WJ���R�j#"""��ɨ��(���o޾��?���[m�A�@���fF��!r�	BF����o�Z���M�U2a�:l1��B���S2����ϱ�P���Z0w�M�$,���Z|D�%�tQ����I���jk�|�7#@�$�+ry�j�巚(n6f6�w)J�/ Z���W�4�Z�NX)K�g�ȡ�H�k8��r��A��u�=��Ak��HU����J���̫�6��܎0g�S`Ο(̯i�Y��ȏ���~1�̜>~4ո�бP�P���4��ω��D�Vg�8�}��� l)i���dm�=ķ��U�v�D��?k,���c7K2��6ˢ<_iɶo�Y�e�+�]]��.���EQ��4����x����yH��� ����{��b���6�Q�
�+Ry)��\��g
L������:� ��j�T�'�z�0���Q�$�%+?cFD��㉉Ë8� ��/�� !�ZS6���ͤ����.yҎ��v|$3:�B�~�z,e88��%�]��=	I��Tw(Ax�ʖb^�����v��R���C�N��A�6��uy�X"J5��dj@�e�s�8�9�<�����q�玀��3�	��T<�K��׉֚�̮��cg.)J�a����}��"���y�:�ʭZ��|e+��$)3sЕ��4 �,H��A♘``b�R��	���ÃKO%�f�pG�?(K��_*d F�o��
���ۻ��b�h��ہ���$IO��um$D��� �+�I�bŻm�u���-^]5��4�SGv�J+Ief<�������`D���#L�޾�]<��d@�\z�����'
�D����krVȓn���Pk�Qk�oy�v�ECq��c,��fe"O/�F���6`:�?��BF�S��@:�h��	�)i:��̝�MsMv�ȓ���\sAf+��Xҋ�,��.�R����:�%��!����h?]wKŒ"&�iM�j�"�:싊��F�;&�H��OG�}���� �����S���L�yc�T��=��X���������uؔk4;H
��%�^�� 4u���8����|�T��Hbr�1oR�$����.��7FF0��M[*vӆ�׻��FH\�F#U�Q�Q-��<.	�Z@��9:��	�$9-��Gw��nPV���Ri���u�S��v���x���ہ�?]ʖ _��s�'tku����Z'����Ay���Q�[w���a�{��B��A�:��~L�mU�p����Ǭ�S�V}�$��9�cH ��E�ofX*�wF�"C�ן���������K��� \T,SNnM�J��ĪLp%΂E���1i�cI��s�)���?=��_�z|8Z� [>���鱗�X�T��Ly���(�¥;��|a��v�P;���<�^������[�g,����-�<��{!�#r0�%:�#��Y���g�Щ@Ѿ��.E�hܔZ��#��<8a��F������Ж�$Z��*S���Y|v�_z��ւ�q'�S�yA�:o/"l��RO�q{��{4 �r��Ch�D�6����v�%{��e�I�>BC�����i����P9�عRK`�֣� 	��d��(�o�V�;2`_���a��M��6��J&��OEj@I�f*Rq��B�sΥ"��.�D�p�hP2e���h������/�u�=�OS�HMXYIϣ�*vF���q���Y�,]+{�2{0��s�+���|�:�*� h2����[����X�OR��b��+�����o��a���7����������Zs��M�����oT���ͫW��p�Ȃ̯#��jZ���=��܅�A�G@�7�=|I_�(�(�G7�]��n���:�]ڜ��v�-�I�R����k���zJ4�t�<�o?ޣ���A֯�N�j	w�����"�s8uݭ��c��l��̾gg�)#�grl���ڑ�/�	�3O��s�����4��ȣ݆���gb�~,mά��NI+
(9�k�GFU�T���X1A�X���~�1��~?�"3�$K��t�a��Eц�)�h�T���ʿ���N��J�� bn��'tՆ>/E2�9�+�D�gf�^�;Ej�TI#��j\~���ٻ� u΃�� �3��s(���Tte��	q���m{�L$~��ɰ�ĝ�����]��_N��������+��n�4:�?��$ك�#a����$w.�R�a���/q�9��n�}��M8�=&���1V[~�;=3ӭw���.��
��W�`�NI3�W�������c�7#/f?���i��5�U�� �/������e$�����E�W��%��T�?�R�2������۷���w�c:"�(�|��V#�V)���8¥#3 c=;|_r�����P]�H� j������#2`q8��4umf���r�v%�&��}�h���Wf�U�R��퇕�.U\��>��|NQQ��
�S2�����N=��朊�v�<��~aJ�k��O������������&x����9db�m�bF���*$��Q��ޑ#��w!����� �ҝ�e�+�$�� �6�U=�}��*���> ��k=�m�Ce��y�@c�J	C�2�	�o�^��$�Â�1׾1Tbk��H�|���#)�����ho�cY��E��M)�y(��}�(#�J�q�*�.��8����;H�u����/��¡%G�Xa��ao����(��~�|��mv?�~�̎B��¥��\t:-�B0B�{�b�mLIF�w%�������AM���?"%^���ft����MT����cT1B��*gh)��9m�Y/�xD�Ey�;6����Bj=�ֳ�������$��V�������1�)!�g��#r�8�4T֧��O�.��"�H�
���4��e��VH��q�o}]M]�=���q�3�ԣf���䤀���l��56�|:��&��>�н��UH����bÄ��̜�ߙ�:8k|܏N���L/k�3��b�sM��1cX/R��T= "���
��ɱ�d���#�E������c�˫	:tp�z��,������_lX�!at���s=p�>j$���J��Gn�jG��ʶ�|늲����;O>�z���rdcY��'�Q�]L������y�6�o�5/[�(2�x�+E�=�D�h��eS�5g�R^{F�|�"�2ע��Ȝ�׸?��ߌ�1�C�,Ayu6k�ۍ)��,���z ����R�06��w:)�:y��EHB꿌&�}Y1!f�1ğ�P��ђ������ʒ�o���`������4��o�3�
���^��8����PK   t~�X'�%( �J /   images/6b7f4d85-4146-49af-b1bc-6149946ceff8.png�{eWA�' ��n����	�`�=���!���!����� �w���������9s����o�����PeEiTd"dTY�/00+00���!�tJa�?ɪ��w&!�g$;�o�00���/�nsկ���N��N_m͜���0`0��������Δ���{�p&rY	1U���U������5��F�v�Cl��6%����;zk29��-�<ֻ��	q��@A�������UVWe�u�n/vi��If��4��H��?�3CG2V��d4}������	��	����AiЕ�����7`��m�/��&;D�-��hWB��T�#@�-cߥ����%�����a�Z�o�<�0��Y!���"G�3����,����]� ���7�2o����*����j+��I
b�n�\����݄ňaK�Z��nEGt�A���o�< GY"����Cmy��ߙ���"��M@x)����1R��U�?�}"�a5���i�1�'_��bA�[���~�W�����V�Y?�͉-��K>r��l�EfA�_��q�E��4�/7���
3ݹ݅����bM�>娋���dLC/��a:c|�4``6� g�����]����V��ֽ����v�뻉���������ވ�����_�hnO9�-a���q�w�R4����[�ǝ�k*%����y"1A���里�~��/�#�C��ڷ�_���d_��G�+����FA�{���?�i�_#p���'RI7�O"�L}xa㤢�9�1�v���vvS^ޔ��u��my�J�ߎ}�:�3>��dAt����Ȭ:R�+YRq�66�e�ie�zC�z��0�9�H7�
N����h�Yf�4���@���2tVb�@�+���:�ӊD�R �F��\B�Vi��M�9��1U�����X��k!T=��j=���,4�մH���Q�P8�H`5�Nw����8V?:�S�D�����N������f�>ߌ?�?�:k�kI�νc���� r|p(w�`���Q������6�[ֽT:a��>��u��s��|x�Ps�}���J�ku2asS����jv;I(�{���ԑ7�o���p��A�L��T�Ke3���2⊿.�--�m���f	��M�ވ)��D�o;�y*�w��Q����j������yRm����x���������6*Ph1����t��n���|cr:RT�g,1��@�ܬ ���������F�Q�a�y��j�R\�*==𓬎{��&fxN)^{���q��P<�3�cj9{�-;�^i�f�ݠ�.�JO�x0������q'I�G�c��a�XAe��y�+��T�v!!��&9����̂� ( �;"(
r��7�E���ѽF���~u��|�1��ns�!��ف����t�9ﯵ=$����ș�{m
I�\�V -��ZA�O�z�AZ�D9��3n�hmeLFt��@�)ү�S9gͣ��&����r���i�+~̀�H�pl�/M�F�bI�����Aݏe��@��L�����)�e*�兄u�8a+�������a)x������x/,D�/�^-�΀+�P�`3hW�FŇY�$�!͒�ּ��+�Gu����uOqEG��(D IԈ���.t�9�뜻�q��w}�*%���mk�E���7�!���3���#� ��\j���7�)� ��сN7�m�s���2���A���i��S��ޯ�-YI���`#?jAZz�<s�_��~����'U�-0�b2о���Xk�!Pe㓖��N��&V]Z}�_���	����{,�M�E���T_5�E���Q�0!7s�t.a�ݱ���X+\������m�U������P�9���D����*��Ʉ'P�P�"��l���!6�rƪ�m4Z�K��P^�a!e��J筞�V�ϖ�B8��su&[�K�5#��3�����\L��d���T�YfI�e����'����8���</Y ��5ľ��2���n^��	P ��e��"�1�c���(lAL�⋰"sԄ��Lt~
)��"� }I���*d�4a���cm�'�u0f�տ�j���`����A����V)�-�P<b��Xuj���.�Ë�8S �sF�#���@gf�W�5bx_s��/:�;
3b��u�nL�,s0TKB���#4����T��!!&�\��s);���kp���D�R�>����U�5��C���0�;��o����b���Ci�7{��x)�7c�R겄��Z������UėH7�Š�$�O'�����d_�ZAT�5�]S�#��)2��6�-[�p�-�g08�7��y��E�7�B[CT���s��K���Xϳ���Py} �I��yߋ�?�>($��u_qZ���m�Jր��#l������ώ:�Z���u�Ƶ�Z`�֕���{ c�@r�H~�@֞B���RV�� �ӱ�`���H����뻄�����ܫ_�6�G8�0𣗂��P�������u[W������ִk���Ae��3��Yɬy_8q����N�T���G�OO�r��5uK]#
��څn�D���!�a�2��`-�(fu��Xtnk�L-�2^H�|oÁ�ѥK�$E�!k~��t�V�e�-ڟb3�`7pE_w= ��q~x�����j/�CI9	��%ݍ^���a��;�uw��2o�(�����|�Z$�p��&F�rG��(���֎`�x! � �˧����#Ϡ�[�;^N-�����P�F5��^��SR�RE��{�ӡ�V6J���t՚��U�AR3��D-UE(ڂ��
�i���7��$t��?��*��u��^��K����	>x�]�*��No���Y����`.��]�WY�0R�ޠgs̰^�ʰ[�X�$�J�e�G���
��Y�j��{�q_����Jh�ߌ����@VN�����>�� ����;�4#����ۍW���0R�:s��㮭���)���IT*�b��ﻌ�X'%���Ri��^o2B�=�"&ms������2v�n�T�޹�u����~4�I��`Igaz�S�.���T�7�\��#�9��~�ϫ��\(��+a�p�R׽R���+��'+��J\�Jt�GƟ1j�����.�?�N�A��T��]A���UF�S��K�f��da`^-#P�lT��&�I!8ϛl�k����B,L�����;6v���UR�݋��-W:���_u�-���a�1Iaw���M��`��y����{���՞?Yc����H��5�Sh��G�=B��a7�4�n�>ӎ�������`�6����ϧ��)��)�
�K;zk�)}�t]�y|�0��#����Ue�k�\���,X� �77�P�f���E\�lvw
Eh
�L�yC� #ye#?�;WYlR70�7�6Z0�z��6���~<��E��AWU�x�m�a7�`g0�[�^]��/X_�ldN�<��r��XN���BYl����BB��D�A�ehL����ˉʐ� �7�"J�>�
;^լk}�
�i����m%�Yː���`(;aa����t۟��������g|�zoXYWY��L6�xJei8�Ǧ����F�QE�1F5X@j�r�Y��w'�l*�B ~�����T[�^�	L��Lۊ�8F&4N�����q�<t.�5�%N�9���j�;�g0�2��_��Ni�l�$4�r�����lʍ9�h�𷦖�"��o�ӿ\���]�8�G �k�j����ځ*~ ��:�f6R���J��R��e��(��b���Z"�-r+B�e~*����g�W�d��-��TY����φj��a�#�6��Q���!��_�������/�h��*��B��I�#[IH�Y���g�Z�a�� u4٫ۥ[��9wΈ��H	���*�L�/0>�D_�>��K�Fq�p}t�f�'�����֘�1���|}wzvn�YS�$j{lBS���E�hf�ud�(#�
U���?,���LD
P����yƒ �*���7S�j �i���&χ421n\�
�k��]�y�O��ŁhI�R�;�'֐g#Z#a���W �v�_��vh�Ǌ�7�0�Gr��گ4p��%X�J�F�[�c�7��N��''���)g�?0�w�]Oq��e�f�e�BQ�U�zj�x�[�p{�ȣB�%@S^C�DU�� �ь�ų�����WWHB�4��6^�ɉ�[!�#��,Y�4�oh��.�*��m �(�1��7�/�-�c �ȋ�,8�����!���������EI�,,����Z���c���[��=�غ=�B ��e	��I�\
#lTp���fC�zL�q�}�w=�:t�X^�,^��
�\rK�^��`������+������%ud�Ō�&O���sQ�PD!R��D�x�<��G�H�9�ε�� |$p�X4?�Y�fm�%]3������7�O�,�c�M��Q?��ԗ>��!���z���qut��������fZ^�'�w��b���sT1\
�&:e �vH���������v�`yNT�yIQ�)�J��ƈ��~�6�9Y+����3^#Z�O�Pm����Eg* ����n���2�ߪo�]h�Q����&F�Q�����ek������9@�q���������F
칟��7���ӽu#��,o�^�ê���@vEU����(��t��Ԥ�nV��l�#�j8u�G��aQɽi�4"���@��OC�!)JŪpel�H�������(�X��Ad�-5�\��H���63������i�ѱ�E$EGf���R#���P	��4ڒ������+�^%T7`�UT�S4lH���w�`*�����-�Et�P������*E�W"��+2��1.(�v���J��×�ᵒ!	��2v�Az��ϗ%������'T�"EM^��jA�η���������`�cw�t�F4Z=�K�����kf�q����	1�J<{����W�e����?z����(�뾃Fc���Su���s*ߍ+J���l��������o�-�-�N˯�k[�$��RJ���f�
[�h�F"o'o��8�J�`O 7{X�*D��k��U�եZEG$�_̓F7<*:����BC����QZ(��u$p�α�^f�Jl����C�&�I�Ka��Dj>��E=� f��X2w��*i�m)��4��/�$�Т!>�P�{cN��E��ɇhU��g��KN��D�r�b=f����� ��'S���ҀɊ�:�د$��=� ���@Q���B�f�G���H�"�h�������%:�+�uia1߃*!�VZ�Η��5)돩������*��PvD�|l(��[�qM���Y�c�j���+�����}�oP,&&�Y!�zM�����Y��5n4�ҡ����Φiʿ�;'��ƒ_�VcB�9�]��BSxh���?�a�h��>:��
�D:{ok����'��ĵ��R�>0|HG*�
VA������{Ϊu�P�����w�����C�c;c6:���<��߶��$*�5��X�u��rĺ��u����y�� C�-�v�v�����o���Ւ�:.@���D镋A��Y�H ��/w�������봱Ǵ��ڣ�i����~�|����,vE�d�Y]W��1Y!8��g�̧"Z>ҴFn�������H�	( �L�L��kK/��m��eU�Ë$�޽;[��vk�}�C+u�[qk��+���8ڢ�V���������#�Ep-�o��SCi���LX-��p��z�+�h�z���IW���s�
 �X��	_�4�e���/�s�j�Ļ����Q�3;�;�3�U�ճo���BD�����"�\�kM�6�����D�{��i31�������U]�.S5y ���J��x��3�����஼�8T�+�8-�QM�ܹ��/��O�-><,�.�W[���Y	�^	�JIΑഥ}�X��X+���l����gь����_1r8zTzG�*6�Y��?O��F<y|:�����S]�%���(��gK��O��.�V*I�MM�ܣ�/��j��PE��I}��}t\\����!a���4?͙bLU�`;�]_�6����q%�Џ�d���ŵT^��p���qDW�g_|�8E��&d�f�	���4B���b��S@���m��r�vm�\���@�/*{ҽ���j+mnA7��ob�N���5��F�zи���uMa���DsG����q��N���s�!6&&*^#�
�3��i�*liE���t��>~���}�+�O�����h�x�s�W-����tZm���=&]O��U���:�G��A>�BI��[�tґU.O:&ǉ��ˏ����:�CmHJ��,�7� ��bzs`�-� �6��>;ɫ"��m&- �-�~o1���:X
���_u�!{�1JR�	�%�C�-���H�#<snF5X�{��9�fX�G���n ��o{ܑ)��J�Z(��<,��S�	&���ʵ.�ce5T�n�s��Sd�+�=<�\Kz��ۇLn0d'�A���;h[�:]�f���0"����9��x����R����w�0$Oz����h��������7�Y�"zZ^:���y�O�JV6w�Vx��k8@v��-�꿻���x]s�g�=S���Y��R8`�n�>�:�œ���PŸ^V]"6�Ow�.J�p���Ӊ,Fމ�B���z�3Gx:<R�_�����9�O��r��^��0~��3�pR3��V����*�?$��4���H���e%)�!U *O�7����*0���(H��FNj��ݴ&���sGN1�探�����,�|�0HJ��Ō���%I%�c�����$���u�`�S���f�d�\k�$8�K�^K(����-Bs�W�3a�a�\���/$G6��<�څ���H�j�4@�|���B�/x_j>���4�&�����[�ͩ���I��/a��L����^ER<�]r��!	���j���}I~��r��~v۪1
_�c�o�5q]����.�JA]�PDfnh�{��$p��7����a3���Vd�r�b8a��&����|T�[�UW?�*�3�z4g�hN��h)b����h���s�B���5���0?e9��*-�	�Ƀ�����r&�鹷vK3���*,,�I�I����A��2BB~��Z�S�n]1�YX�r�4$���j4Ɯ���K#���U���������9�^_�Ǵǈ�-wF!�'�r�Gd��+T�V���ߡ�eYݻy��A��ɽ��݇fz�o�O��緬u�J�nʯUf����N!k���5�K��Y���~�1��֍��A=��<�߸�I���a)vJ:7X�E�����į��a�u靐�I���l�A6�g��#ϲ�I_�Ɍ�B['E�/��X�J�g,#����Mw=JY�9M��2[�y'e��a�l����|(�y��1i���J��	}n��r5����"��_�[q���X��n,.�>���[)Rٞ��*S1[��_�����-ɱ--�R���ʕ�mx\U��ś���H�0:�bgn����֢1��]�IxJ]�kQ���2��\S�X�{�Y�H���t�X!j�<�ȭ:EtD,���V��r�~�T��Z�Ͻ O�]_�}����Mj,Թ.a�����QYh(��y�!+�}��;�b��B��|\}�z0%e\/ �ӕ�}��i�{�fc��:��'1BI?��6�����~��]�6������H�w8�O�%)�����S��� /�h���c��[���ߟ��5�Ѻ�_�*�4h����Q�����݄�>ݠ�x�2�M�m�ɮ����i�>��e�̜��w_�Y�n���|��h�X�yk5"�&�3*�8i�9�&�@(b��sz�v��{�����k6K���I��n�4�c������S{6jL��@:����z�^����'�g���NJ�x0���Ϟh�����B�ⷭ�r� #��Ϭ�LE�t~� =*}e�o����b�B��1����;�V��u�j��e�bsq��O�������=���-�]���Rw���9�y������Z|��d0�Үs�Ren��^��<����^^��	���<u���G�*wW�ם���nk,��{4>�'2�5�H�@)�SWi��0�N|&���~���!��{���_� 5G��u�14w�pX]m"�?S�~*T��M�q~��8``4gb�c�<2ޤ�4$����o��X�J�m+ԣ<����޳x���b���X�U�:���x��e�#�.��hn�	��\�� ���;�����yS���}_N���&"�$�k�����(&)��}q˘�~�~_����aGf��~��i�(��>�%Yv0�q���o�]��ZMldS](O�$��.�J����'�~�/������L����Of�IO�^�n��/�@T�a�����0G��?����!�T�WC+��8�y�!���e��Y�z*�q-����8�[���ɔ-�Ui�	*X�.LH�u����%�r�'�x����6��yj�u�ˍǆ�SR�l\�2kaɟ�߶�	��չ���wc�Y{�˭��RU3�lGSC�ǉ��j_6U�'���,j�e���v�l�( n���w���)�Q�8ǻ���C'���Wԟ��9����sEK��y�����g�R�Dv�Vݲ�Pz4�ڣf����tn��/քϮw�������K�ϧ#�k߅~��홋��3��qR/��&L�ɫ��
����ts�?���/[��D���=O�\��>Q��4-�z+LL�@@�:�)s��d��K�֍�62���K;u�'�����is��?��<̔���[]�#1�X7A�w�	�*	]G��ѣk��U=@����p�z7��\j�{`�<�w�Ӽ�Μ7�:ʬ��n<���p��BSZ��%��z���A����JZ�Xi�t��OQ4����dԠ:����B��RBL����5u.��{凃i��\�gB��-F[8��2�QGJI�9�
�)T-`Uv�^z`R�+07���k����δbk�2�ԏb�U.0[*B�[���w��������!ĝ1�|�v�+�(�f��d�|t�2��Z��z:O#����+�WQ��G+��k��I�:{��]�����C)vL��U���|���=�+sFY>�Iw��̂{��/<�y����l�?E��Kx��5�4�iy8�D9A�F2MH�f,%f��-�Tg��e�1jV�td>+�7�ı�YH����YM�&�ŀ�����S��U��h1��z�!0�f��E��� ��A��ߌaY\۝����e��b�	�Q��{LSg3H�U��o�cY�S�s���nX^���oZX��m�e0�2S�_�0u�܏Kc�
�
��/�	KgH�^��>Mr�P>_� �w�T�K#�$NZm����#H��Q�x%�s�m����+����j�aTR�/-d���|[��|��J-��
��s�\���O�IsQ���"
��rH!�iOA.��zͦӰV�׌��N�Ŀ��SO��cc>�oÃ�X?w���9!!���&]#���k����O�9�+�XP'�N�����؜�I^�a��Ȧdu�_2M��Z�؅O �E��¥�j�ZwuPA��lE��߶��n��^+�%��?��������\�&�^�K�d�i�u0FKW]�bz�LP82b&���Fb$Z�?�F���/��d�0$j+��	�
ms����W�'���9j]h����g#��V����_�04���n�}bM�B���;o��$Et��Ui�6T�!P_Η<�8NVq2<��!u ����RT�h	�q:�-6��bU��UR�U����8h&�C5��Z/�8C*WW�ݩ�[I�ag=�9hBn��Q$�ad/� :�/3o�%p�Py^�-£��w����r���ᘥ؟���\�O�������j	�H0S��K���*05�T�ܱ;��E!:P�o�fn~�ll���N�x���pi`OoZ��L��\6���} �q�p_VP#�׸ǯ Z^�v�p��Vk�tFx,�p3?���m����
R[PA� �O�x�^D\3|)�59T��+$<m\Ӟ
)(�KLg��}��6v��4�J[�ƨ�ष�%�=���53��>����}[i�	��W�VyR?���x��d���LЬ�-YF�����nAI�p2�00���q�d�2�D~F�z	"+�jT�@���4��5ڣ0���Y#�R�K�%�5"&�p�9���'�b��/�K��ľ����xd��#��|�����G����hN�̒�+7.a"�4D������.Ԋԫ.O_��.��r�Ω���V����2��v�%Ρ�v�Ưw�g}��R�rEa�}(�u�b���=���	Խ�
fuI�7���EV��mnm��#���ᔛ��7Idy�9�]�"�+�H@X����!ۘ��FO��Q�vA����!��9V<N�~��:5�=���y#�Y�r�"k'/�tz�+���~c51�O�f�I�v���-h��KZ�0��4�c]L�[��<Z�܄8��&f����E��+�	�o{]��)n)Խ�I�H�����q��hhF��x&W��ao��Fp�g���HR,6��zx�L!��?ځ T�ğ!����,K����Z��ؿ$^�73���x��ݳ���M�yx۲��$	���`u�zU��d�o����e�3� ���QC��R�4:xb�����ڴ�YŸ'��vak����0'#�UB+/B�X�-:�ъ�!�\<���כ���Y�_ӑ�:v�cD�ȸD�ͦH�
c�ó�i���X�5�q��qX��z}��2f���:�"˧���Y*A�`�Z[�k�U��ԇӒ$"�[j��
��J��q�c�~�e��"|�Y�;Q�R�z��a~��� ���&��<űcF��+��z�ot�vx�c ~�5g�:���"�D���O�2���yb��ࡴp&&��=vn:=2��@�ꝉ0�*&j8�/����IQ���fDة�s��_ւ�����"�x�J��K&,�GTx4�ў]Faf�?��D�2�X�睆p+)ߣ)��ϟ��)�ޯYR�X.�H�)@"�mt��N�T� 3���{���I�n�q�E	-�z�ϖ��E���%F�×��y��B��@k-֔zm�$�we������"X��y�x���E��}̢V�zX��ߊ3�\��'�p-f�g��q��P"L�-�(쇲U�n__!f���>����1�ͥ�mvF��7����v��I{|PQz��[�gLvҦRq�ӛ�!�9��W@�4�gl�ZLl�R�3����P��RW�����@�,�?p����g:�!;�X������% $��޿._|�G�?p{!��Ww�Ԟ\o�x$���������rSӝ
ӓ����M%H,�طTb�'����OLS�w.�O�Q�a�1�ShF���]�T�	v{p»b����6U���jy�㡧�5q�G�1E�BXC=p3�����m���4��!��J6�h^��>��������}����z��C����������m�{�A���b)�4��';����M��،[���]�7װ��Tey�+B(i���M9�d�x�Aڣˣ�ͺ�����;�I;�F�"�����r3��֑�C���H����`�.<U+b���g�!�����B�}���(kz���d�U��i���U�����)�[-κs�Mz�������!��~+���OI?��7�Ћ�65�_w	<[�P�|�K��F�	b/���S>ıS�j��U��Md�_�G�jQ]5IʺL��Q�հrCB���Q�0��9�A! uy���g��M����P���TB����H�i,�����T�;��H���T�`��=@>]5�ڼ(ͧ+�*%�m:��6�!���46	s���ãcZ�͟�{�簔��~֪�&��������w\-f&�����rL��	_�`T������:�G=�ni��+��j��s�9U�ٙW��}N��X� SH<�^wz*���@̨L^���o=����e����d�3�w�d�˓���b�2Y��'�Wj>���+��z�`NBxJ1��NV�=VT�,�79���L������j��E�ޚuCFi�N!{Ћ�"%�q�!i��Ľ��)|H�V֤m:�]�}�b�����]������@2�Ta�����K���Ds`�j��0���)�e�)�V?sh��i��끤4CA�Z�����Bg�Uĳ�I�/����V��/4m�r��Ӿ� (F�bq_��b�Azث�^xHB�_,����2 �"`���UŬ���̣��ڐk!St5X{hTIX@�܍�ɘlغ��$���);c�}ar��j�Vb�tr)�n�Fǣِ%lU��Y#W������S�V��-~UӬ{:պ�g]�2�	�8y���o-&~�b�d�`�L��z<i�l!�'��ſx:W���z� w{l-���=�l!E��E��>��=�dj��k�.� y�h�����XO�dҞkt����o=e�����=�§�G�Ft
)'w�u������u�Zc�fb�)��Б0+j�Z;�}�<8VF����o�5�#?t�_q��Z��;�X,|8���A9��H�ò>��(�+���E��n~�Nғ˝]������*.qY:v�`�� w�(�ڧ֣���Q�C�[2˪ވH�f�K�t�d'��`^z�Q�K�Tp�%���;���7"Eb��t0�l!@�6J%QFA{v0�&ѝ���O����'H�,�M�/���[������f�r܋��k�?�j�{%�W����]���8<��3�b	���W�d��B��f�sP`�$��:�Y�:�@_Ӈ|6}�(����N��,�C3��	��<L�p㕨Lۏt{xg��~5�u���*����cV%�C^={�(�h�c�L��H52Qx:�J��M���Vt��7��\�,J�9��D??GG�����Tn��z�_���6j"��ː�Pn�V����=����{��q�L�S9S�h��vH���"��A,��Ɵe��W?���纗���i���J�֡��\9��c��h�Ȯ[sH�������	k�TkZ�z�Ttz�=�煤��I�1	��٤��7~I�$��\O� <b$Z:�YU+��D&���\����u
�lk>��r��I���f���F����T��V����'߱c��%��Vh^���%��)���������{����>�j/h�����*�reMO�J�������R[RqlȲ#�:U/������
�
��
�6��yl��U�>�(�Mt[H�Iٯ�F#�#�_�2���zl��
!���&j�7�ٞߴ/���}�\���|����@'v���.����ř��T��Eww 7��q�����_o�5�.��=���>���DQ�j��AU���ٵ�,~��0l�����䛐B5�)��L�U2�M��V�mi��$��&�I��B��lmcŏ�����H%i�*��ڷ]���[d��~7�6@���L:�q�XJ�4O�(V��p08W��BU) '�E�1/�Q����{Ls�67��'���~��J�{������y���m����*�!Y4	�����D��Oز59��BŻ�o=sVo��c�׏FN��"��{f;�`���OI���6�rg���+���Ŷ~�y����.\�ةl���/��$%�b/R�<F����zA\���֛�Y���Q.s8L:s��ں�g1�!�$EG���[��;^���ަ\�ɶ���N�Ռ[C��Z�:ď*���U:�!��r��gE�lv�6x�^��,�\�%���ǰ�2�6~�\UH���/�(��2b�m�����E�yJovsZ>�D.���7H�������Z�h{��7�qtŔrF ��H����g&�_mW�����mL^϶��l�$���z�7��������ɣ�]]��٥^�x�Џ;˱�b�5Q�g�饩S��AM��Io�4�U�&͖ ��q���=��e<�W\�����t�.�T�K"���W!�t�W�_-u�c����<8d�$Y!|`�P�����by�8�.�O�썴��
�iE��<�s����C{�:�d�)񩩩�������Rȿ��٨�)o��zZ*8_����ƄĹ���Lb{(ټT�|�lv�wtE�|!�н��Ġr���l����V,����$ۅ-EV���_��f\V��o�U�^ϓ�.��^ꪃ��&$�~V���.��P���|"�#M�DO2>��$����榍P��.f�����Gq'����\�}n5�S|\e$�g�f�ⱒk�1�Y��f;��^��mxB;Z�_������|"��%,	�35��:���o^p���3�>����"��Po򀋗<2�SDg#3b&�`���^L	�����J�x.�N��5�7����Zٻ#�N2�T�1-7'�o�}��ke06����6Pٿ>'Rq���&�C��)�u�jP	qK	�B�ú�&tO��E6z}��X٭��]������x�<n�Oؘ��>�E���&q��`�>�}�֢����k�$p��f$�=ϧ�� �)z�we��E�
�dV�ix�:��y�^7=,�W0�v஢f�L����Z�Vɛda~���V��|�W��/�O�I�|�Kx�#c��ñ�H�g�%V�	����v��LȄ��i��{N�R��?�S�L����+����÷G���p��|g��.�}���a��2�	F��#�bTa����o����X�;��I�|�?X8�W���<#�Dٛ:Q&f��;��H���u�M�^�/�b��
J��S��ϩ�[Α�K�wp���r�@�wZ���ƭ"��=?hV�毌t�o���I��;]���r����v���RV�]����>�tk�R�7�u*��Z�f��$|���#�|��l?{����r�E���x�~���t;: ���QxT��J��0�m0���Eݽ���U��"��X���DZ&����+�KAk�2�j=��板�J�a#���&H8����G
������/�,gv[$����Z��ൺP��z/�7Ӫ�[��R@3�����=w�vi6~����y��p0�~�
�[)�l�94��ڿ���S5"ĥ�I��n`����ܺFx�`��X.��O�7�Y(�Ԕ��X�jr�c�͵�HR6����n����Q��h{�d
� }��vN��mؽiTį��O���;�$;�xHܻ��U����$�� .4/�4bϟ�Pk!`���/Dv���_��ۣ넞\�q���@-�ƝC.R_�Xy �s�ǩ�89��[u$���E�X����G�cji�Y���.q�Fe��u2��_lA��1ZL'3����q�+9w}aN{��hJ�G���d�֟�D���Z�ܘ�,7�	�W�nI(Xc ��x�A�ѳ��:�5b��5�Ӧ~��C��\�����b+܆o���!�*��kQڴ%d�B#���o�+�{
���fnO�1kK�)ͯ��0�m�|Ӯ/IOۛ[�f��YsQu����[�\nZ�ߐ��⑿<=��ｊ;#�����s/� %��t�*�'�9��m<o	��/���6��΁͢=�)uy�����`תqx{j��>	�1�N�I$�i���#.�y::��S9���v�6>����ۯ�U�>����{���z�S�H�@�<����'��y����l>�]�"�M#1W������ҪYcw��V$��*��!��U���IW������z	�ƿ�C+�u���ĿW"��J��հ!�7'u�7`���^�]�9u�/w�-����a���t��HHp��^Dhn+�_�+L,$T@�|F�x��yJ�"�z�m��Ơ2 Ŏ����7h꥞l�����x�lӈ?�;-ֱ�"���D�D�TL��',xd�ސ$��)��{���������e�o7��cf�鹺KZ�I���8�0��.曻�8���&�)buOg�x�6���8��5��pJk����wlw�5�6iP�w#��U7�P�B�11�]JER��a��IB)W=�9��)���k㑮���#�^�SZ�ˡ��)&�G�237/bϭ�6ݢx�����)�E g�\T��:{q�:�I�>aM<0�{n���9��n��gg�ַ��j@i=�L��n���� ˮ/�X�n��n+F�Xq�g�y��5�^�eX��Z���?1l<�sKM�9b�(>���)T�#?���Y�eb�@�H�|�-`����r��x�e�Q�>9�D��-��*@��L��ƹp�<�d2��}�ַ�ϔ��l� ��*����Mbn�V.񁒠�E��6W�_n��h����_?�L�_�+���v��z�^_t�X��r|v��ٹ�����QA����l3�w�<����=ǔa�B0�8pv�=��f^�V����昣�������g��z30x�8�����2G8�6� �ɖ��a;� ���z�'�83
�ʙͮ���1��/;H2i�3�~�k��iNZn�B�~�
�l�T��G�%�����{��@I�,C��>���h6��8�`�q��K����Opww����=hpw,N���.��8gsꜪ������w�?Sā�M�}�c�"�F�c#O��w�9�߈X���]�Ы����K� ������r4�9G��v�X�����<?�T�+}�\��Fjo�\��=N�Ŧ2���=>�0؊p�h/۪�L�3X7�;9\�0���M�?�:y��t��\!�n*Zu}ǩ������u�ܾ���g�Vr>�%�bߝ�{H$	��!�qR������v�W�����9y�����>Wf[Y�aHI�;��;����V!v�γI����
:��:9�BK�d���2EF��.?%��~tW���U4Xc��lh�M��k�+����z�T�#Q��r���C?XDK9� R����F�d�y�	��l�	$d�[cZ*�6�0Ǟ��/�p�o8Q���'���:��p���1Z�Z�-L�-���.�tS�>5A?�kr6��^��1�d*��Gls�Y����u��~�����V�}���t$ �@��9=�߉����z$oF��f��}G�/Z�?=�={�
Y�l��S��0w��0�^���=�\xb�a'���2]��S�s�KQ�?\�/?�������-%F@�g��i���1�	���� ��0*CW�b��afV|5�][�2��&���KM�ޤ?>�'8�\���49�._qE�u��� �^�I`%k%w�v= ��q�)����H��z=`:g�:S�Q䡖8"S�=��X|~�j�H������(%���L2d4_^{v~Ǻ���6�Ft�H�a,Y�Ҷ�լ���Ҿ7��Am�ۼrY V��.���+R{�^�ٟ�P�Fүkc�p���+�5>���C
��-�[�k�Tz�n��EӘ�6��޼?]k��Z�O��7,1Z�q�.ߡ{�U�X4^��)՟&�+��j��"�Do�Ƣ8z�y�^��:�x�T����;M�|���|��N�HX�qK��i��p��w*�"ѣLm�;�� Z9(^�ow\̶�"{�
�7Riu���V4��-f�p�������8`*��[

�����BF5�1-���p���B������R�˗�bЕ��q`-�������mu��D�d�_7�0~���M��Z�f��h�H����l������g�L$Z�A@-^�2�W��89�@B�^�9����
���[�4W��@o=Y'�aa,�W����M��a��F��:�:-j���$=�@g:�5��g!�Efs_����0�e��m֒ꠃ���c//N%���4'"Ita/�y�ϗ�/7��>� �(�Pmu��oO ��|���x�R)t���qP*ǂ��5¢+������&D|d�.������e�C�}=ѣ�O�p��Ng-�$U�:?�4�����{5��O��0���C|na�إ��	�y	-��)�5��ե#�H��D� ��;���JJBԬ�ݪ~���Ҷ[֝��{V�ww����E��Zee6���3���ͮ����-����[u�ݳ��/t����uKv`������X�雧b9�6��3.���pGG��C�d}���h�Ԙ����`b��c:�j#*�N�(�`�;�M��a ��Tɟ��+�)���-�5���/E�����iB���:}�������^V3l_�ۮSD8V�Z��Lӻ�!u/ߦI���������k9;�����j9X���������L�$b�g�$�Q��jʶ��o�(L�T&�O����)�'v̮
2Vz�^���;��h{����wo������y��$b����Κ,�X;Խ�8�Fm_n,1�C��Z�J����3P�k�j��g�j,}��.R�}U��g����g dt��
��r����m�IE���.6���l��8�7�,�Tlr2≏�܍��w����uc���_$q�!���ȹ���� ��~�[s%d��L ������ C�0R�Y8�/���m�M�<w�����<���B�z_s�۶kpn�b�d�g�e65�P��Z�BmA�'Ɠ�F��.�H���"x"�~:�&�[���D⑖\�/B?=�I����uqc��|����`��oVӣ�	�B��5���o>&�7�>�,��D��w'���|�Q��l�ƻW��m�d`��K8K�|�����Y�:z\�V���L���3.[E���{P+{`?�$�А��#��F+vMLG7aqO/�Xg�y}@�鎱�tRԢn���%Q���^���С�C�Jܒ�=�o�wǦ�v7l�ö8c�<��t4Y��}�Ӆ��TulOX�᳋�)q���_4���ls�ˆE�V*�]�p��4���_�E{�4��S�B��n�+p����|J���!$_����`�����W�r߻l5������P���{�������T��1���@��_+N���է��k���Í|�[��]j&������v;2���R��ؼ'jG��겁���(���[�+���*�smQ�Z=�<O~��m��JZM���X�Em$q
c���9@)�<	����v�c�/�̺�rv� m�܅F\�^V�hŔ?4MV�0*�.;�xUHb�\����8�9���]��2j��Y	תI7���G4��ɬ[l��[C����˙���ܑ{�}{@��Gy����F�3N�eI�ց�*�Bj���lm	�;ӭ�|�5ֲ�o)�#�B�-
��	GOʼcF!;�&W�I5������{o���{��Z���QgP��00���۝�"�N�7�%���Pl'�^�Щ�[�t����(6�&妭8����$��1AP*�,z��?����%2D:(�)f��PRS��z���/\�~b��d=�K&�D�w�-Z����>���mM����e��X�V��8O[�5Z�)��[j�_v�GF�N;nxj3'g�ߺ�D�q��"�L'ь����C�ׁ�UZ����S�4w�S��{�vn~�:��e|�X!�O�D)�n?�uٿ4���Keb+�	6� �H^��9�~�x�5jd��.d4�aC��i��8&d颧��G��֟�E"�v���y�d�b�يuh��W&P���ɚHFQ������������n<bI����q�K�Ӄ�[�]$������u�ԄY˩� �E�,�_%���̳ A��'N,�0��?�`�e�MI�I�������ֵe�0�����<\���T�=}����	Rݹ���v�+��^�q���r�k|����FN�ќ@5AX&+�*���G5�k4,c�n���;�ۨ�+��
��4әw������������{y"���߷��\��ڄw�I噯��B���P/P�D�ݕ�_k�,�{��Ȯ ��i�\�T��_����΂5�Vw�e�6O�<��J���љ坵)<9�����ӈ�<MH��ko�IVOI��tc�j�;;�
[�=�篷n{�{�g���_oK�y1�C�L��[b�xY��U2v{�a�V7���BEN!���R� �M���'�@#x�`� �[�au5B��c���8�y��L�
��H�ԭW?�|] fL�sVTP�&�ݑSo~xe�9�����c�#B��/A<ܓ�����5tJܴ��v�'��u��[��)՞�{��C�>����԰fP裔;�ƥ�]m&@�j������ꊻ��%u�X�܅�O&	zTc��>%Ѭ6~�A�ܗڒ��M�=`�q+�~����ѧ��ao�@x�K��+�ڜq��ӥ�m1�����H*�v1���Y{�|���TǏ:�'j�ui!wua�Ȉ{>-팬.�s���$pwa}�xc_�yL�!���k��/�6���l��^e%wF�3��Hװ�߄�Wviݯ�X�O�r6��\j�o�����w��F
՝? ���Wui2�Bc�_��K0 ^Z�G�=��~g�{������]�7C�s��l�չ�0��IT���A�t��_�G���p�Y�B��E?�)%�}ؔ�8 
\��ےNo{U�Qs�|9?�杍�}H�_�V<�:�kf,B.�z)И�	�*XB��B>��:Dd��h��ϖ��R��V�q%3�{,�6K�t�x�=4e�U�q� N��丹�n#��d��(�S���C�it飼�����N�դD���EJg�O �#>��%�j����ϐ��L����&�1q�D����_�Lݮ��5x<�Nu�,Ô��G�y��C��1} ��C��{�xp�����������&�E5|d{4�:�Ӗ߱���\ �����I��R��⻁a+�[�I-J��(�]���>l���zh��*�*�+$�i�u���3��u"�Y�mi^�īuɷ����4u	���u�]��7Lwbz����ڛӣ~�)B��ׅ�ݎE~���S7\l$*l���-8~�2\�xMT7I�P���v�GKT��D�!�W���S�)��?��sÑ9�]�[H0ԫC&'a2������oV	�jŎ�Bٿ���$�uz����o��2��A��&v/�C��[2햯�	hz������ߕF\�?�̷hu�ٗ��{���^F;�F]��2�`�����r!��u�D�4�z����܅���-���!�43��1b��:��qh�N�Z]�h�����T�c��r�Y�0:g53�jF6��-�����jTW�����5���G�Q���n���	�G��ɿ�)8|�>Qu6�:g�%��¬z-U|j�
��-��λ�y]|D��W7~�ǖj��-8��� ��Oc�n�4����V�;S#�f���S՜I1@6�i5�|~��ɑ-p@��=�#�8%��E�K��Mb�2���A��V�Y�I9W Br��ؓ�o-�l����z�]��Z�~ʧ_o9�7�h�������C&�4�*'W��P�H������&
��7�u�H��M��]�|y<������kj�>��թ��`����]���=)����Xm;�z���UFj���o�%*l~�I]��9���1��1����NZ�����٠�}D|a���z&+���ֶ�Y}iB'��1���_�i�Q��&@�E�i�[o.��j��0���<`�D`�23�U�Iϗ����d��!�:~*���Wy�[FI$օDg
��qik�e`�uu~w�c���o������=SyK�~�y[YXK��H
�D���w&(b�w�V��cͦ���OE�t����i�����ق���K(B�K�*�A��Ǭښ���Ϝ�R��ׅ��5�6�m�i0��P$W�I�����!���T\�Q,N:� �u�ߤӖ�Q)�T�u�>~C hF�oKB��͎f{�����3?�LS�Zk"�l��;�e�0F�u�u����N�����)�q�֑��R��տ�7��V����ƣ��l(��zn�L�^*�^�y�
�Z���9zIu�e�����V7p�)���U� K��y��䴘���>��C����t�Y�ɀV�X��/��.p�ۻi�e`B__-�u%����҆ ���_Ok��0�^C�i=�V�S�#����P���˔S~KS$�l.e�v���܌��oG��]�'~C(ѭ��*�I�o�YzI'Q�/�m��[0���,�͈�)�arAp&4ä́�ik��8�V���g	���2r}��2�8(��5�.d7�6�V�f5-���O1����_K|�x��E���m_���N�-Z��Li��X��J#�#n籖�_hU��F�U���O�o~�a��o�{<�^4i4>�������������k>�����E���hO|D��i��x"�x�"���qp>����m;�@�t�e�ֈ�zI��t�֘�.���Ϋ5{`�m<�
�XG�C[�?K�}���Zﲌ'�4��z����=�*�\� Oۙ���� ���o]}��~T��,F��$���̈́O�f�튮�X�!�����YS/��o�]�M�e$ҁ�R	4�{�m5s"~����K:�>��%M��{�	j��&���뵥@���V.!c���]3!r�~�c��Qi**+�o�<G�O|�k�#x������|8L�,$O��0��|%��z>Cw�$
���I6F5��
ɝ���OPי��b�/C?���< F��%��єם�O7�o�-n�r�'IZ�X[��٣αB ��G	jI��X�De��*�	����f�G�u�v�^����-��n<��L�"����c�� _�+�?��s�M�� ��v7A�����º�7�5τ��5[3vr6���h��1۔�&~�z�N��X��6�O��oԶF��U/���mzN�ȏ**3ȹ�)�"[���HН��r���d��$7����51�V{?�}��$�RZ��I�ҽt`�<�חۛC�=�>fɲ�ʫ��T�γV8\��e�M��ND��\v����-�pQ���an���罴����+VF�ĸ#p�P��i��(�"1I�Rڠ�����ؿB�I�O����%`޹��c9����D�+w�����h k������v`�:fv�����3؝��Z~bp۵��E`#�s"�<�e�W�A��(�{K�PY�o��܈����͖>�G�N*��O�Ѩ�Z_փD0A�9k�"/NE�r� ��"J���R�őqV�҉C�&yD��<u�6�"�eL��>:h�t(��x4N���UL3g�����%s)n�7�M4�y)	x>�˛l�J�Q9���s���.U�K���L��������L�^(}�:���g/���J ax�j��ܧ�7��̈Lw����ኑ��z���$�Yo�/�l�(�i�xq"s�Oj�t�M�Hn��8r/]�Q ������P���/��7�ҎAb�m���m��/f0~{1w���D�%�*qε��!t��� d��p���3�t�i��?|n��c҂���Uma���4��n�`8}����,�FHy���u���X��O7��7R����-ODV��\č�v~�{a���n�=z����q ����1\���~U�tהa,��xX��8PW����d�3}�Y�u�����8)&���>�(�?pc:�\$����)�H�m+-�L��Œۗ�v	�SV����h�����6^3)�لTg�j9̿���$Z�Yk��Y��)��)���׮W9D�N�P�V�Ƞ�O���3����n�Yc�&)��zK��G�3I���/�������z�0��6L�CT�qпVs�j�e�A#p�y"���=�_���M�����I���ѕb�Ns6>�;�V���-<�3�}Xt%UO�*m��ޗ,o�h��)��	�ڙBڎ�m��u�h����Φd�n%�v�VJMY�.Q�M֍�7��`����\W�3n-9�7�����idm���� �ε��P���z�o�m�0������T���ѵ6�>?��g��a;� �l'�էӎ
������1��?d�P|����.��-LT�G����$��;�%�?�P�����9ڬL��<��{KBKoJҎQ�#&H�����[�$����.�۴�L�S�FZ�{�1K[��ӌ�N��5�V�}s����\��_�ʍ=������_�I9���#�t����x�u���@�u���rs�x���^�;w[
��;��:r/�V�v/溇؊���P��⑎~�?��.���|�!�.~Gc�mKw�sM�P�p�\�i�������_(�V�h�[l`�	���64}� ��6��_e�����#�`Wf�)R!\����D���!9}>�N�i:�Uߗ�ˀ��9�����<]��
����a!�j��0�7��M�?��\�7�g~�%�)FX4��^߶_S�;��4�9�K0��fX��(Cl�lۗ����ɓn��5�e�T_�̿�����YK����O	H$��G"^�t��J]�x+�缠�$2���r�זL7_8GWz���`w��o�˽;����h
J�뺳�wF�|!�>&�q�>��Fz��B�x�Ќ}{Vl�4���^��Yjnxx/�x?o"��P��iFt��~w�˃{���h�i�����*s�Ϫf��9|��g�c��r��_	Fb��Lʵ�B�e��l�E�$��o*�(�J;�i�F�+u�7L����z�P2��֯�>�v�\T��%
�O���7MؖŹoi~�*����x�+�֢�joM�~�+�6���p\�|��9 @xҺP�	zI4j��;��c�i����Ȁ ]������IKX88:N�Ek�_�*$D&f&x�`�mN�̨Ộ�)B���I��{��:ܸ��<�u¬P�s���t��n���1�_v�e�%�[�"�ƙo����ȷ3rߘ���\7� Q����/�m~��x<FQ����'�i�1���b\)��)ۘ��0Ԏ�3aU����"Ǧ[@�o�^ۡ�紘0���<�_���pɲ�m�˴W��J�q���e��Ȅ�P�~^5e��#��AЊ�U�#��B�cW���8U(��ǝ�����Q�K�x��#p@y����;,@Ֆ@�'L/�a��p�I]���>7I�=Su�=DA�DǴ�[Z��f0ɿp�O��N����E�G�VّNZ�VY�؊���F�p�r��uw8|퓼�^�dt���3Z��S�r�5��Z;�A�	�`��,�M	o����y�c�WPK����f�����Y�6����"��U�kg곾��Xh-�mrÙ��*�C���RA�K����K�|`�X��t�Q�y��Qjy:����&�jX�G"��~�2���'��Fԃ�b�.m�C
v͐ԛ>Y���-�Rv�����vh����|�9һ�3�����6������Ԅeoe�p����+��fЭ�lXSWa��`�\�=���e\X����>׬W�M����%`]ҩ��.��N-���q:�ky��/��9:��	��
�$�1fV4j�;�t �>/u�ט����c}<�|i�����>fM�5�%H�r0b��)8��Sf���=mS����`�P��|$0�g!�'���2;�n%�T���7_Z�ȁ??��;��xN��8�G؟���w�z�p�J� �U�,_����q��cF@�Z��(O�������Qc���B�MGL)��8�|'��%�X�J�N��*E���>y�Y���w�)Ŭ����m��ly5�q5�s��r�%��b̭;���	n�d���w`톍���-�	�cҗ>��d� Ӟ�W�÷��R�ƾP6Җ�9���)�8�"x۴^T3Y)&ޤ'���l�K���Չcqwb&^�9��3�,�C�:�Ag�d���l�r��~��Aټ�H[L׀���/�&'q��6�t��}V�
�������ZVO���D�L���dc<o�C�vk���ǜ��xH/}d�ҩܿZ^��y�iԶ�I���6��'Ơ��R�j�4�Y?���y�IA�YL+��0󽲄�K����aH���d6i��{�l��W��|�n�~1ǃc�����|	:y��	�zB���e��y]چP�%�7��D��.������Q����;�^��w�Q���9�
@���[�E�L��M|� ����kr)��0P����m=������������U	6��m��X]���!Xߨ׫}���F�z��*Bo�|L���Gڈ,z�e�L��T|��<�[cs^�.��/2��4�=7�'R)���?�o'h��[p�����r�D-�N��s��8�4[�-����w������dоl�>ON��
�@z����9Q��,6b�?�E�Nm%����U�c>�^9tb�j��+>)�s��gaa�B�X	S����g����h���Ox���)��2����~��J��p卯#yl�z=���c֌��e3�����]�|-�hqu�����y�������I�V�? ��X�K+K����Jz�q}7�4ǭ�������2d���z��Ze"�p�x���p����?�����!�.�y?,^�7���rˀͅ��1f���(���iH�B����[��~�k�o�Oz[]��������x���Nr:
�h�˔��gxթ�t%�H� �W{6$��~=��Fnw�t��/�x⠐�J���컡4��tO�ޤ��N������������Jlℙ��c��h�~�����2��BřĦ=�+
Qh#��������4��)m��0���%n	������uת"
�߳�2��r��������w.1�SFv�C%��w�� &�c/A.�9Ρ�i�gg���1�*+n��I�W�Ӈ>�+ێ	*S&-%Ŀ|(3��X��Tn�ݻ"~�Яj��w��`�uZ�I"$13rG~Y�l���Y5ط��~�[��tf�^C�B�qU��O�m5z�Ό�=�Lx�d�3�ƂJKԁfً.���>�a���@i�8��[1��/���۸6�$�Y���(U��o�ީ��$�by��,�b�y��;φc�� �/����Ϛ��k_8�"�ܼ#���O��9�u�]��ɣ����^��/�eV��Wm�]�8�ށ����5��R%�t��`aֵv�~�\�D�w,�h�������*"2C.���5�^
�i.Y^��P�s�(���cM���@w�'Kݬ�g�B�����F����Kr�H�޸}M�.Xx�y���?L��-���X���^��*�G���i�ؓވ.�
oz�bVGk��2v��7��}'C�)l���h�9�u�J�X��D�Q�'�K���d`�v+¥M��k�"�,�/<m�c`��AU`���Ky����q!٪�e� &;#Q���!�}Hi��L_����d�0h*z��l�;XNe�������6�I�n2Ȧw�۸�����͖{��"�?6��A2�y��GI�e�ٴP�ˡ�V������'+hr�kI7�v�=�\{N�m'�*
���5s�����ӎКI����ٛ;�uv�N��5���������r�[�p����&6,_�_s+roŘ�N�_��"��j��-\<�t(�\?�UYC��H��,Fp<�4]|R�]-�掍�:tCB!s7
�ŋ3�4�on�;st~�:��g,���m<|�I��?����\��k�F��i��-����d�E��((���Y��`"�ΐh�K��{��Z�0t� �.�C,r(���j7�i�x��;��o���ۍ�����v	�2!�'�,Ⱦ?7h�������Bu��n�����j�p�]���%r����$�iQ2s�:��V���2d�$ǯ�O��!N7�#4	��ڰo3�ğʣǛQ�8�t0#5a���J�?��ߴ��{+�P�r��K<�̇���1_HՏ���`y��o�$&�� ��	�ki�u���y�9�6��~~{;{[��Y�E���zi�-��Š�*��_�Ҥ;x<Kj�4�VL)nyt�BЀ�'j�H<�d*�.���E��'�ʁ����y���=�ɲ��>�}��d����N��YY0�϶�Z@1� �i���xRi�\�cxXd~C�K2����8Td���՞CӕL�1hPѺ���?�`�����)ԴT�o���B���<|tu��+oM���{U4�$s%#��]/+R�J
�5c�U��խ�}hC�V����)�}�������������:2t��v�~�-��S�>F��R����9�I�^����#
���X�M����$��3����[ɲ����Cǘ�:�r� ��z�U�DS�Ο⨏G���3�� ��C���'GgX���mw��lϣ�3zƵ�п3|���#��x����hi�+���T��k4:F���7�4���>(	XTl���+�x����������I�j�����6U&jv����59���yK"?�����|��%��E���xz���d���}����d(�OS�fDM�8c��vxzsv �j����+_\�H���~����q,���S�C���A�W�@��|�T����kp �5D-���?q$~}c3/9;}@�	\�Ż�L>��E�/��Vp"H�tHW��e��T-u���4X��ޠ���p�\߾�Ň�)ױ������x�S������1����Y����삇P��\�B��rh��-�a�[�X`D�R�u+�Np_�1�����y\Ͽ��;��(x9Q+�;�o>�6(n�x"��N���S��s��p�:��^�=��v������@�����1�5��Pv˘�~����ﱀ��#��8��<����?Uj�^z��<�������U{M_�p�LKj���R��t<��DpSQ����%O����������6hn�Y����.pM#���g�;���Ks��VvK%�wh�u%�"NīQa7��`�d�����;��R���Aä�W�WK��fd�縔��aXc��)�ؗ�QH,��N���E���|֔��f��U�,�V0}L^~Q8�?����O�x��Gvk��b�+�]�ꈕ�l��'8�D�� ��p[��<B;h9~*�zۂ��h�.:�>� :56�  ���Ҿ�y^�6��B����'��َ1�l�n��wq�!FE[��0}�{;U�F��.�ם��\�j7��G:|қࡶW �՟��T�rK?�G��A7�K�tu~%�B7��_�$`�F�3�\d����*��6�)�R�䙧p`� ����O��	G(a2�Ci�%�>��[��ԿL�U�>�v-�֥�3z���|�8c!,�Pec~��j:?[n�`���o�Z����Š��&��e�
��L��Rc�8����	�	(Y�MBתȐo�:�`�Zkץ�嫞G� ԟ��� :��<a5�A����H���2���h�Xu�b�}����.W���N���b_I/_o|�Y��
i�~�x+>"� U����l��ȖF&�i�U����Ernk��ԁ���M�?4��WoJ�u����tS5|Pe�@{���B����P~��pk�;m�q�U�{0�4�K#&�W���깠����#���޴c���r�#��^
�O`���f�ɣ�%,7���bA�(b@M�������6�ĩ@����|�&�j���	�]��3qh�h!��b����������3eol�TNr�Y�G�hH?Mh��xd_�"F`=�C o��fdƨ�ư�W�K�7~��E֍[+�ʎ�w-2m�b?kj�@:�;VĬ�P��x�:�ن������=G��mվp�у�hl�6P9KoJ��OP(xFV���9b�\z���0�I_�Âlt����F�tza�w
Ǜڎ��i�Q�@�};�@|�eύ�B�z44�7F�
�������k�$x����l7�6��z�ڳG�����ܨ5����'��9�kg���X	ڎy�Ug��$B��سX������J?3�Qo��D�Zl�RQ�X����fbͮf�%�_!=N�����D�ьJ ��?�pu�4ߢ�o�~��̤�^��o��c�w�G��|:|s/FSw£L�� h�xl�$���g\�X"��,'�_%F��B\�	V~bӗp��7�B�c�
�m[�2+��t��q��翎���'�I'j�~⏚������`C�j� �{���t�N�7B�ܝw�;+������\�\]s%����z懝�_����OT���OF���><�(#��MJ�b��}��z5����8�g�Q=f�,_���gsua?�U�C���P!�ՅM���
V����S�mx[+'��O���Ƒ��m�Lp�.���]���U���5�bo�}@�.�Y2�j�z���5H\�?M��74×�ջo��]�͢>�8�~&�-^�?t���K�z�7�9��@�z9�B����x�g$�_#����j.��[���Bx���υ�[��ٵQ����䋍��
�6:�T�1e�-'soى�����R��ٸ�9�Ã8]�*p��g�,3�ʪ�h�����U��0�~�7�Q>^4�D��*�e�I�E���`fN�e����Ѫ�E���48Dz�>�Tc7ʉ�PC�8�P�^�S ƈ�&�C�������J�k��Gu���ޮ�^��aR��:���$]6���9�id᧚���'�)Y�cw��ݐ�׮Gdx������V�*�q����K�o��l#�>Z���{��B#���(4�������(���V�x��V��Z�M\�Ȋ��i�oث�H��&P�՛�/_z���.�S_����61���=x���WcseG�ƺV!�G���K����-��҄
�b���KVY=�#s�KЌ3��xN�aO�q��1o���,�(O��X�I��w!9�~����z�+�E��E�C+q%�~�_¿��7��m�����Jq�s�?	2b0�7WcO�˔l:�Y�h�cX���
�2�6���?�`�w�~�o�$	�O�&��F���Ƿ�n��=��bgs��}o)��.�,C\�"�x�i=�G'\Qq�[-�8ɕvG�l'���*�B�Cй�)
�Lg���D�A�D��I�T��(.�~ ��<6��a�R��e���|OQ�r��> ���V��O���sT8W��!�鋡�-��.�S="�?�!O�@��,~��^��6q���-8�@ �3.���4Q��!�}L]���K��ׯ4"+y��f�r&l8#�����d��鈼Q���K�n�~yE
ŻhMj����n��/��΍�T���2m�,0A�qX��$�t��z�[�̷F � i��k���^�Ƭ/�߿_��#ȨW�t���\
`��$�3��*�b�p��B��Żr ��RR;��DO��@"*
0"�0�[v��RJ�U-��V�
��������U�����'l�Kۉ��H�⨡���V�"?J�������ƒ΅�_sSw��3$K���W*��)~x�Xi�K��=W�W$�Bt�H��W�������
֨܈C���:|]��6q�Qͤ9�,��Ƨ����K��
�2Pb��B?�wT�§�?�����sfX����T����sxn�/)?6��A܍f�W�:߶�Z����,�;�}�ֽ$e����M�P�Zˇ~�@�H�K���ܕ�z��q�T�/;�e6e(j�ģ�V����GN�6�.x��ʄAڎ,��HF)�����]�<E�C<XSv翓(��k!"�cp���r��I����� �5�����L�U/s��R�VYDB#��������#����ǹ��Yt��xQ��S�}R>|����ʨoGW����u�l+���8��平�򸸑t*w��C�W�v\�Z)��c��¯����Jcꪴ�G��9o��FL���� z�N�[]��6�DXl��s���C�P*��{�	�$({��#Q*�F����,F��v�8�f���1%>���_݈+�0�c��S�����\,�2ooP�td,0r���a��i��?q�Y�����@�?�6�y�f��>�dp􌇛�yH���sz�+��/J�>��y � S�wZ>;Ky��*s�%@�GK���;��������YKѮ�R�bv�g���Z$!�Kh��y�I�l�_
:��$1j�y����ۊQ+�̲���� R���j���n�����,�d�Hϴ��V:>��{v�"b|�D�,*Y�����i��������)-}������y���@sū�X^��oD��_x��	�f�݅h�'p�]R$P���[ e1������:zR��y{������Ώ�;"G��pB�)sB4��:>�K�����9�xS?�*%oH}������c�#;��7s�#�)u��Qbu��`��w���i��+ZQ&��4��o����0�;b����+d�f��t���\^L��Eh���}�?�N������Դ�"���
�/B��%ϥ�WǺ���EVS�׃��j�������⏅H�T���q�{��P�h��<V���)��*�o�_W6�x	��&~{U�G�2iC:���J۷V���;�PފZ ����6E'����7��YXS�hC�)��Ak&\�&��?���wH\�J�7>�E�-��$w���ǰ��:�-�?�P
���ǧ�; |E6��&f��M?��`) �A��!Z`m W�̴���c����s)��!�	>pv�ZP��߲D_�hǼ?����# ���64s���4���Ç�@��R�1ZW\n��q��*�4��X�'�%��^�_p�v�����mO$�����:tqY���X���'W.~�����8��g�"�\4B�dQ����\$�$� �j⿯Lc��'�͜�Cs�x|�칷��Y�DR��lR�i�$#F��E��ܦ7֕�FӀ��ި�H̦�.�\��Ah�$z�߀,�^�xq^9��)>σzS���\�aِ�p�ϧ�����H(kiR>��{|qaG�]ם<��a�Ra(Y�ᬣ3Y
7�A�^�s �w9i��E�F�?����z먪�.ZEA����$��C���K:����f#�ҽ龿�9���c���<{�9ךk�C��Ü	��_;y5������<�;����4H���}�������]�<�w��u�����Y寸5KYN6����%��"�� $R_v(��x<e��)�TeG�V�|<�1/�pm �L2CL>��J��=�±��*�))����||�^8��6Ѩ�ya;=2r�dd�HY�].P��<B�f��KX�u]�J (
�8���o��?ͪ_�]�R�>[�J���E���1Qwv>��7"�7՛��,�fE�~n Ax�IEL}y�`6���Qo�2�%*/����\^��4-_+9���x�
р�H��!��óh���93M9��3�ی�b�e���w�n�m�X� [;��d��ݞ�?���5��)ͦ�;R����-�99wK
�״*���G�z=�M�xOe��QeZ_D�T����!5�^�=L��}�]�OKqӧ7Q ��Z&�$₯ g��l���.Y~j�'��[��h&o�d {]�����vK2o���R��iy�ce��+�q�w(�M*�K�u:5�Hk1G 6^xR�o��Ȼ�M����p$�թ���E!~L��+�v~T'lqtٽ���$YXq����iE�VD�&H6��D�3�`��]���9e��c�Hq��d��Z�7�6�?Qϸ^���P��{< i��H|��W�*`���[�h��M��%���{�.|!��-� �*��H���!��p�`�-�[jh(�X'�V����PL�0�'�C��S��d=���J���_2 ?:�}��rM��Y2�Ł ���K��M�2b5Mo��.�ĩ! ������w��ɺ�ٙ��Ӱ`/.�"gϗ>��)��
��[�ԧ ��s�T�K?趼���	����7�Й*���Ȼ�J�S�3t.��a٘�Z�=�=���������it�����O�-`@�7�f��i7LީƳb�Ȫ8��D�/��b������d��%�'�#I�U��|�����w9�/�:�X ���D�AO���:^�74R�)߰��j��8��Q	�]ݫD���Po/&�2]� �؉���2�E� ��m���5��R:��{,;F[H��ճ�AڬwY3*����2|.3�BW�|mIu�$����p#ϊ >���
�K�!RA�er��eg˲
�{.�&���bGD}���Ӥ���\��g�G���]d�:��(	�ҹ��X3`U*C�5�#Z/#���A���eŜ!9��@�@v���֓�<����n�'�cʛ�g9NL��!#Eq���Ү��Mp�s�0�BF�����R�I+BTu��V�t�Ӝ�J�N��"2�_$̽r�����s�Q��j���I�r+�ۈ�&RN�Hi��PQR�h����n>���f'�v���,� ��kb­�m�
�.���R��8'o��X-҇�Nj"Et?�D%��D��� ���D�K�qF�W�~;�-��K��0E�-����c-/�Y�4)*�q��}Ob��G�Y�C�_W����3=T.���������ӎ��ms���%c�ӂ�?*\�x����T�WI)�:/t�!5c!h��e��٦	ZIeg��9�my9Nԋ�gNO���ڂNj�����C�̕>���š��Jм����~���Y,�l^_��k�;j��p\#JM���]�,��T��C �Y35�����5��nb�k*�SQu���U�������u&[��j�R�e� ��k
 �B�ٴ���R�nڣ�h�<��E�Ġт��V����%��%kaE�ؤa�>�4����1����#z0`݀){�95��s�`�p�vђ����5Z�h�X�D�&3��eh�i�,��H�X(�\U����T��.������������[�s�LD�ˋ��rbr�ϗ��m�g�?������eb�Dx�Ѐ\���	�s;����.آR
�Z��G#����pP�'�$Ǌ*���3�Z�,�Qy�a��g�}kaHo�Ķ\�_��>�Vp�K������&� :�6����*$�\^�F-5�%U��r�}�O�a)�ِP��&�wy���[K�d�7'�J�|����������L����&��f��F�J���7%D���4g�5/z
L��	����
�I��$�*Ei�E���	�8���T���CG�A��UZ�x�1f�P����&�%2բ����=��=���^�˷μ��+6��^F�1ewm{�s{.�)&�Y�q�2.���Lq������틫��c4�|v8<�o��?N. R�A(����<ѯ?�QE�D=���� �%7�L������[��U�U�5l�1�XT��}����S����C"��U�"�-Y�)2�$j�=kA�� e�9�rnm�>�4����wbc�$8,o8N�&47�f�V�Q��
\�̓��>���$$c��E�����ȪV�M;A���Qږ��t}�⢜zJ���Eox����nR�
Xͼ�N�`ڼ�J$Ҟ�טX��ŭ�<z�Өdye_�zX��@ʤ��V��JN�%�[A��ҭd��L�/bS��Ҋ2Su�����m׶�QJ,Ċ!|�����Ch|��F
$�ʟe�CR�Ur��Q�!WW��6y��;�8�-r�'8��9�C't�8�k����]�6L>n��(�A$�z$�$v�FʜQȊ�e*?q��w>{�I�?���w>�43��jL� `�Ws(�a��
!�}�
��;Bhl�xt���>�	A������d`ŗ�U8�rV��N���A�.oP>�yX�0G�g��,g{�x�'�>�Ry�����\��������φ�P�P�mA%:�pcD�9>�쭛��
�^@�t��^�< ָ�/��I�{�Vt���HE�y>E���.OK�F���û���9�}[�I����N�-�԰��UY��ξ�=>��^���Z۱8�D$R���~ș�!u�Pe���&,i�c�dHL 
���T^�f@ν����/&�yB�=%������ҍ�ٍ�	��-�)�� cEJ�B�`��!�d��W���x*�ߣ
�%	Ka۷�ȭK\r#��K�T�����iT�=rj�lg������]g,��QJ�/��!�p�;*I
����^?��e��9H�j�����f��c��'��9���9��)����9�T��r�S��`�]9i��Tiލ���P6G�!e��"��;�wop�W�m����Έ�;)X�c���n<�)������t�)J���80Ko�Y�7A�H	AG}�G|�c�o�1�LV�o��Q�����>�?W���5�n1���{�GTTԢ7M�x4��	Q6��ɞ��l�f�d���1��2���t�.��w��p���å���ɀ��&��E�#,�M����B�0$�zA�l�G�C��G\Nr^�������B��&��vNˇ���!x�䶂�f�d��8����M+eڲџ���?Rb�?ѵѱ<��]�À��:�0��s�M*%���Y}Z��:���l��ט �X=o����8q�1���Q�rаn�7p*��eS�������DQ^����DV\�g�p�~Y�46O��I����R~��έ%׊���iЗ �I���q$g�y�Z�2�Q����d����H�Ts����p;��E�	���p�H���3�.� �(].v�>)<&@j��oO4�8\-�����l�sIAFF6M�NCY
l�6�[3E�7Ͽ͆�����U��N��^�����������Q8�D1��N�DK�ԩ� 慕 �����9kA�/���<>v�0Q�p&���2�k5&�h�Fu�a$�J�м�W#�6���,��j��y�)!l|�i�Y����r{O�b2��a����"�����)�x�W[LBp�N����z�<&�8?Q��$��t&�"
�h�vx�8wt����r��!A�La������~��
���r^�J����~�D�jʒ@��Շ�����4H���B�(VQ(�`x���_�Z�Ќ|�7��h2��~M��ɼ)&��8E��w�r�|��Qq�y��;�g$?�B�� ��PB���RB��MR<��t۱[�O�����\qX�$aR�,	wS�p'>,��@�*ͅ	�
�{���s��L����_|J$B:fLgLR���f�7,�)i) ��%YR�'8��������?��E�HK�Ɨ�US�� �-}
�߀���eq�[���Ɏi7���eùCz���@��3*fBK��oB26�ا�)���=�;��@�%ῷ�"��$E�%7��m�������&`��T"$ԏ	T�&��*����t���ߎ����
�T75}�HA�"� -*���d���YM�B	< *�*㿀$H�݄����`B+��h�r��ņ�����q�cK3g���T�$]U7�$])(f����R���6J��kt0L�e��72�mA�{��x �Y���m)I�V6��/�S'$k�D<L�w��>��a	"L|
ϲ27�JE�4!���a[��%:K
�ҀU�ř���!���8$1V�T&	����@CB�}Ҋ���Cq����n�(6�R�@q������J�� Y�#H	zBE�2�ג�����Y\����<�k�I������8���i��]�U9t}KV���?u>Em�\���P�3�fpi��5%�>�Z�$���0B�ț���f[��l�_A��c����V Rwb���uw��r�D霺�Yx{�1��&��[�����{#.��[�6����B�1!gI�c��(���/���Qh���9!��@�
!��I�H%u�ﴈ7��!�E{߿à��,C�pV.u�g�>r4]^y�(���
�N�pτh"��3E$ �]:|O�*z��u��"&����&)���3�Kt��+Ў���g�(���1��~$YS��a�Zi���e��aי��_���i+8+U3z9^O��,!^�?�S������'���#��{f4���K�9�ʟ���������V-�^4x��/���&ef�ȿ*�D9��I�$6Z�0������;�� �܎e��� �V�ť�Jw�Gb���#��z�<��A3>�w�T�j�:Q�REa
��5�
.لG"��E�?��ń����q�;L6������W9�8�l�Li���To'Q ���
��	q��I��2Q=q�[��J����/ΥJ��L�B���������A{���a�|z�a��"9	��W�}�E}�=���k���5��,H����Ua&5ۡЮ�0@����H���r�(��gx��h"3̚� 8�_�H��I��nӀ���}��c�@
�?�
_K��p��h�!��?x����n�cy�rD%ŧ�T�����V`����G���Tw���̛���U���-� �.R�=�^�R1idԼ�`�2I}�!E0`���(��O;a��,�]��v���\XU�{��*-�2�6J�vF����l���ya(�>&�%��u�"��̿`�IȦ��� �M���w���T&M���?���c
*� ��'d��\�X`ݎ5_?��9��I���Fu� �GU��eTs�d
�LxoI�h~֨�w`,6,\�-�k�S�5F�5l���@� �YN��Y�_�-�(F�e����a\���"�D��>.H!�do��+�X~����1��6��/�]�����j�ޖ�2�/�����v����d,(� �J_�@<��� >RpyK�+�?�,5���Y��[�m��餏8���긼�d��[1K��c���v��u�U�Z���_rd!�P�w����T�'S�� =�@Tc�}��Hɨ��F�+e�Kt��E-Eb4@Z���=���������^+dG�.��[�"�wre8��s�j4ڱ�Hgh���ch�n1%�~��F3�u{���'� ����8�H<8w��4��somv�t.e��+a�|D�@}6�U��&dT /o��q��z��إR|���gt���q�uX9#j��!�;��bue�Uم@L{gc��
��
����g�V�]�����=����spDQ=e��y��.Yɀ�k�ӏ-{<5�|���>�I�{u���yQ��8ձ��~��B���!b=ymF_-^�C�6���,Rh����(��/B�BP�$�.T�}��	���VG	&��,U�i��j��m_Ct+ޟJ;'���bG��'Y�|17�W�b��L=���s G�]�<z����~��6S��~��`A�@�O8���Dl�w��h(f Db#Fb�ls���F��}�C���&��0���6��D��?̧9}^�e�2D�����d�u�?o��y*4�����f��D�.u�c�!+.K�?L��<�O��j�LkI�(L�J=�wP�e���K�k�'����Q�k,�[/��O�- -:��ϗ�G��9�H*7���06�O��?#��w�f>��g'�9(BU�>�W��	{����t�HUW����LXHZ���P@[��m�֝�ZmIx/?Z�te�O����PZ�V{��.�26��K��N<�Q�t�ǼC �����n�U�Y�2	�θ�Ze����:;L�N��o�S��X�
���5
�_q!ٌv'6�}9�ro��V���^�HA��0c%��Y���Tz���tj�nP�����g��
(���U6����h]���a���ǌ�<6�����]}��MG��I�|cR��H-䨳l?�`2�AL��M��򙨩���6
*�at?�зJ�$�o�kQ"�%��r�42��J�PZ_z�����1)�����Կ�@�i���|��&�Q���k�&3���"L���n���JFC]};
>���?d�����ag��f���z[ ,B��v%4�_e�0j	sT�i���,&^,2�g��'/o���ڄ	6��o�\rOE�%� �$ɼ���qhg��(�6�D���B��K�~ҩ���`W׷�j*_���_�K�X6�J䬡�/�Y�Ja�tO%���<%v>�)@3�㉖�m �a�I��N�J�eۗ2d�K��꛽�������I�Ӆ��V��]\ø�o�w�rqm�x���	���YO+�~��q����0�ہ�sF?w��ZD�������k�#'(��6+؀i��n��F�@wc����e�Rz=��Y[��U&�I�0(W[8Ͷ��Y��Y�t_H���PD.��̚"V���:GM���Al5�..�{+G����ba"�ԓ�+a�I��!��ʡ]U���3�T��G�K��� ,AJ^�5����1��7�N!]��&w�D≅{aaF������~��3ǃʺ�ߏ������yec16�^��E�5)�r��E��_�#��j3c�}��u��'��Lg�z��`�����;�
)���Z��t��=cvto-�L��m~�J�XNc-�Ƒ�2����$P{(�O2���Dq�6)T�'b��܍d�|�j��_�� �&M��\�d�@���f�`N��y߼xc�4��(�4�a����c���3��@3�t�G�,KS}�i쵍����4��3��K)��1���%��������%��
}n�9��'ɪa�x�S���+ϸ%��R�z�ժ4ACL;�&�݄S�$;���g����GGLKH���\9��Qd�Jh������^Dr�F�C���u�|���#cr٨��#߿h�t%���w�.:�38��?ٴ�6/yh��\Q��m���fG{�ƃ�����>�f0]�?#��R�����g��+g���˘�A��EȤ�b���W��Wt�ԟ�5��1���ӁI�vX�u�������:k�
��ф�w_.��ſ1b�fZ֙�͢�����c>4<s������9���߆�3�*��⧽�����M�=>�̥���A�mC5y��E�l҆�֊��5�5Q� _�$�}x��"��.�ZS?7l�ך���2��ߑ�Њ�Kpڍ�m����$h�X:P�=�a�j#��
��r�?��Lf���u���Ȑ��_������Ė��k��`�::�����CF�q�������-�a�F"Kc���z^��B��a�O.13��ڠ�k:��E�1A4��]�x��-У:�||���ۯ��<�d�o]{к�]tCJ�b��%���Na����q��K*���V5\�4W�ox�L����V�E,�hT�&���}�PL�y���«�̮d�.�� T |�Ș��М'��.�!�el7�?�������S�w��FP��m���uX�sѷPT��@<?K�[]~��݊��F�p�}4��*:����p	>�{�m����H���O0��
�~#�I��΃�E-_c�J�u?�6�Y.�o��t��pʉK�h#b�zӯ��]�
v���\��g͋���2ds�Xe1b'(�=p�=�νt���VH^�ksj�X� ob��@�-��4P����-��WW��|��_}	 7{�!�@���#N�=�0�J�WU+��	ڪ2�vS�\n�����Y�ja����R�&�R� �SU	iIT(�,?�"��v����/�l`�gky3s�(4<�e���H�%�)��b�;i�lr:�ԡ�,�|`��Y��S�Ϝ�c
>"5v8(m��n�YQ|��x�v	����V+�촖O�)�����.�v����	Q�κ���c��[�3�E��c?�v��C$��PP�YIYJS��A��2����l|~�G2�Ï��ܑɌ	�૫���0�%W^ɼi�� 7<�q�i���AN����"��,��H4�e�h���٪	��R_�cʌ$�b:�j��4�PP�CO+��=�:�&&��Ғ;ad7��􆳂��7�����3������Ӣ���v�;Ode�x<5���dL���� ���6_T7Qis(�P�.�M�O�	��t$j��^9�
��`Q2�;���ނZy��t�|fm�^nf����*���ӛn?�Q�6�y����,}v!Xkj�$~����d��V�g�Q7%�0H�������N/9�&�f�e9J4�a
	xF��L������Wr�f�0��I1�DPw^����+҈��<Ȫ��ZQ"�q�~�9��b��D��}�v_��A����kr=�_��d&�����m�_Q-���\�cd���V����5Cd�zʣ��^e�z5N���sf��[n9�U�=�[22�e����m}=�ǈ�H`�f]x�st���X��Ň�1b��=g��>t�6���V8�Sr��,I�n�S4W��XZj>H��j95}B%G܁��,�BC[�8 �&Yƣ7?�kߚ��<�xI��x(�^���W��$��ٸr�4�y�	T�Ay��vݷ�9�|��'����[�~x9�ߢ�9�F�Nrۆ�+�:[*m\6'�W�z��7 �P�@%4¹7�F�HT�o8 �㐷z��`p�������D��2»qVU@<�y��f�����<��|�G���X��;����]�v�k󵵬�"v��c�� �C������E�x���5���(*��p[+Q��꠼�X)vX��4�F/���'W�ʥ�I?��J�8�FK��O�Mũ�%<��!�T��������ͭ���T��dNW.�����X�'�\(�l���v�F����<������0�М�I��B�Vل(�0��G/ �V�W��f�3��@#�z^��.�>�)ԓjH�Ⱦ��J0�f��8<�g�Z#�.L�����｠a�(C���=h��g:�����_�M�ˣ ���'����de2�W����U*�2)oQ�W{�����~��W��έF�G���§|�=�_�b'��-p�ݮ�İ�9�����yW�*�v_�ҽu�t5K*�2���󡨩�����ef��G�貲�~Я��ר��Qgz@�AQ ���ͩ�ѐyy2�߯���rul��VzI d'����i_s��5����)�$wFZK� �������^����'�E�'?o)d��8��C�� :��!���V`0�0gq�c�0�{�2q=��b�������F)�ǿ�6���U�I�d�n-6oI>�h��P�����Q*zY����*?�%t[a�.�[b�x7.
�d~�(��jڌp�9���W�3� �y��!B6�.W�POZL�Ɛ'��`Jd��%U�ی{8��@I��W�E
"и�������w�z����]�ǽ���}�#S,T��p�_k����Y�㑀f�J��m��-NLO�(�0Hp��~�pU˨Y��Z��<�#u���V�=դe�k�>�d��2��gI\��߄�p�9����t�M�KB���^W��r�z�͠'�ȩLG=A��� {7
<�Z����Z�ڂ�d-5��^��H.~�í=���ə"�9��C´�U���&'�A�+�ք�!�m}6���H�n�6��a����CB=/������.�0��g�5#��j��7�0�/�m=����|��o�&2�*�V���5���1_�dQ7%��U�e#¥^�/Q�Z��V����`�a��4d��	.��EE�$���=
�%���sͼ���7tbâ�G:ě�3].�����f*N
~��J�6�h��xy>�%9~����$�H�ۀ�Ľ�#V2�K��샍�����cv��˟KyG�Ǘ�	���ϙ�pY�''���l��d#V}ZE�~��҂���һZ����k�	�G�!�M�>s�������#m�9����g�1/��f���2�]O�a�bb�L�k���9�*x��|j�*L��+��4`��>�ܾ�];���^�>��/;I�,u��C�X��Gh��8LEJ����]u������g!Q���'�A�w�_�^=����K�iu�hL�{ƫ��q0��[0�����B�L��v���.�FA}0�� ��@i+��=d4 ��O�z~���Jo����ߙ���qi_}v&���_���2��{x�W���{BX�,X��zí�p�R�ѧ=�X����NG}�_Yo�N��1/x��?TV�����Z4��XJo4Ҥ�a����Ir�H!��:�TK?�|���fTʲa�p��)�H*&�\3`��刻 ����]z�����w:{=ӕ�7ْ�>H���R���D�O^��S�%�܈�#Hjӟ���c���)&a���$철8vm���V sb3��R]���8��weԿ.�t4������T�o���]+ڶ8��߉�F��{d	��= @�JP�ل�aV
1�_�W���G��z�q	��V�ƽ��T$�n�����f��<Z�͎#�DUS~�ɓO�~R/u�2bq��3j�ox�y%�6��GHp�k$l�R�;�i��e]|}���2������/{�ab��t4|��v�M5����MpRMo�q8���|C�Gl�vZ��M������DR:ޤR�ř��m���3~߆��ʲ�l�}����9Ў���J���ڣZ���k����dy�6x]��071����&����ѧo�������� ����뻜��=�I�0���][Q�l�4�������87���-F����g�!��.�+
j�@ڮ}4L��&�Y+���l��L��~ȷ��mȀ��{�Jc�=ߞ*/o��7�d�0���mz��7�E��٭���}7vO���j8��g����}��]�������PZ7�����{�f I�@Э>0�ǰ÷���6B{m>|�H�}�2J���yͪQ; _����v�Q�R�i������S��NX��<-�Q���0˓ߐ?s�I�1-C��o6:��Cr� ]�`E�0~��<�|U.�Ԗ���1Y�^�Ra�Ps��*�]m,�ߒ��\8��ǫ�����LBZ�� ��j�2,բ]�5v����A<윸�>����qB��z��:�|�jx4�Z�I�:�Ѱ���Sb��iczNAmf��jF' (%�^��e]�Q/�.��0z����}��?19�M�X���n���/$��OUj_���%P~�����3Ǉ����,�C�_�O����N�Zݫ	�6���z^}\����A�,̙�˸:��1���y�s]Ef-�����?����$W���=�
�	���F�o�]��Kl6��u�֬�~�(rY�ӫ7l`=������y�73wO+�������[�쥛@��a�j�r� <�7���me�()Y>f��>܂�-�1�$���MmS�<����@>ޢ|�Q�8�����z8s�f�͒:�\�O�k���9G����2N���)[����J����P��/rjF��G
����/�R䎲i;:�1ɟ:6�pX���mo���{��D"���<�ִ�渓��z,��H1m�+7�x	/��x����m#	o����Q�����˩����ù�E�G����y,�9)Ҹ7��� �*��d�[{��B6��n��6,�������:d	%Ƭ���xU�<"&$a�
;�cz�2"����d�;��&���ﻉ�el����|������,��o�9��Z}큱'�<g�v?�D=��y�L~���@X]۪�$��?���.�v��<�۴cs�ڀ��m��n�_�1$p��T���H�v�a/�N��W����ϙ��� ��Ͻ^����S���X3����[{{�SM֦��P�ml�.���P���N�}�6�fﭷ��)�u�k�����vk�f�*<�޻�&'#B����G�֯H�P(1x����==��KD��t�DM�/�ǟp�r}ر,ֽ�-�d��!��t�"�QF����B)���ӹ�����<��U��%�b��(OXy2L��˟:�Pty'&���s{,�w�'��)�UB�+�B�Y�@�q;XI�Ak����0d{���ȋ5Ӳ�֜�ǚ+499�:��Uv	�� �ցYE��v~����KkdF22~��}��S]Â���[���Ňg���/[d�b��T~cM���5�~+�Np��x�O&��^wK��9�)9�����/���[�qⷩ�wW4.n�HA����/dԆ�p)�\&P�	-�=]��X-"�3m�r}�������߂4j�7g5�0����Y�v�'f���&QCU��lA��#��E ��ȟ�,l%�.8Z��j�����9(������w��4"��*27��b�f&�o�v�}���-?��{L&�oK%qe�q͵-��K�	Ρ}�-�$֏��7��O�<��{8��d��P�ҭ�#@����������������*C��Bw�����^�=#
��6����><ك�M��6�� ��H�vў��X>/�by���V�yCl8��f3�d8 ��^E��W���n�@�>@�[����-�GE-������T��D��l�c�?�9�O?_�t�3�FK�0�r�����h�KC`29���G�<��ў���#r�5��v9�|���$����$��|-��q��g� �O^���@#6ԑjx(�4���D$3�����V"l�'�S�b��j����9ħ"�zIF��5�?���*;i=����Pŵv���R8,��tu��܈FĸJ0Apjy4��w��G4��qvm�k�1䴸y(lsxy������@�3i�$M;�	F=7~�!�ɜ;��?�*nA��R{�X Jw��&y3�1����9<*��R�sz�hx:5z� ��qA ?a5�H㱃{��,��{6ظ���x�\Z@���M�=>_�p`��[b��u���SW?��O;aA����d?�����e`+�Ӝ�q�Z��	��!X&�!���7mE�Zb5��51�-���� ��#������Ҵ��p3�ƯX�!�<%��+�M;N1V���ǀ�W����/��C���v�ϻ�M�Z^���lԗ��UD}�l:w�\xf�Mk��ߩ�G���U�<����8N9�V����*�c4 �#��lNp�����Y
�o���$��vku�UNG��e���'
�W?�s���|}��{Õ5��pZ�i_�݀<�j3����uu~�� O��kB�]�kJ���>*�P��������a+��T+�tn���,�RL/p:��O�H�2-o��ؗ;�7�b4�*W��\3�	��,@ʥ{�_�%�"�e�͜�ƞ�����M��'��޳*>��cա���(WնA+t�Q�g�g�30���<�K?����}�T�)p��'f��?�� O9�\�d�����x��?�@ek��2y؆��3���)���n�1� %�w��|�N$c�]�i��+`D��h��]���?c�囤d��&U7���ڭek�c�E�	����p�4��0��1�f_�W�#�^| :�-��[Uky١��*i}�=Dm��шȊy	�
"~Ԃ16Ո�*�`��P3ff���D����l��	�/k�k���(�$�����\���%��ԍ� g7"���n$υ�	�|���vl8K�PJ�Q�����*��0�Y����S��.ɋ�!I".�$��ō��t�N�6/a9�D�F�Z/�S�*�����C���O}�/.`�e��Z�X�`��Ԭ��շ��0-��|1c�a��mD�Z����K!f����s4d�����.V<@I��[���Vx�eώ�˨�n;?.be������g�=4��W���-,%�#3v�enc7��',�l!�U�G,��Y���f�R-o���v3�%�v�_9��+���4�oY.�1�Y!衦�.Z0��� �a� 
«��y���چr�롅��ڂz�W��9K&Bگ׿n�r,�n8r�4��.�R�j!��Q+�ڭ��mz��B}�*����2��~U��;�����9��]xF4�������v;���E^��co�� M��ON.1l��0��%��f½T`�[�x][/z���/�׶<���6��fl�����u��L�>)h��BU��i"���0���`��pQ�Ұ˃OQ�b�C���@���Cʩ�fj��	�
��Sk��"M��Pū$�� NQ�鵷5/f��ݴ-`�d���8~th������SI���Ǖۥ��>�.!6���إ����:ۍ�.d./wL�Ϊju$I
���嫪�j��G�t������t�Za��j����L�"�'�GyJ��ؿ�[�o���̟&pTB�<���[5�R����Pe��D���3��[hz���Ҟ�����KW�)\.����J��f��=Fm��MMT��e-2�,����d���N�e��F(�%ϗEr�:+Vײ~�� ��P�*k=��?�g���v���1+m�����w0�g�7��J���x�C^4k\~�l��2����۠�M*4��7���z|�m���}q^�g�i�F"��ޘo0EU�Jm���~�d��uj��d�E�\���(+K�[Ϙ��/flbE�K�\L������Y�����R.r�9��{W�?@S�3�2��	4�
�M:wT?��9K�iLɿ��S�D|0 �fO�j_�.4�~�剫����=(�nG������NV��p&.*�|�UZ_O\U1��0����
�E���e��s:<Q��*�1�¿K��1z��O�G�5�4�v��s�@[W&Y�M��sk���%yĄ��t#��S�%b'���k�Q1��	�K�W��vb.�<�n|��͞;�c�W^V��Yz��z<���X��`�^u���ET�$
}�����窮��b�G�#Hx������x�왏J�����v���ί?#��D����?Ku��������� .�����V�T�`��澱0���B���6r����~ԓ�g���y���Q5Ɣ)Nέ��-�������lA�c?_�I����ӗ*�<��no?<��%T�V�ڧ���W�׽+�Û������(�}:���*:�Y�Q,S��X)z&�d�}�W��5���B�'�K�|kjk�û��1l���q|4�:�����`7UX�o��/�M-��Vb�a�*��S����3c8fO�}b�'d���^'oq�U�[;�=�(���7z<�������V�3��F���B��c��z������o�$�Ւw>k�w�h��9�����-�M�`᮰l����KB�26�A�zi�c�~U��#�+9n3<�c�Z岇X�*fI���6��*�����| v�}A�ѯ?�䡶�b��C��;��t�R8͠눥��v-��(_��\�dkC�h2�_í��ъ�I 1�y`i\�İ@"�=߼���w;��p����sL����O���o�ӡ��ݎ^Q���e74�@��Z�?�`�~�&4����aȄ���X�}��-s��.iVe�UP����P�y�.V'��K�_���7d���u���g�?;���7�c�:>Ҁ�=6C*l~����O7w���[*qy��O�5���T${���j66|5�`��d����ڜ��8�:8#u��]����L�#�ĹF��_�6od~U��"T�q�J[_y ��hb�}?��k���ɟ�����O��kkm~}���%Pg�5�|!G
}�X�������_t�F��������;�Q�nuo+%e��:3�}�/�a,P�KW�d��#��a�-tY���	=�w��kmC��]�ß�<����r�Km�̈0U���{_c�bN��,�)��E?�JU]7�N�:\���I�%۳:m�3�}���e@�`|�X��`=Ȭ8�g�bȱUdi���r`��4�x{QY�ay��]IۄC�9>�n�mC����|^�AO�v�W��}��(V\���(od<B8��}���2���}fz&��#�tʵc��|r�9!�W�
�;o�*��:��@=X�޺��C��o��?4]ePmצ�S��S��ݥ�C����C��=�[qw��Kq������w����nv���K�=3[��m�g9C7��p���u��r�S�h �Ğ�5�n;67y�ʹ�&��GE��Mj�sR;ZEXEdo��̩��79�x�4w��wtx�X.-,]��g��lB�?Dns�2=w�H���5>P�q{����1�Z���~��q4��7�x�`���fz���{���e®�A�	����|S� !�[�U���ǃ�m����]>�ϵ@���:kTc�����6�-������Cqx�V�会�/f�hs�8%]�������@ �[G˾	��UO!_;��VX���oRR��f�9��榗v��x�}�����2K��r(���x�9���:�c\оW:�L�g��`3ܸ↍�յG.�<� *���(��x͡�h��js��.XИ�G�������4!Q�D>*i_����<T��)c.���]��sH�RT��d}�i�B�G������w�xHHӎ$��l���Z��Y�����N�}�Z5􄸃�{�q�gW��i�{�:?_�f�K3wa�����*��
Eh��_?�� <�����|�l�=G$��3U*_�:�P� �����Lb�$�t�,9����؁�R�s��-��-a�h4k��ղ�ʅ�j��6��	�Ѹ�����t��d0�C�N%�>�d��"J7��eT�i��]����O `x�@�M~�\6�f}������rYK�����O͔�f���0oz:4� y�j����9�J��3�lbp�,N�����m!��\.%7�tר��Էq9 ��w���]/�6K�!=>�T"�7A�rj����?�*qFL�Z��M�D�1�cvx#-�x����l��~ ��u�Q�7�����dTg���O��xQ�
H>��0��5�1�~��Õ�>0}����a�5�~��L�=q��t��8^l�6}��|��	'r������;z��ܕq�p�d�Ȗmp��&���ͯ���p�c�'a�W���s���˚kP�˾-}�%l7��1�f�4j��UJ�A���{w<Y�1�;��Q=�ތ�w �g��!�`'��QK���8j��Wnw�����\!�ر��<��M�]Ǽ�����ʈùi�+�����gv4طR�n��D��B~~�W��Nl���[�>"xC��*pׁL���׮��|�k{rf�m��W���Ԅf���ק�i2���r��di�'_p"��U��r���-�XM��T�����1���N�K��6ݥ�B��C*�p#��r�����r<l��k��C�@awt��իW��^j0s�����?���}V��K��)�񱈷�w� K)f���ʢ�9���쥇�' ֿf-�ʝ}Nu�ؠ*�2���)Qwe��ύ�^����kخ��iq)ۜt&Xy�����Ԝ���<ЧR���ѧ��z���P?�Tvq�g�pU�^�������])����`?��<�����]�^��1;xy��ۅ �GD=�k�����ߝ+����B�x�lX���$��U[΃�0#Z.O���|��9!k)Y�J�Q�>�p2AC$�)߽.O����CK[�U���3��?���`M��$�����a�֝���*�X{�δ*EH�~]Ӛ�Ϡ�?� �$��ӥ}��M�5�\�A؋�l��ԛb)g����8���a?���L��8LJ[�v�Ѻ��<�}����3��#V���j��(yy�}��"�o�HQ��*�_�H����(Yi{�7��y��E�2����̾s�z�2��x��j|Y�&�7Z#v��#`��C�2�V�f�)T��������<��oND�U_(�U��Ժȼ�z�y�W����v� ��Nj���u�/o���0����o�	_o�j��͑W�xچ���R�S�Q�op��ݥV����m-.���2�u�@S��e0��:;b�Gj��_�꫈�#n��s�$�g�އ�2��h�;��;�m�U������%X�:�\�TS��|�2{��l"��9�qx�gE��w��qR87��]���k�Y�n�nq2"`��J+�q���h�xєr93���ħOB��=��UB���p�._�(�`�9-�^���ܜ�('��TH�6����m���n��)b7X��~���x �����Y�&�,�_���a��{.bˑ8����;{>�˓ʺ�q�k��R��>��v��#����9)�/��u.�s�_f�������D��t��������*��HA�;5��� ��ͧq�,�z��F��針�9��4ĥQ��t��(��0�b�c����U3��^ߋ3�LI2��Tp냻��I9������M,�����V�OgW�|�@���\v��WO�O\���XFXUD����=�4��S�UEx���N)��S�`�DEMm��5���Z#�q_y6+l#��<V�n=!�V�܅�D�xV�6֎����!��1�A��27�:��?f9�YoD7�Mfş�c���qC.�(�l�oӫA&�O���et"�n}:�ޛ������X�7��b�w������t����|�ͧɓ֪b��hq"�N�2]G�N�6ƨ��FE��e�Ὕ^{D�<9CzQ�O|X��ʴ.P� 0k�X��F�h����,�MX�7/jg]�%/�b�2.l����%_Ժ��w�UV�c.<-�z�/���J0��9[�\��PxMh���
w�
!Yf����O��)@Y2����ϥ�O~��<z� ��|�S7�k�n�r<�������0�}7��D�c�5����
X��n���ǧH]�dn�܇����WXZ��M��·.g�8Ey_���$�j|#�*�Nc���oQ�l�9��i�=6�J�-�љ9�iy������C����ɒHt�;�����\��I������;۳�3!����}��q�\���V����{�s�9���,B����vD��9��L�x@��Y_�y���36��k'������T���ʉM���c��}�F�g���j4�46���o�>w�� N������>@���;di�G���F�6�����j6��~�Ǔ ���oN�MݬoԜ�#\��K����+S��Es��[�+�o�'�a���A@�f����.R���Pflxy�l��É%��J(���lB�Pm��`#����ko-��/B���p,�X���7>��y�|�!����w�'�+�ɦ��J��a}�@`m��[ٸM��0���*7�Ukh35���}w�c�AJ�a\��t�M����s*9։��y��37���"7Ї��+LaG�eF��Z��%��z�]S1�E�r�"=��#�e�A?�y�H?��F1��1����MB/�љ� ik�j��ֱ�O��p�ӭtc�rn�7?&�r,��r |��#L)x��i*�D��x��a#N1��C�G����!��F+�nݸq�{ٻ�{`Nj4&���;ވj@tZ/7術l���&�:Ķf��7�䈒�E�-���,��,�)��CY|<� �$�	�Qu�,�����vS؝�	o͓ߵ��ȩ�0DuW���i�)�	:�*�2��5�q\��I+cI�-v�Z��#F����t)S�6mI_Q�m]p��������z>��
�GӹvDEo��˛+�Rr�k�;��P�]�V�)x�ukN���v����{5BUoCu�?4�Q����	��Zk/�)c��� ���o������cq�k.�;���J�ɍ3��|lvG���OC�Y|���@�g]$�5K�[`�܀C
"1Q��Y�(�4�}�0��Հ���CTm��R�>��S�>j���2=�o�(��H�򾿽��)ۙ�������V�����o�o	;#�={�ɡ�Z��p�㴔���B�{�%vg���}�����YO�%������� ~��h៮BZ��_��T>*R���d>Ჯ)�>� i�"�씚��1��;���rbO`Z�������R&�z�8�������u <��,�D������+N&Zw.ws���q�ڻ��8ӏ��P����c��$�Ǽn�+�
rU��Ӎ���QW��r�/���;���Fawq��s(�:�|LDj[\�����Z��u5�F}bGqD�/[��5ߊ���������N���G���F�>�R7��P��.g���[�R������H��"����L���W3C>4�xF��v��]t��m5'�핒j�[�j��O�|7k ޮ���W�hX�������I?R�j�>/eZ�)�1���CUC���$�9z�JĖs�ڇ-�w����,D�z763T
��W����b|�R)��b՝x���!1ha}O/u���o��T=/��E�xE�7xB��n�y���_՘�Z�
���&d)�a㫝-��Q��d:.��q�6�l�נ�'N|�n ���H����r��ohq�$��ӳ�����Rp
�솦���]9&�m�4��=�`t	}��"ug��ymZ�ޟ�u�qA	�K��").��n�O��Pk���t��w  ����G-���/�$��/;>�S�8"Fp��jh���T� ms��-�h�h���rt6HP�K���AF�G
�L�z������T�(	� sd�Wo>��b`{�Ĵ=�l�6�| >�2�X�塵��X˶#2������{�;�RN�/_H'�z,�!����3�8�eˎI��6�-u\�\�k�w#=JFD'K-?gb�+�Ⓑ�� |#����n75ڂ �l�Z.LJ@��1�wԷa��w��t���Y`
�>��z�#�Ǥ_?/f�~��x��`�j��:��c�=w?h�O�W��ꬲ�Jgtݮ��ʿ�_e��xz�����\b�O�{�����ӕ�`�E$�E����A�8M�*�%�BSph�s!�q�row�GM=�7,�y���&�pO �^���D�L��Gw�<���S��%�e���bG火R�Bw��P�梩]�UTc�+Ry���zeن�~C[N��͢��Qe=d���oyz�����J���;ԣJԭfm>0`GL�b}�����?T&��u1=h�f)�kl~���!���x�wQӗ�2`�A2��h&���H��@Q:Px�G�U�G�|���W_�)4Jͪ��K�<�n?ϧJ�fљ�"�v�i��r�F.�6���8�H�a꺶A�Z=���W���i�M@0?J�j� �n�s��*��ѼS�I�h92H�v��"� Th͜�"g��I�Y�^	������������j��8MSw��ʾ �zM�l �+Ĕ,	H��R���ڏW��d�`���\]�W|b|�1�b@�s���^�a�Oa%�?�����b�q��Zk/����.Sb�.��᮱.���)gqj��-���U'l"��� 4"�f�#�4��T��w��qa�ȓ�s��0-V9�0\�lY �캩�{	�$�K34O��'���cs��O"�[�\A��5��VH�>\�M�5_#�������v?�n.�H�ַ[���dI�3�15��D���9,��Ԕ��:y�E/`��[�o��������n�.潖^���+���Q�N*�z�#���rD�4y/�1��|��7ۂ�e��|�r�'[���~�z$�p�ޯ5j�7�5F����Q�)�h#��s�ye6{��/�{��pV~-�n��X�{����C�6
���H{Q��.��%\4��i�Z���s�"6���8^X����/�a~@�"�m�o̊vlO+׳t��5�Hw�F؁f��j�Ӧ�����t��hf������{Š�>������]0�G�ڌ��d`7X��°�x��ā_��cT�劗/v�՗��ȋ�7�7Dl��v�V��7�{�Oflq���M��a�Sf��@�q�g-@]ycz�6Aw�~�@Fe��	�i�{�_��Q����pqV%�\w�C_�)^�F�&6�04�1#�-��-�@f�`�o,�
���ZV=Õ�%�[�d�8��p��x�ؙȰ�Y���Ft�a�i(�%��^)��Tj�r>o�q��g�.��i��OS��d�j�o�5�ᄳ2���1�U��P��4�e��Ul�%훍b'x��t����so�s+�g�E�g�,`�u��@z�S8����gqv��D��� �_8�\���J}W�e�9���#�� ��C�x9-�׭�� 	��y�Ƹ.���j�b�>��w4��1����M�u�4�����u{�| ���*QU�v,��L��߸�4В�&�%�J���y��L����� k������5R��*T��I�[��'���sڴK�Dg�ܬ�2����jE��٥��,2ùے��ݩrĉ�B�j�k��u�@���Ew����Qj��^�B�\���/�䳼u��㐼/2��E���'������¿�^Ͼ<��������JKu�� #?��l������ٽ����'>�Rq'r{8��~�7�
0MA���N�6Må"¾7��Kr��~m4��v��uud$:E˭韉�_�c:t<�oM��<���r��'V���aΘ��:�L����@2?z���2mBk���V˝ŇYL9({\}����f�7�E���cy�$�l�]��dٟÃ,ٱ�y�P��2~���nBi��J���TF ]+��� �[��(k݈�8�!��#���NЊ��L={�"��Mo/_M��IHO�țm�#	}Ʈ?�v��q�o�t-����ꑾ��$t��U�>�RU�8�*||.�a�\ʪ��O	��`^h�̼�^����I�{4�*������q�z��tT�'X �}�r���C49݈z��Ҫ��w���z�_	8�&q(_��I�L1e�V_.F-�w	J��P�j�[R��FZ9�6�S��ժVۤ8hf��#`z�Z�
	��3��,9���~�"���lv'��ߗXrܡ)���lU2�]�T�MU�H��W�#�}�v�J�>O�{�+��ԏ����ã�YԚ�M��n�ȁH�2�I�D�����VYzi�,X�d�#f(q�c	w�n��Wb��}i��O��`��D��ϝb�[�)"߹owu�IϬ�G����,�.F�5*�P=��7}������vKL�'���k�R��(*�6��Yh���0}������$hd�*�x���m��h��&�{_�x�9WM�' �>���+\D�`x�@�DY��}�o�ů�ƠB�� 
;zZ�}둪����͗E�Z��0�ue�_Ĝ@I^��7�3p�o{��+a)�;R���߽�o����0J�5��bʽG�%M0���Q�,���Z6�A��g�h�+@s��+�[R�k���}�o!;0 ��5"�jf]ڝ��:ߤS���Tk�%�M����w�3%PO�\����Ϣ^5Q��d����Y���GE�)���N�2���+���7��e~���E����xR%r���ŊF�N���t��߄X�e�X9o���UBʗR��U�w�ꊉm�ګ��nj�o5\`�� �G�_iqa�V�����p��s�0|J�'��p|�ճ�~�+oJ��Ȩ=�d�݈��r��x�/:�n(Q���|�rpA � �b~5��˹,�����&Ý�� �?�{:.s_2�(D֢7�cD�-�����=�j�ً#��b�����~���|/���K�pq<9sV�ê�����Z�=C�����I��7��֏��W�;?>�&Y�<1��0�G%�?�o�zX׊�^2/�����W�~%�TMu�͉ì+Ê��.ѩC�8D�)Vj\��2�Dp�:��k����22�4E�[Q��ڳ��l���O�ztt]~rc�{��z_��`��y5�kHUOH�����$�qZ�C�/�-�f�\FD�)<!���,~$��y�f���q�*����R�����t&?�;�*�M{)~�A��ӛF����N���kS��A���w�&�>�e�������9��n�  -TwQ�G#d��� .��z�.������y���p���j��E��O'�PO�t�ZVW:[��Ӛ6�@��Ok4�Q��N�8�\ns��#�[b�M�"p��T�I5�,`����At�̸���%�M�'�)��Jk	�������ecd�R�����7Mk����ˀ18�� b�$�P�'�izW����bHW:BVD�:u�Z�i�-�~�R#4gh @.���VG#��ڿ����!�u��~7��)�Z)�o�H9���x<j���џ��;��xm&���7�`j~�Ձ56$���ڒVƃ|�C�y��peJ��߬�e��w~'ʿ�	SJ�Piv��9��D��=_�c�y|�S�~Q{�<R�P�p�����)��l3w��(�x�*��H�~F=�g?�-l.�㯻\Ru�n�c�d��S�à�L[2k\;��=��_��z2�QJ��=�zZrZ���2w3���X~�/r�hj�+��D��Q8��}{�A�I@r�����7Xņ�eٖ�:�bx����S��J�����n���P�谣�{j;f\]p�W-h�U���uhέ���k�d���d�P�Ot
����@kz�Z0z+Xj�\�AW/?��j/��A\��F�CRҝ5�n�%%۴ID(_�;����e���1�Pi�6��W�1מ�~qw�C�mn;�<���o\B'ػ�ד��d.��M�-�k��l�dr�H�t2�vi��c��t&�C�o-o�;�K>\�H0�[�� [���%��^��.�Z��]B:5KLw���e��bT�R'ghh֕j����7�So�3�΅�
�[r蹀�]�K����Q�MM�SCt^4H�=T��b����c~�Pz!�&K'N���ţ�*#���#M�X̋ޒ��`��q�d؉#������� �nHt2+���.{��]J��x�(����(�$��`���K�@��k;i�Pyw���J��^�Ԛ��x[���'}��X1�[=N�ۉ�p� �=Y��F�Yس+��p-�7_�I~C���_QI�Sp��\�p�Uۆ�[��	�dy��1�wz�I�T���C_֓�Ci��x#$��P� y%�I��n(q��m�)��^o�屖JF�����v��8��t��|�i]�a��NQ e�p���e�~��\�(��֡�=麛��O��}��P�a�?��j��$��0/�X�}9�fFwt0�K^�AY��gȼ�o"R,�ё)㟜�F
���$ԯ$9�f�U�YՃvp�_����;aֺ�)�t��U���v5������Y�++4A��dF��]������C_�9:�P��Z���v�;�� F#A�)�QO�v��f4�̢ɢ_c�B�VN �����d��n%��%�v�=�%U�LO�v9����{Dk��������N%�}@��ـ0yU�ݰ�l�ހ��Yh2�>;Prjį�p�_�.�CeE�Y���M��(�	h���v7y���X��5fF�i����`K�[�b���o1L8��Bŧ]r�ly�6ѐǡ(��2�Q��a�[8	�������*���O~�MN���E�֫�2K�v�vu��]T��*�D�Q��b$��_¸E����9~	�2�o�l�2�n��BHZ�9��#�Jx��6���x�rZ����̪它a��4�9fsILPjد��qZ�.��N��ޅ�4����8�&[��sZeS�<_fk���qqf���{xX,t ž�T�0,���V
��̀~�ｃ����3����>B*L~Mi
�5~f�F��T�۽��7W�i-��~������l�Ͽ�,o1�N�������oMV\�k����Ӄ)�j2Q��.��|��^�.�R����Ѐ�y��xig��>�������O���'��O�L�ڪ��S�ĝ�Ԅ��(cՅ&�Ӫ2�'J]U��^sB���6\�Zq2��^�>04xA�1��o~��Sz�M9���nudS�s�l~t���1Z���J��MYNW�ʢ�}���U��pɳǞ��� i�|D����հwe�WEz<?�Î��:@ϓ���� W�ǹ��R��s���s�|���}hL�l���0�u�z��Af/��Rȕ�ͭ��o���'ժ��"'�5���� ͩ���4�:����.����f@�E�rJ��%�_���-ͽ����}�f���R�@x��U���d_e-�FPbI�C�|^3�U�c\Qq�,YVq:�RLԍc���/+�V�^�D�՛/ud�P���D������Tݔ����,��f`�ylŃt��Ő����׮��=�g ^���ĺA.'~�w��yЙ���d�q�CZ�-<��i�����'6F�G@����S)��*�3�2,�8Ҁ��ʰS1X(��7�Ad��Q����J35if�rb@��o}�j$�S"�:�l�]|��s>*�xy�&��C�ʴ���|G �o�z�a�aų�p2[����*?���.�7_���:J8�#.%n�5��#O���$��+j�J�>�I�k{՜��v�_,�/�S�Ɯ#Oh4�N���U�^�2�4Fؾ��NَT�8k�on�N����D�%��i�	�Um��a�^��|ncHj�(�	�Yϙ������^���#�*1�:��?m��1VW���Hﯣq'���l�A������FOh�IШC2�D�~�w��'��� �JB|5�j@��?g0�@�s�㴀�S�c�������4�F�ՋJK0R�;������}�����s�[��bR�:����2�������ɤa�w7ş����0#:âT�1?�M�s��\�XD�����C��v����G�F�	HSJ��\�\=��}�]1hp9�y�l��@>(���XH�d��o�֦cw���F�M�!�����zE� �+$�91U��x�E�:fW�����B���萈�O6���x�ڪ�j֨N)�� 8��֠��ɸy��$�~S�����P{���_>�����\��9f��(xU�/�lV�_��Z�"| �9�6I�s0
��ҡf�L��u�'�Y��?� E�J\y�W~��;��Ւ���=���l|���}m�)��O���]���=dH�]m�[_�^_�1O�{=u�M��g�ng-�˫e.�7�_�V��h�_-�;}r�0_�M[	w;6�Fm S_�r�蝧µ~%�YUt���W*���xt�d1䞈կ~�<�ٞ��I�t:<��)�=�ݻ�I-5"10Ñ|f��|�����o{��3��H�B7��R��>5F���ɮR)gYVlµ��b6yo0�2:*�83�Kœ�3����!{^���$��fg£CJ ��FZ�wV��LJ��ƞɺ8q<�6lh
�P�R�ou�������n�顰���	4��#��W�w�4�
%M1Z �B�i�.�~�Ԑ�Z�h�"���;^��S�gƞ���b�c�ϻ�#��Oj��{��+ы-����?�U+L/�Z�`
�j#��9���eLU��K�Q�8	mM|q��b����+�x%g��r�GK�д��a?b��r��u����T�]��JnG��>�Mr�N��=��� Be������F����~͆y�c0�)�Eȸ��,�;IyZS!�ܷ5��� �9��6�Xt=����_-d/7���t��dH��PF�Icp6�N6��C	�/���vۨV�1��X�t���N}\*��Z$������|�M�8 ���!������^����}}4(�NV�R����KF?Y��;;:у4h�q�YKЖ�~���`���]i�34�N,�
7�dr�U��Ⱦ�^� 3;�e�&x1�o$�C�pc+[J��!<�cD����8��7��C�k㺆���/0;Cg5��=�qϦ'ޏ��3'�
��44�yd��g�����H�W��[?�ה���?��4�?��V��iXk�&U�x�����I�����T69��{�[�q`���os�iZ�<.��P{�΂N�j���1���_y�P�U��Յ���qb�ZL��>�7?ʹvw�|�9�:�r�A�η���K&����>'7�����d��]]5�)�]�
�c)�ަ5�8b	ݺi�o�c<���C"��.���@�c,;�t��.��_2��ٔ�S����A�������Y�d��aHZ@�Ȥ�d��64�R:���)ܢBP���#��N�YH��,{Y/R�v^��J{��>�8a�kqN<�xj�΅j�b�[��d�[VVg�j~x�p���N��n����`�L��j���Q���OdGf���x��jZ�n#p�AGLP�����S�0�]�y����N�R�{��5������4pH���V	�T�Z��Y+aR�tqૈ�?�HtX�l��l�e3��Y'��Rl�{g�0���p��n�Ѿ�=1��'>�W�I��WUMJ&�BW���JÆ������0Ȏ���j�#�+,m��D�ʗaH�q���q-٩[{V���P�&#5J��|>s�zQ ���V��6͒��eV�T�	X��G�wd���\��NF�D8Z�-4O���%��N����硳n?���k�����;�Wx8�'B`<����	+��`�Nc�.+� 1͸0~����.�����u.����\7R�h�f�{&�},�K�Ҋo!��'����)�4B;�_���e����������,�.p������х$5t"�6#�>����K���W�Vf�4����*�O��]M��-��lݏDW#Vq�mB�����ۢ����֭�~�	����$k���#��~�x2�����@*��nY�#I����z��)�[��P��bٍu�׈�Kwؤ��9,��c����l�?�6�z��R�)��(mE�jB��x1"���C�_M�KͰ�`�sѿ=��*�#�=�VL��Xދ���5��g$������5�f{�N��j�R��R��t%��S�Y��G45|&�z��`���x܊��D��U�����m�)<w��Y�e��� SP�-DqJ��@�M��#o6�]��W!��2�Mz"����K�h��J9>d_����G�����N<b]gzh� H��
�34��}�Jϕ�<��n[�K|q�vi�?��Sr�ϯ@�&���ml`yT��}��l�1]C�vrBk����i[��j8Dk8Grٌ���IH�
C�`g���v�8;��ڣ	���	���z%<^��߶(��~��v�)j�!��|n�7�	/M�|���_�����u���4��5�*�pvf���T_sOr�s���X�3޷�������م�I����͎d��o���{���Ajs�~z��ft����bj���M��s~�L��XU�b�-M���������u�䢄$���/;�z���|5dxe�*`Ɂ�������'FP_��q_��� a�V�_N�;�#V7��ˀ�47;t�TOrDn.f�`;��b4�u4���Ǒ5�%�q
����z?;��)Fh�Ǹ{,�TW%@x.�N�<����CNč� �Vd��ց��(δ���i�.��yг��� Ţ������� 9�~�3��on-���� ����_��FH�M_�y]*��pDn� �ů�?�Y�I������L)���]���kU�up�OrA	���-�U�u�%��p��(t�J��r{}12��H 7�Fs���e�`˼���l��&�������h�"v�+>�"��2o����C8g�Ø���*2�pw����0���)��}�������H>���l؇,	&͊	FT�M$���]-�ƨ�k�	�v*��|S{��d���I���gn��f�)^����W9=w$�&P���O$�e.?�s�������v87��t��W'��٢��i��IҹM��m�g�ҿ�t�!,����{�kx�9S�b�h~�:9m�QO&!z�-1�X�.ӎ�R2�<n�汊@8�{�N�����=/�����t4FY&M�O�(L_&�w��sl�J����� Orl\\�Ck�� ���jJ�W�X{���*���=Ǻ9!x]I3�F��/lO��v��\�\�Xsge3���'v����K�ϴ�m���ז�I�d�
N�kz�h�ƿ.�v4��Z$C1��2"*��]�i��]�!1}���*�11�i��k���zn����X�� G�譋��������6�C��Y�C��k�o�K
t���x�ӡ�nu�<���u����-����_{�'��FTᵆ�``���X�+�Y��y����ݎ;�a���FNF�b�Y��3϶���-l�?�Rg�7vr�F1Ae��>������Y�Y���x�ٙ�Ն' �o���rEQ�fkf�RZ��j�K9[���syS�
0L��i���`�Q/��5MD�=���:�p�0A~���Cc�dS�-r����T$�<+0�)%+�â�$��b���[Y�
��OOg�$<��8�B�)���¿1�KZUmT��;�-�7f��"�*;���;\��F�[!��-���,8�5ܗ�LI�Y�"�h����ټ(��G��au�u���
�0ngm�2�-�s����#�4'��e���׾/���c���Z�V�j%jS�C���!Z�=S�X��2��KN��`I���yO�zf�i�L��A�eh�����-ޔ��j���3���%Ņ�f �ߨU���Md��d�@;Y`A���>�p' 6t�e�n�a�<t巙�޵ޣ���+J�W���ÔJ_��B��>I�R��*�����>(��z�G]z�����@DI�$��:���4x�,�9[/�%`S2���C��ި{�����_w<�6P�A����6��ߛH�l���^S2�����u}r��A+�{����B	XT\�p(rs���?<�8!T��mӢ�rt���
Sj�~k|���TpB��_o�L��5��Yv��>�:�ڼ�ڊ��jW.2E���}�a����Zh^Xi��b�QU����_�w�]i�,��S�_��_��0��+Z�S6�{NV�v\t��F�@�C���c�r@{���I0����J�?�e�?�DCV(�<���R��v�U9I៼c��zS��}��������!�j�g�+�}�,a�{8�����}��Ʌ4'�����w0Wu����C�17�@�_}I��K;C$TC����\����׫e6RCf�)�ߣTܨ�=b�ie���kא#a�M�T��t_M
%A�g�O?�_��'?e]u�z�"���<a)%Z�'	��(K[�I�[z ��t���ާ�Ί���d띉S�2�.��^Y�|�[�nY�R|rDowE��Ր�єf�-x>'VN9�IT�Y���=h��q"�L�:�QB|��Ȓ\���2��=�L8�v;>�;m�׮�Ԙ�w8B�8��YH޵Eo�����3c���u���7 ���~��55�-` |u<���N���5ғB�ɇ�k�N۽B����k�s��!�]��l��A��������k��4� D!Sv��F9S�GDt�96��R�БCu�hK���Yw��cI��p9�]����]����I�izE�4=A��6��3b~d-'��Z����c�����%�Z�������x=̙p�-�db�y�<������փ�>ެv�Zn�����@1����	����͛��針ȣ�J�'.��_'��Յ��e��HKہHV�ؓg>��|l�Xe�К��r2�:5�ϸ��ء�*(��9mgMkx�0��c�V�%��Rp���(��g (�t!��w��g�,T�߳&���[�nam "Q~M^t���.�.X:�>S 6��>���'����j^�N�J�hS�b@�e�`_x5�Z
�>:m�� �?�Y6�}����f��ͪ��3�,g��v�9�h�� ^�RQ�|TZ�{��Ԛȱ��Bd��ޝ{��n� t%���%�ő��k��g�<$6�j�h�U��F��@�ι$X�d�H�WN���s��ϰ���J�'Q��2�2�_�٬�Ao�f�~�G$'�(I��*�I�V3n9ɮ���`H���2��*��|�2[��WB�
�qp� ����h��=|����ϰ�t����z�J1����4Y��6�T��`��ꑡ��6	]�I�##����R�[{��Yj�>�VN�^��:C�=%�!��O	�(k��&Q�k�����Z�+j7��/o
L9�t<�_WS9��9��YK�<�SL�cb�?'y���u��bR��3!�4��m5�#ˢ�8Y2���7
�]�O�y�-O�]<p
������X�� T�kK�ң��)���^��>ioOj��8�V欆�i��B��dK��O�7�AF���A��3�߼�|�M�{BP4O�l��*ޕVO8�#-rv.�yeh��n(���&|�_te�\�-^�l�3�DG�4R3:��|9�¯D@t�s��?��o�:(l\m0ĻG��8l�p�ꃖ��ܗH=���`I��Μ~��⣿�*
uR M'�:��͟�TQQJB��bQS���?�޲��&h����	n�ݝ�������	�$8$��;��w�w��<_���G�5�]�UW��=�ȕ�rH�RP	)��������u�E�V�`I�,��r��xx|S��ϣ����p��S�^���-8���4��>#z����1U�LB�@h�N�w��d�g�P���=�ZR��6pӝ��#�&�wԸȦp��K��S�����=�?!7���a�3$��q��Y*�L��	����i(�R��GW��d̦��c�?�юf�:��@�[��է^�뫺!���(e%*Uj;V
��99��&�LH�n��+��(�6��P����T�:`K��)��	T�ꕢ��{�k2��ynQݘ}^�4����&F�������i×�9��S�����9�Z:�}^�쟛���x	a�'wr����\������6� ���"���R��)�"'��e�L�����iq��#+��Cߛ;#ܛ{=�������[�\�|�YI�|�f�O���A^�lU����^��[հ�t�2����o,g�j���EvuD������Y�����t�/���|��o|�g&�<jR�2��ݳ�I=��0A�����؍@�;��o�Л���4љ���5 wT� 	v�ְ�}[���8F��{ �b�N�d��%���?�e_�6�mSYDBT!�n�D�9ɓܫ�}L\�i���Śk��)"���ǉC �E�����)�jkJ{�i�dO��5E��ܵ	al�ޜ��1]�b.��E� ��	T�{��<��M2n�u�u�dѯ��E|1�`���M�k��+����!�#j��u���1]������B@����)w�a]�}�F���:�����B�	EzR�}TAE�8����Љg#���A��u��ɘ���]32��h��yl�[HpҠ�7�p�fQ�蹪6�� �R�U�\���G�C��}�ga�+x��]w7���_���PϏ=���]^QĿ]�|E����-H���-��G)S���r�
�8���}���7-hYYS/���em>=�����]����֞^�����(�Pi�n-E#n���<���d��9��8;:�JI�N]*&�H�Ч��AS'�.��Rs�Q��Rs`���>��P��(�f�'�˹�������q!M;雁�4LfogB)f�Ţ��Hn��p�[�RoQ�����G ��rך�Ϟ>�?ss(����wo��+QAt����k�!�x�n�l� �^;[���Iy9NA���e��T�^4��=���6���Q׉p�����Qq�SՉP7�At8o��05�]�<�aR/�l������N�'�|�R�̔���ڛ���P�4�ɲ_J;5�C�8������&�q���2�{���K^�������?�K_Ï�W����8�_ecŚQ��q�o��"�'�1[�Y?���Z����~ї�����ls�:T�,�J*̑
B`MX$�Y`�u׿�^�,�!�^��b"�'�,��{l;��rPs���ߓ�X��;��B4~\|��s�����6 �ۃ䑚�BK�J�zY���R��|�cq+3���Ci�����W$���r�!k���aC�0~����z8�|�ձ{�]�22��^�ƺE��sr�M��:Bɜ]��:[]zz)�e��o��:A�W��m3ȝ�Э�j�M��u9Ym*x5FK�3������ƒ	5�h�ʇ��V>T4��d'���v#}-�w}�`A��ts�Ő67���c�V�����C��l�j�p[��
������d�1;ߒ�L����?Rwެ�E��u8����y�$M�l�s��{FX�����xp�`�sJ��xX��˳�&��?�Мq���6���_��~#�����.��>��P������ϟ��g��,C��c�[�^c~����׍]����}�}*�\��H��ͣ5�����:���mu�r[���ࡷ{*UV������&d����K�����\1���c	�#w�*zlһ��7e�0.�����E��k��o�Yn����w���!u� ����H�5|!�_'��`����AW��.rv]��r�S_���ޕ��ݩ�u�n��Z$0��7;9�Ի�[�H%��*Yh_��{堉��w�B�
��5�4,>X!D,/�^��'�*O�t����Ŗꃡ%���?��S!Mn�����FUX�����W�������m^���u�b��ϯK1I�����hB�A�R�fgÏW�F��{��;S���5u�1(��O���	���=��&f�lل�����_ř�'�q*Qa�͐���c���y5=�1>k��*F��:�P�1_�(Wa���������I���=�u��~�qJ�y��?���N)!���E���9��@��g�`�����=�a�W�5l~2|iJ'۴,��=��j��e[���C��J�����n^tH����0a�!S�v�4@EO�P���eҕ̙��D��ڰ�9�J��.	iN�K%ǀ6&z�k����s�r{-O3Q�e~�O�ě]�L��B�jh�!ň��!�E%N�A@�̕E�%"+���S��!ߩv��t�~�(|����Y��>?�����uځH�f����AP�%q�)!���[v�;�a���vW������.J�g?�r�@�-l��L�/F���7�Q6c_5h+�+�%��ͤ��zv0�$o�r��v��]�57���Ю<���k:���M�ߤ�]���D���҉�VX&�BD`GV���	?��2��wL)Ks�q(��T�u2�X��v�6��Wڟmj^&��i�2��~��e'������
|���wz���Ms-'�ߩb��Ur�Q���l%a�JhQ�I
���Wth��폮��N�*;��*͖�p���ҟH͞�0B������q��Pm�a^#I��
�qs&�(\0�?�L�ֶ�Y�$C���_�f�gr0�1�2%?��Q{���0�
��N6b~E�͊��=���g���P�,QׯU�<|i�J�?��s��aX*��}b�����u@�&U1�@�PlB�@.�26���r�q����^�0ňÇ��������Z�uZt\��^G�}����h��~g�i���{1�U����pʚ�6K~�����d��0��J{���Ђ#+'�Y�S�Fݮ��9m���M:�,� ����c;?	c�@����R/.�$sc��x�oFA�j�O;1��VY��z��}�_t\�����52D�����7�|<���2]w�Rn���j�Ŝ�����:89&\��2n��ǈ��V����T`��th��ա7˄r1�/�����M�s�l1M&��gM*�|R�{Ć^��1}�2��}��l�x��e:3\ݱ,�Dt�l(�)�qw�����M֓9a�����_�����Ǡŝ���d �A��B�!Y�MV���R��Öqv#J�Rb�*����Q�~��~e�$��W�1���8�R��<��m�|ZL��Q�)�j��/1ܱ�Io3ʽ�A���w� h��-�/�g������L�3��ܸ�+�HS�Nh
�����/�v��2�����i}�g�?�}��EunAc�3���5��u9P���0�Pv�_@R��#�D��]�qY��ۓ;1jrPw_��y���S��6�tZ�I��0Κ���ډ%����#�6H+.C4K�-�V�^mٝ�~�6~7�@�N��UB�2q�,���6�'}���/�d�@���ƃ{~NB��qڟ��K�J�Y)��+��疶(C�.׎�(B)�Ag�w	J�ɏ�iM�BP���Pb�2s�Qzq�>[��F������8������۾S�^{m������� {�Q���8�jN���$=�M$��H�8���ݷ�T�=&������Ze�5_L�R$�#U;v����޳����/3E�򽧤	��.�W��U�Z�@.��J�8���.���X���JH�ӦNa4R6����$�3z�De*H~���jzlk &���Kn����������nA��Hׁ�nvc1ͅ�������凁�6
�� �����e��*m�9w��!y]=$�1��T�I-
p�^�z8b�Y6�p�d��h��l<���-�싹�3BM͈�.TM�%-I��3>"1��Te#�A�'S�v��>4�b)�\�l��o��e���4�������d�&$��������h�pK��630�ֱ�12�rܞ?����ZC#�f>��W7\�M�i�1C�
.Bo��+&D�ZhX��ZIO�(��1z ��kv��m�{z�ZE�/��	���8�P�ƛ��hbQ;x%������,�_�j���%��ag�V��&������Μ�/�*]
�^J�6B�&�h/:��$_�G7N�q����%$d�֏VXS��%�"Li�z�y�v&��,�b���
ĳB)�$J���$������~*ۍ˅�9'���9G�=�W&0��B��]����M�{1I����՘x��~_O:�O�P�#��Ρ/ݙ�}��d,⯇��?���iN�5r��t��E �b�~�$,G��
i_CC? �!)�2�%p@��[:g� �Ӊ�gF����Ә�eO�jm���g7Z&�:�8 @"���L���C;�}��N^B�JG	�i��#۝� y�l�7���b��T�Dn`^D 2�p���`��r�	7�*}���D����r�p���J�s6��F�Ҟ_z��Riv���0�8mL��a�� ����8��"�!er�mwi�8��>q�tUa��Sa�Fhx�n�S���?~�b���bj�Bjh��`����&?�c|L���n���}2�G0U2"qEJ*�5�� x����?%�1yLk��xp|(>(�E�	�����@NQ�yw��{�6�R�\��^��\� ��K���G>�En��|��*�+auzɮ��Y I4&@a�V��R]XɋmȔ��$5�)h��p��p�3BVM�v�q>+�����(bf������[�n.is�`���慻��'�Q��B���B�'_����y�%L)K�[Y9�G �!a�5���2<0�i���YWo�f6���ʵ�L��Jv��y�M�0y�+��Re���26�n <'P�s>���(i��BC|�'�,M]��w��1+"'5i�E��z�B(rt>�ަ�m.��2����Ȅ��x��T�q�5Z-����,��`ѯ�Q�}E�ƆXG�T��Pn�E�}���8�����ᩱ�3��u�V�eK(�BFቁ*��[���n>v�#�x���W�Mţ�	&��*�����,���	U0��p�΁�DEŗp�} ��$ ���6�п���y�dXd��<�a'�䈺`��Gpg��c�0�ap���$Ta��ɼ(]�2��%��K�7|�Uf2�\xO�ݞ/s�R�_=ϔ��k�XE�*�bEꐅ�cG�x�-���e�����22J�}Ā�ʇ���b[����$v
sÁ�CzXf�/ϕ{�`<��$�MG��i�1����v�5�?p�0F�M�)u��<p��4�V
�|u�� ih�؎�ÐF�����Rs�ӆ{���E<q��;�>���"���^�Ys������s�6���rnTF��:��������pQw�
G���/Ɯ��o�B.M��	G������հ���������
���h��N{Ӓ��0�Kb���و*P���n���s�|�K�q����,.�	���pʠ��ī>�������LJ��m��E�H�Nu{2���0�����aA�Q�cL�f%(M;M��l�Z)_*��x����u���l�}�ѐa�R�r2����2�T�К&r��5���k�����U j�9���g�I���Rt��&j⎋�߸i����UPn�����d��ܛ1Qq�%�R[��-|�D�A�s&m5��[�y$x����&s(z����ۑ;�dC6pa?"H�����=<���K�Ώ�k��.��G�f�w$T l2��&e���j�m0��8Y����T_�Q
j����K�L�͓qf1���D�j��d��j#����O����J��`��7%�Y`�.�[�$a�[2:��tݸ�[)�fqrA�?��#��=A��Y���4W��Ɂ���6����2�	�/=b�*�a]?E�+�"�LV�۴�.W��������I%\�����8I�p�\���`v��NR�o��۷���;M5�=[:�JB?FE�,
E��^:^�DD��1z�#8rtK�8YP\���G���:\�W��	Tu��ۈ��ol��1�#+t��k<7�T��v����Y'C��_W�®�Ųn�D��20�Lx\{F�:�Pi�s�E�&}�1fn�)L���z���%pa���I��&U��{\ԡB�v�/� ?�@C���"N�e��'�8�,�D7��[W������4�^�Fb�&��(�>~Lf���S�099y�ݸ�>�a�h1U��c8������{!o�P9>}V�,�՝��l�m���i�mN[��VT����U>�U�����;::z23G��4մ=ھQ$�k��o?�:�ʪq��2���m+w����mИg$�j+��_�KHT�II�8B3�����5Q��p�q��p��7��V\w�l;U����Îp�@��R�5$��vd�za��@��r��2��]��C���V.���6����A��?�;?Jn�:�U�b�L�^�B%��N�����n�(C��m+���� ZWA��1�㊋�����&妁<��H�XwF>u.|�ic)��dj��_&M�8Q�Q𞤹j+y�!k�R��Q��,P�}d�q������/�w�6E�܃����|���?���u���A0����߈��o�D������V�?�,[��se!�j��\����?W&Cd8��ϕ�`�g�o��7���Aso���?����e���H�9N\d��G�B��V�Mҁm(��m�,�l���m.Ň�V�-��ކ!���@�~5��w��0���a��_�Ԍ�Cf-��� � 4���9A�A/K�+�S4�P��n�-�n��9��9Cߑ��b�A�e�A��vo�A?*'�:G�p/��.���?#��^�/��Q��fy���'�ԇ�j�Sm!���{u�3�=�$Ţ�V�׀�X�cm����HX��0���ͯ�}v�bE����\�S������E���z�QjT���D$	�m��!�VV:�zW@���)�(��Q&4*J����ِt��o\��d`e#��o'�!n��-�!e�c>ټ@����G]H7=���;�#J�F�dO��ŵ�@�Z��M1b�c�%1�ax��8k�-^+%�����iSP�L�v]R��w��uU�$9`z���ҔR��g�E���hiW/N2]�H��7z��p:�F����W�=|����t�0���%��#�hwXْEj��@���+���"��D�^��4|i��Fi�j��̜��鶚G_�3J��f��+]�[�������u��jm�a�n2|�7�r�`�Yz}�O�1 I��,4�*�-4��0[��r��A�3�

�7��`�-��L��3$�P�Xk�s�jp��0�2�ߊP����B�������f��D�mym�r U�bCZ��T�DP�@����m(h�����t�ʟ�l�>��?�˛d�7)�J�FL��6��3[/��F��<�{�J&����ӹ|�>7�dR�[��¤�I���Êj;l���
�<��׾,ա�P���'���-���.����?X��N���`8y�Z ]��E�'R���d!>��/&nz��:���cTj!�;�YO��猌�[ؿ5¼�U������بY��{��T&o������v��a�7u(���:8�{���?��R�g��z�Q�Ԡ��5HP9��7<�H�N��=��!���>_��\�U���k�iT"=���s��?�m7OF�˟�j`Fj���O��fA�ڌ��iM��z:����B�xF�|��U���F�}�� �A�JFNn����mX�t^���1���CR"i}�Lf�ha���z���6����i�w	
L��t�����H"��q�9	iT��(�z��p�k�*=0��Nd�j�a>����������A�f;)&^>�0
�+��FXl�
�3�ϐ�ⓜ��%+,���&n+�&�����-���*ؼ?�9�I��rAQ_2�4�0#I\��W����kNz`�7oN�f�G�s
E$�K��N���� �ߺт�E��S8Y)E^�
�A
Cd�	jytG��(E�e��J�=�QL23.��Y)Pv=��=tv^̴U��gY&���X���Tx0C	xP�X�;+ݽ����K�D��~����� �P���m��[[ڴ+��oneAo��W����j������G�׏��:�^�xM+,7,�����1���.�;W�g��?(��E�lC�J�C@��]�H:�ɉ��Z~V�Ej����#N�<��l����6U$"��E���M14�Ra�YѸJ�����4��5���pߑ�@	X:3}q����Rj��A���������7��֝Z�vaL��{;�,{8MA�ů�%2��������{@��-��� �3`Am|���Q����c$i�K7ژh��|��uK=�|Fd����Q-���}��{/�P�x&�7�����%���M�{GV 53RY(SЂH��f-}�1��"�wZz! �z^�b|$���O�N]�E�')���g�R�Gw�r+)L��r���I;H0���,�@���4�j�9�H'r���� /S4&�zh�:z�{�V>�K���p
�qR�^1�mkJS5�|rWz\�P����N[l%� ����G)���.S�m��Ò�H�A����.܀��iZ{��6I���X*�O��w�.E]�M�rpl-s̕'�](��R��8
�!��⋍!�Cn��7��`�����9��7f`SI7���'d���Xͼ�,��lVy��'�\$�V� �p��YS��G�р�Yi�{W@92u����%*�#��д��lݩe��`K�� }��X�jɒwg�z6��r�lA8���ʕΪ�=��8-Ԇ�G���H2�e)��q/]��
�k�E�-a�ʇ���!���D7�:ŕw-�>Kn�u��^�F�W��hv�Cn�O;����%�/�^���Gy��~od��_9����3ؤ!��Fl^�4[j��<g��`��)ڙ���������}�_v.D�B���f�����-� �8���|tԐ��M�`k;������r$N����i���C�v��P`s���m,q�#P,y����f�2���w�(���_��T a6:H���$�B��j��R*_&��JY�����ˣr)����D�A�u����S�W�BL��@�5��4%cF��<�0̩��mIן�
˟=�^�;��7mT1<(��[P��<��|ީ�Pϸ;A�k�	���s�r��ZV�d:�r��ľ�ok<PE3E�Yes�A���dR;�"U�;�9H�t�K3XzT�qD�w%"<�$�]�`�[�N�@�&G�_4fu/���f���0�� ǎ2?���uv��{���u�GS�Ƽ\Q���7��"~�����s'
l��G5Z���J--���s4��´#YUN�+$=�ϔ���MI�.���l�E�v{mݲ�&����Hm��>������bN ��t���o���Ċ/�#F�^-CͳW��s��US���p��A�·v!��0Jɔ�uc�	���;F޴��,��Mu$P,��%�(qN��&	R�J��}םH�°��H�zrJʩȱ� �"��v��$�@I�`�b�����{�Ii�/�'�q�+-`�âj�/��A�9��^��Ϛ��^�0)��.&������)��TB��ͨ����0@1GSV52��ƪ)T��D��b�����i���Qh}�v������e��{g�Tv����C��B�)�|�{�[��]E����=��w�PV��I��V�&���}Oz�i˥�"��\#�URѐ>�6XӻE�D\�(��̵��KE��w�iJ�'�kq@�q�� >W��:[v9���N��\>�A�iJ�����M�����fV���_��I;��*����x�ۛ!�dWJ��"�1������z�n�:�n�"˸���{Ov�����l���&����<�&�N��S-���R����\8W\�]�~���[�O>եuъI�4�ʯ?=os���9��q����qVy+� �}z'���q\-�
�8��QQ�cYJ0���Գl�vz��S�	$�/z�~�����mZu �M����]f��F���~
��j�G������ D�-Jt}�e{�9��h�S�.�֋��R����?B�v�<�n�l�xA徱���X9TCS�̠�Pr��~��ϊJ���2��Z=/�Bx5X_����/������;y�E���8|:�;���zЀ$&�r��LF�쭟r�Xx]9(ծ�P����m&[U��_sI�~�,k�n�T�-L�3ඳ�����	Q�Ɉ�ܰ�4�h��]c�76b��\�k_�(���i�t��5��qÕ�}��s��5�t�rS#K�8�P��YU��>�Ջ^���I��<��X���}V����Ե�m�NT6�z`�(ㆮ��W�h�j�k@����ǋ��Q](���wO�7���'�ݬ��4O���=���(��~��ـ,��ds���ߕ��fu�5?E�rٰ�շ�D�q�څ��8��η5^U؊?�~f���>�!Q(�CO�,;R�>��ل�T.(��S5{&s�w��;��}�}iL1�g�8 s����\D��X�P����9r}���u< J�#���%T �Ǎ6b�W�0:�bʢ�� }e�CA_�<̃�s��߼�b���Z ���RI������|��~��U���f���2�������C�!�¥�~��40V�v DW2U���\���^�X�{1٦��o�ކ��5�&l �8��%Qsm���e�����y���?�����Z���������(����g��u�ͨ�{�I����U��p��cz�*>ej3��	1]�s���)u�=�,��\���!�ݪ�Ӿ�[�5���FJ^n�04��u?,o��U���IM4���o΅��v�+�Q���0��Hk����K}��{�_�:��k_%F&�s��Z�L�ue�5y'�T�P�H�Lgg�p��ױt�֞�ڰ��>T���C���u]̴�%}�^��e +}��''�4��k�h�b��W���=&ݚ���|��pl�.[v�pn�#>]/C����z�������.!�G`�c)i��hkH�6?����<~Z I��:=N���O^�rC@))���n�����T����*+d�z��*v����3~?z���v7p���G:��t-Jƛ3hǘ���|�j���@4^�*w=�=�xG�9�	�������Z����뮎.>���*"����w5��#��-���ޕ���q�>�0i~|�E��e��zRz�q�4�O�Qjڠ1��ן����Z���$a�&�[�$�L+~�޹���u�.��^�C����Q;�6����¤�#��\Al�$�R�Z������
��?�NJ*�bQw�
00)ev�{��ӪW�v;�G0I��޼��T��1-1h���\j���)q�4Ӓ�z[�?8{��?�!y,]̒@`���<�ZB&5�0+4g��T2�[��9��:K�Dã��*�����نW����%�=AP%���̓�b��5����.��++�;'
�lh�4H�,l)�{�/��x\?t�l��#W@�T K��( �/o�_�5Z<I�ަ���;w�S�Rcqf(�;Jei�Z BM
�.��$��s��[��Į�����u�6�[��4���LQ�BSG��&���=Q
m��`@���3�b��K���C�bO��f�H�o����2����'	�� @��49T��x�遂K��E}uKv����k�,6��E"ڲ��	�V�vO�\��V�CW�U��E�("�şj�ۥ׎�]M|�ZH�;�׸�^�Cj�\I��hDE���L����I�f�$c.:�:�&9���QW�N�ci��a*��T�B#q����+b~5w`�avoX�/������j���6�{Aʡ�1�:A��ex�K%�C[bL@��w��xT�cNb�չ��$f�},wO�LgT=���q�� �]|�7]P�̏�9#>IE&ru�{1���f5x�2F�W�w:���S����N�m�������E��F�}W�w��3������x�Tt��,�Є��w���Ӛ�_���y��<LMU6�W�ÿ9�����x��f���5-J��M���*�����_DlӞ�(|ö?��ȅ �I�VH�JCo��Y�F��8����9�-�`��B����r���B/�T�5&��~�OnE1K�q���1N�-�X�y�>BWW	]":'�\:X�<�>-�Y;��z΋MVBCn��T,����&`�k&�Cw[Y���oq�_��0u�Tʜs�>�)q%���[�AS�D��3��g��&���b���Y��0�:�`q5�u:*5���a��8)�u_z�ār�El��ȋ����"�>�M�6)��;�����|ok@�|E�s <@h{��X�01�Y`��v|$?��?U�FB�
�YX��� C7��j�r��8����Q�F�B0J×�F�қ�����W��k�Ê�+�qr�Q�C`�(��)�5͓��mU"L�~���	O��]����o�~�c���{�sa+"������@k�0���tT��
��_�E4�ܬ�i\�®whW w�S�7�����o��x1_�l�nYj��H+ڜ�� �F��3��:�!�ب.�ΤGw��Dym"-��\:3�ˠ���[*���$��y#�׭�?CA�(��f;����n�K��i�fZi��h�קf����
���)b���#�I����s�b�@��a�q1�5��h���$����*�m�J��1c
�-+�T��]Z���	���K��J��A�2�1w<4�02�G�I_�+�:�V���w�8ql�EU���d+�)���Q"�B"�
���S����Bt�s����}%��s�լe������N4���o��(q��IwNP`��?�� a�A�+�V2v��e�fI=/�լ��B��4�[(` �b+4�K�f��Ca����\V���2������(�=�_�H$r�_"��VOQ`K�?o���~C���}v��s�@�l#bS�0����hK�L8**�&o�nt0$�PY���xċ���$� ��Kئ�c��*ES��w��>\\c�����4����ִ�r���,���h����ooj�M~w$�#����_�*+����.�Z_6�Vq9���\�ԃ�()K�A|*f �!I����҆�G#v���uk?N�7����as���Z�z�'�<+g��oJܚZ?�4����Q�L�U��x����?�V
�m�;
m p�����x�P:2�U��{x�H�KV�)kO�h@�?y�-H A�D�0�G��k�ry�y��(LAF�nv��6�M�F���?Sy�Q��e����:S/? ��������q'���X�����{������|����tX�Xq0\k�x�H��z}�y� ��g呚oE]�GG}���J��	7���\X���^Vź�阀��_ǜi���?(�H�M��O��P��c����@'�T����襸�{6�R���t{����e}��+�v}q��n�U ���/��ߌm�
�pq��M���	��cM�
�2I��{�a�E��	V7��mKQ���~$<]Ѥp+��-~�7<W�?|qr��f
i�\�!V2X�M�bL�ԙF�
�9
йJ�>_��u�:y���r��E�"���`�4u>�+���3�!+��,ac���!T88V..a�!ƽ��&��G��ւ�zs��ًp8L�Y�s<�F�
F� �p�-#~�TE;â��U��3�XL1 ��%��7M�>�Y�l�PR!Է+���ҏ��6���l�U�j)�	���v1E-:�pZU/���Ms���agM���������D�Ѱ�_rp�mG�����8O�Dg��G��1T*N��s�]z�ڽ3b�m�n�z�xi�?���*��:�,}�8��[����q���8�~=�;\�^+���Ů�¼�ɜ2��X���To�(K�)S|��$��p|��d6��kZ�UI������"H=�6���y���*��92���%�27N�er̜��1EI �v�E�.����@����Q���:�d}gp��6'D�A��_�ώ�\q���y�N>(��w��a����(H1t����&n�Ln�/l�"]#��k�$����2�^`�����Z3<	���|�@���H��x�(
��*х��N1dx�\���`���Xڥ=�C|�OT?Ԩ��������M�)s#�co���Ĺ6	��D`��>ˁt�A������d�/��f|�١�O�-�F��S����,f��]y[j�PR%1��_3��<����p�/���)�-aQCY7�L�NH�(�!�[���UpY�	5�E5^0H����B������m�9����� :¥N���o�{p�LW�(���$n�0}�x���<[�rӶqС�<K��ފe�,.mB�j�L��?��.�i_���|5_��cخ+@��S�H�ט+H���.�{��C���Q�q����>"Co��y
�&�_���g"�.T(o�� 
_4dQ��s�?������p2���o�>��}m�r�;��k��o�d�iZ��7�B>����)�:|ul�#bU)�e>6�c�����%k�R���Z�|�Zׁ�l̺7���)?1$�~ 旔��W�ew
�y֕���"�HI�;3�{.���`�($�^j-AT�FtT��F��'Ma��8j�:%�t����
�zT��k�q�ts�1S���4�8�j�N�voW%�P�:r�|��M:�J��d�w6���@��]�Q�� :H�$Ǝ'����Ihg��k��ג�`A'�|@�����%Cl�:[q�\�t��Ȗm*d��ɛ{��A'5�)��`@Z��j����橂�77�<�w~ A� ����k��Q�@4��p�6K�)�,ﺓ��7S�(�J�d,D@E]�l�|��"�i��ز��|� .���i)�(8nޖ;����խ's3�nKN�'��p������tM���u� Ch���SD�;���J�ɗ��4���I���w_��� ��7�+랚l9���PV����{��RN�����'dv%�$*��f�lŬV�}n�)��l��ov/9Gv�N�ЄS����v�u�m�$w{�p�!�f�q^��QHԮL4���gM��K��ă�ҏ�o2��D%�����0X�S��~��j6x�x�MZ�8WN��7C��D�>;J��'���(������w6�|�"�ҤS����=3�];�B�^�4]qm�{����<B�a:N\'�m^� y�TI����h6��_����ͱm�,�<)~��o��7A�I�@ ����f�@hͣc�d�Z�ܹ|��9!FSO���k�i�˩����F���v�b&b&mԽ��Iڸ�N,y�O\�p�p����?dt���,�`�r��6�ȞjW�7I����T<�k�)H�IW�<;����syyޞ�3�} ��c~����}�l`(�������h�0�VJ�!]���t�[j@�lO�+?b�5���oα޾g�A��r�L��kQݮ��Sr����X`^�Í�"�}�1ur���~�qa9�M���{��/��C���V�C��5��������i���(S19d����GǤ�y���i�]�	dQ�k+W��|�H\����������W@���WiE����9�n.�Q����^V�87���TV�(�뗴�<W`S�qwW<�
�	x�	}��y�}�Y�z~v��ONΜD����̓铺��V�X��u���~$�xb���6�]����=&K��N��nc��*� �(���!�N�M���!e�G^~p\K�ˠ��r��g^�V�Nߡ�HF޴��i�-JF0yB�ؓ���qH���4�3;/��k5��g#�æ l%���|���J�Ư<�� �^��\�:��y	|��M<ɳ�(�����G~r��[�u��B�E�Y�����7����|u%�����%��Ѳ�8�S	�[>%��G�iK�s�|r�i߁І~��yun>��	�2@��v�"t��բY�TZ$mrM�":�/7���27E�ǝʿ�"w	�,�g�����>�}*���)��<��#�����@{�r�maנT���w�Ȇ	����~��!y�(p�x�
�<)7%��ݷ)���ŷi'sF�x@��a��UfC�rV�2�=`���4n5�Z$[J���cq���7WQ�mrf�a�|5�	��'�夵�u��qr�, v|�j�.�Ty��|��;y/=$�T����=tn���3*J@v\�V-�wWW%]������ֿ���锈��3��-�y�kޖ�{U|�>�*�=�d\eS���t���x�ǽ�M��o��k,qɍ.�a[	��G�YFŵtݚ��<�w	�!X�.��\���6���ƽ�ƹ�������j՜�j�/��p�K��ˋ恇��4�$��S�~6��r�cCy��4�c��T��C����!��Z��9k�B���hӦ��j�/�P�o8sl��]���&��|��D����A�� +�T���ǂ�[�[:�O�J,����Rp�Rcu+�-l�*��l�iK�[�	��@]o�6��oN�Ku$h�h0a���b�0��=�WJ����Ȥ�c������E\����cF��������uz��N�Hܠ��KgQؐy�f��m��'��(%�����F�Qv#�sK��l^�b�n�Vխ�[�_G�;F�����|�P��&@���at�r���:3�[�P��39�����W%��+���&��2��f�t�(�[��np$����B�Û�x���l�G����)&5u��i岷��B�ڝ`n�T�q��:0smQ�H���M߀©`�5GTi���N?ڎ�;]q�9�����WC��lн<������+"�~Pc�v�'+�O׺��B�h���}��N}[%?2nK-F��&N�! V򜮃{��!�����J�;J��ͺ�M4'͔��-�R�x�񯭻#�,�)n�Ǆ���ESF562T� 1���U.�m�1�I��߇\B��$*z�	i�E-eD�q��hS�(Ӧ����8,�
髬'��+��Ω`�$�L�9��BZQ�}x��j�:��7���N�>6,����9���L4MNk��4Ư�4���|�f�v6�ͫMŐ{{K$�h���D���[�P�%W��l�0���+��{P]���p�:4� ���&jAVEFg.��$� 1��ĵ+��;4����+�����&��*����?�
�ξ�A
M��j����S pq�vxx� �a����zDȝX���߭������jgYA�XMPO������� QNx���6�V'�@1$w��t�
���^2�����6�*��5c�z,�5O���6I;�1�uٯF5�<�4���i�F�&�����r�sԀ�b..����T&��wq52�L0,Ԃ��������L_�3'M�f�|l��x3+�Eω�z�Ťy����?`���r��H�_An�9 � �ykaZ�D�x���[���M��K&�{��Yc�H,0�t������yh�lnD��R5�9�j����p��K���MJ5��(�x5����L�9��f,��s!F�KȢ�1|�`된}r�f��_��M]剡��x����j����pp*�WAQ�u��{lv���n�i='�Dg[n���F±�&�������G��IB��ot��`P�z�EXȃ�C�_2]�
bN�P*�6+z2X��@���(�$l���Lx��5D��fE��̼�QS�롰��dd�o���#+���z@n5�&&1gq�`r�ô�b4) ��-�Чk�+'�%O;�a$>J���;��VW`������9R�m6�?+�=�|��z}��_��T��:��iz7����?�)�z����n�EnB�<��}�d���Oy��N���ɂ�|W��5�pK3�R'z`X�G�g��/g|}w�j��؉��H��z�,�5�p�p�}��g�AS�]��^O �w<��ɑʡ�����I��*_[�����?h��[���������k��
�I5`� �O�`����0#f��`F�f���w��+|�.�y��{ޞ&7���T�ö��q[�[�y�~��N���iA�N�3per*���f)(z��vd��ߏ`@	~ߑ��ޠ�u�o�&������3V)�$ ���Х�+D=�/�g�&�
��mE���8���!�����x9c�?[�F�r���`��O����}����/u OQ?;j��]����`oȅ���f�����mK���r���D7e1cv��K���[U�������L�/�{y�X�
Jn�����{}����b%?���r����'	�q5W`��W���3����e��z,�ێ�&����O$�[�L�h0>�L$��@��s4�A�\�6Ic�^���BǼ @hG��%+�N�V$\�ֳ�"A^〻���Xbc���S�h�O���%<�H��Q�Qm��D]/��h�8�C?C�%�8���fN��)�6���S(k���\}Ӱ��KS%�N�6�|E��Q<'9����]�K�@���=�[����dJEc�(|����m�
o�&Iy`�2������p�����A mc!��F��X��6e>Ɠ
B���x��Fa��0MV<d�L��Y/��sC��jAi�1�n�U�Y鼜$��U4Z�n�2���%h|e*����y�~��72H��{�|��{���2�:��,_��_�p;�vB�;t7K��-���k��]�������(���@^�N�A��S�����+�4�k����%�:lm4Q4N��!���X�)���t�P2E���>,��-�|�G�ƌ�O�� [$#��T������7/[�꛳��3�������n���u��2(�'�w��ɫ���� $��t�r��Ců�QV��,"�E��r�!�jQNf`��3G`;<�El��S|�/u���|�*�ǸN�̽V,g�Qz�x^����Xv�
_���|-���qI�:�9���v0XYɩJ�R��k;r]L��?��kيf����޼*l����=3D�'�gX<�g0J2O��zIa����1m{��F�}�WW�����@�r'���n��v�Y���62-�3�aq�_�Ǐ�(��N��3����J8��e�pp��iV��:�R=<K��\�>����~0��H�rt۹����c�/F'd�Jqh��V�>�^6@n=��C!:�w�M�J���S_�2c�b�h��f�HĜ�j��L�����F`��l���|Ң��|�@��d�[�2n���SuT�Nb������� fhc��Xx5�["���0&�?q��A(�u<�w4�+�;��.P���o7:E��� <�;����\EJ�R)�@;]䉂7���]w�;l�A�V-̙Nw��k븝T�hǚ�ܾ���i6�vљ�����aWb��%��H�C%7�h�s�qE�\��ڪ��
��#~X���/�7�cun��Ac+ۀ�����≓�Ep�Fr+X>^-����%2dZ ����p�u�9E%>�L������ 3o��6���k�ÒQy��A1�'%߂�}
� �o���6���*A�Y�;�����!�%%����F�DS��6�qy\�N��Y�Ϲ�"�\w�����F�u�8�05O\�o���锝���8���A5\�� _o� �5R��r�*-������P^N���Tu>�����ϙYz��`�6$�(Q4(�~�Z�~��nC�p�:�=�n�k���ȸ��i��X!2��Tj�Gi���iky�W���YM�9F������8~gNO�P ~�3�������:���A������ӥ���/l��K�s�@����3t�
l��]԰���{�Z���5�\�FM������̥���Z���k-D��.���� ��J\~�D�aa'�m�/W>��B���������X����EwD���9aQF��`Lrޒ��]��0��¶o�*��B���4=w������d�s��+��9a�~�� ��{\\4yA�����^���k4
B�9V=���1�X����њy�]��{<Y��6����]�9��Ǽʡ�W����ҖJ�w7���f�,g��t��}�{?:�V��Ո���Ʊ��h~ªi�x���b����~f�qF�2Ei�}�����1�y��g�D��)o�	nRA����Χ���C���>��ۘ�jo��������͉~�:��$w����,vY)nҲWy7�j�e�j������1�yֿ`I�̿ ?Gx	���$�)V��O�BAH�`�������$}K�v������L���c))	;��C*�8w�hg��5i9:��*�����r��@����U��i��&�ۍ����m�&�7�?�"'#���sL���l�!�,�RҴ�[�6
ꛆ+ڂ[���+��!a�*檮�j��F�j���l��~eZ�9eE�
$�[_����/�U�������%ɬ{o3mC!Im�D��]�%�k=7���9�Z��k��˻���P���'#IE?��/L)W����g���yާ�����*)�+���}��"�zM��>��`�D��S[$s/�{�qp����Xé݂,>"v��Uּͥؤ�x �{:�i��Ak�DQ��D�fk����U/��m;��sH	F��i�ZF}�<I�5�h=/[�i��i��Z6|��#q:{g=��NDG;Y��^��� u������b�Z'Y��P9l?*�r!�V*'w���Ϗ�@�6�>&��'I�}�Ч6ģ�l��G�HE�띍W�r�-�lO�@��3�'�fI���tG1�'�n�N�")#�������>��#���8��ZI���9+)d��''���W`���]/�*P�i�0�~楘�Zv/���lݞ|��+����y

۸�
�M�?��.���}[ ���`���T~jh��j��y��f��4�mt5"|��|l#���Xv�Y�-��H�4��î���*�H�cJ>��K���Z>�OnyUYZs�����׵����YO��[�x��|/�I�n��8�X|�����\�)笞 �zgIN�&^��@���(������['�뻽�^=���>J��v��lA�����l�E���5��k��̯�D���=:|�7*PY���Ӣ �_L��Noΐ�a�LF,�l���v:�f�o5�C�E�i}3�G_DwWV=�}��〘��B9�ʏ8��P��~PiT$s(54|L�o���f��,�_F�BM��i�������p~���|0�����;\�����v1l������a�2�T�p]�"kq��jf���u�� _gp�"PvdA\�N�K��QZ�'������øy@�O�2�a�v�f#����K�必}:A������q=%��&�9v�?���;��>�Y#�K+��-#���C6$\~WW�9��ߌ�ȓ�����q'c�^J��BM�lG���N�����I�,�ID��)�ڦ�m�t:~l� \��\nT~[�Z{?�\��\_�r+}�Hj�ab7��W`�	���4{?�议�:.�[[�Y!�m-(��h��Q)��#�4��ax�Y���W�.P���'� ���z��|�QL��bSN��B8CT��l��X�Am�Ԛ�O������!���YD��Ù�O�D48^���qw$��e%�s5��R�&�+�8t �R��9�됖bS��(�������@�� �m$c���j���UY,h�?K�,��e��0ܔ�K��L��v�9����T�[�ǔ��{׽f�ẖ�|XI�!�q�� Gi�XM�=�[�<$oW����o�����$Z��	dB��}���A��z��CF7�(�w��o�4hP��h)o>�+��ڌ:����|���g|��3��[b�I�Ab��DO�z:�R!�w)�*�5�H<ݵ�N_얡i����v�f���Yjp�M��"����|a���2ʔ%b=W��q���}5^JeY��8��;!��ʅ^b�|�6G"�����-~=��|{����|��L8�j��v5�F���W�U2l�qʟ�5�=������qr�ȉ'ǆ��?})���mcSѵE�0�T�H>_��,R�wq������Zl)�g����SQ:^܄��$��ݱφV�=�4�IV~L�،�|	hr�v�F�a�L�q�ԓ)�׈��٬�-i��kK'�m�4�o�r�)��Oڳ���hz�����V T����P�+uyP�1���6��)䋣�X[U�o��`��;��y8uDbC̼��ob�[
�RU����,�_X�̊}:���4������||��y�k`�E1�r�P�k���qͪ���r�&�U=lR���m��E���O;����������������K��Sc��lm����|��LD���ȶ�O��N�C�*������Q��"j�xx����2��(��F+zF��Ӻ���G��.�)?�ݎ�O�h��5kLR���H3$���a[��"
K���y�K�4��W+4:���{���i����6}��
VU)= .�J�z|K\$��,JB�A�w�?��kXK�X7�B�M�%�N�|��ƴ�J���&�rc{��5��؂��|�	�L���*X#�w��1�.���6�����K{Gړ��j�>�2�����֕�=˗�~>P� �d)�(��Y�bU�����ٰ�n��؏(�
��`	��j�7�����gA�:�)M��[��@~*�V�s�M���1O��`]���H+M�
qyM20q�{�u����z�`���JDc�k�QF`����^�Wj�E0KE�h������Vߥ��W]�r���>(�')� ��jX<]_8S��(�ܖ����~��u���Ի�������������s�t�і!�u�QZJx�4Y7.��6�ƗeS�?{Y'��4�d���p�T�EC�*��jf�����z1�@ԙ��{v�yg��g���ފ%�`����J�&/��樲���ϴA��oOQ�mr�U�&�F����Y���Rn8ʘ��{��ma�6\��èj_C�b� �7����Rr2��c�����jź�PRS��tF��||p��2�W�J���N%x��Q�E�,�T&u�R;P�.�+%(ʼqA��%��7t��0��vmчY�]}~��c���S�.SϠK��W	�㊳rKJ�x�}����B�ʣxl��Z����{�T�Ȁ��c_�awg�Xa��j��Jȑ���f�f����!	(��^�6�R
�č����J�b�z�|��e���ʎ�����h֔S����?�#d�/�� �2"�d��uMU��6�����`���]pe���k�_��\�AL"��GG��,�w��C%L��ƫ1O��}�$�+U�����X�(�4;EOBd�X�*�6����ԗ�0�m�Ii���K��-�{*؇}�d�t�Y��E��(��[H]�r�.'�ᷜ���Z@�Foȃ��ha��F�s�����ǯ3��BDa���������ʡ���ܖZ��3?��)	3��CR�{��'>��=�7�m���iX�üm�(ptB>�[vB���;�s�`D{9��UT�k�瘈�`��~�P�T� 5���
=��n�U)8�}�S�q�|���B�hMs���H�'�m/�?Mg%��u?25��`��h�r_7(NS)P�;�F�滑"!F��J\Qb˶s"��t�=j�d�n%��*\X�<�U�G��֧�[�'�&�_�Z1kv	pC�=̂5��M��̬�R�>�s�F�9V��ã�����m���~z�rC{�@B|acvLCw�~�����}a�K�Z�]o��h��� �l�~ᵉJ�6�}����:�8�>7I��#K��_F��e���ܐ����y�U�H�]l�5Z�apA��U���l
��D^n>QjY�L�c7?��k�}p��du���
�v��S�S�4^�"Agt65����h�@M��K����)��<� 9�9op�m�W'^�$�ִ�]�R�,�Y��f63���$埊S�ݴ�9����a����]��x]=�:w�����`9y+g|��aG��B�D� Q�fcՈ鱞�ѥM͎�� �� ���z��8�iQW�&䟸>��b_D�)�ܻA���8U��Ü��l��p�G�����-=��Vb�}�3�*�xI�Mn��nzE֎hA����l�M�������:O��Ë:V�.fQw�i8"�s�t;~�nU�+���W�{���Crg��(�l��.�6L�2�`6t�G�{-�G�+Ğ�
���Rd�1�A�������*�[a	����@����=�E쓍���K�|�(��[_�w�pk|'$��`�{'�;Ճ���ړ�?��bpne��jY$��/��1Y��A�\i�(�.Λ���S
�;<M�)����y���4�y���o���o'�Pɵ�/�ʓog#��D��?{��c�����\��% 6�8`�ڐEv}�$A�ȫ��J���LH�>�QF���A"o�2-�˰)@d%��6W9��Ӿ8�7�x���Ul�q���-9�cc<�`H݌X�#�8_<_3N�׈�"��ji����=	f�b� �@I����㩬�L��{I�P�3��j֨��t���y[	�ʷ���	�7v�`Kv�Ǵ ,<�( E�Hܳ�L�'z꿢�Y��� `D�5����z�9}e$���6�㶤����@���]\��S��Ű��_Y�zJ�xB)����Aǯ��Hp*���}��	<��[�j	]��c�pF�yB�.�<���&�Eo� ��:�!�J9�mW��x����׋1J���}�3�Sa�ڸܻ�芚���w�#��߳£��8�j��]�ʉ�^K­k7ii`�Ѳ�Vu"��K��a,��m�Tn�RlOCmi�C�h8˹H�f,�6z�����}u�o��I��9�ԘL�K[lj����y��\��E����H.�Q��pH-�/<ݨ�� �
��I��r����$p���R鍰X~��;�,vCn�z�)9�S�Lv�q�%\��
W@�������#�5�j��iBa����se�k>}G��{��QѰI$���F�%��l���/��OQ��2;.���hr���R5��zaA�k�n�|Ĩ�L��C� �ZQa���9$)����Ry���-q��O�ގ1�<�������r�j-�u-=Em���t�c�%�KS�5e�J�ahJ bQ#�H�yA��|\3�]��`�^�O�@�<qkE�;����j��d,�>}���
i�ҼT�S'��kQ�� �J�E�\�i��R���O��>ސ2�Xl�� �ciڦ%�6��@�g�e�LK�.U�������֣Q����a��K����3j��}.��go��)�De�+M��#1�����9a�/���@o΋ׂ���V���A��W²���`�!��jW4cW��篶�����y��d�+A5D�#�jU�ޗ�mCȭ��R�G�G���܆��~�B�T#�������E�^c��hz�J�!^�mR��ܔ �[�WՑ #��A�F�@��|n~��.�{���媕@ISҟF݇ҝ�r��(�ۧ=ʗ�'�7y�eod0�ɾ��i7�ow�ڎ�	^T�{J�9�wq��V����:ry�"ϭE3���=d|�H{a382���5�����G��n#c	�|��t矃�T�%�v�$B�!)j�
{���_-�2~���q��!�D��n* v_�ӧ���{OC��5�L�t&��"�q5k's,ߣ���}k��nbq�!V��"�Y�tK�I���Nud/bNv���s��I8��J�g\�q���,�����O�}�ƒ�;>I�*d�cn��_n�Olv9������Xx�=;;����W�8i8&^4��=G��t(���H�~�9�p�{*��Z�ΰUH~�5�	7Q�jD=Pݥ俳Ć�*�� �Қ2"�!}�����rt�jW=�ٴ�?��=?7/�������t[|��H2�ׁ�\f�9�IQ��XhD�P���BѪM��1Ϣ`�*^؂s�O����2~sY�E��y=���Uϖ�����织�Oي��aQ4e)��D�ɇ��g*��妽C?o�(8~�J�� x�N�M�-�e�7]�9�����5��Wˬ$?)��}��-C_�4��$�b�ȳ6Z�VT!�$7��j��<�'7 M�EP%-CD<#��F�搩�b.�&������R\�CEnu����3�܈L@.[�8텠p};���t�G�o��(�e�E�?���/1j���Km��=��w��X��M[ݳ�eJƇ󵓄��9��ߏ��v����F^��<���������=kh�XK�'�\7OWPT��w�=�	��Y��LZN�,C[�K�Fc&�:C�f:7�N�g��F?&8�m$�x\y``9��Cҁ�M��-~�����������PnU����@���~J��L�@��l��	��l]Ը���[j܊�x�F�HKi�ߊ��C<�:�l�����ok�}��/�z�i,�M/�Ґ� !ֵ<���Z2ա�O�B�DX��3x¢}s\��T�l��o�j�Y䥉�YϧL�Yj�b�L�?�JuVn��s{��y;�<�ː��&��^�T�?pjR�& �Va"J	+���r��U�nZ���
G�톃O�d��Trv1�3�%VU�JZۆ�(6<GE�~HPuS>�Rn7E���c�Ӆ�3̳f�.�	m��F*�nе}�5�Y�6�*dK7+$��z��/���n�+'�y�O~���/e
��Ϲ�ӿp���4�ӻ�Jn����H߃%��t��&�K,�h0��q�Z�"}��������>��#|M�܁�u4114Z(v=���ɒr[���>6t�zb7W@.�r���SY��x���׿4��[�l�������4�o�o@�4��Y�����tH����[Z<0N1�7�jD�`�����'��52;���ѩZq�]�:Ga�vxY�΂�tVl���0�q�S�Y�ο�Ww�����⳶�E�����8��f����Χ��qG��^i����xN)⿻/�V��W�9O�����������/n�ױ�oZ����E���������^�|�?�|�j��-u�=��v�ר/'
����/=7`�Z9�)�-��ܻ
�q�Qw$�?`��{U����"_����lҷEv׫\0:�@���j2��:)����8^f���	�¨�ޒ'���^�\l�D2��
���@F:'Ix��?�nd*��>���I�zHH�o�Ҿ��Փ��/ngT����'#,�7��bq;���
Ue�<y��{��MZ��\��l�ww��A#}U2ٽ��H��éP�?Ij�GQ20�%�Z�:]4�/����V��(ry�#���N(N��G����
��Db?5�/R��[o{����;�\{KB��}*����b�/d����� ��N;�����S%A���b�����^�L���Nh%��)�ì};y�u�H�iC� ��褹�5�L�}��uM̙���[Ȏi��Ӿ�"9PxdO1�β�,WH+�	'���a����"ȗ�u��O�������@���1iկ��C� Z��=�HV!^A"������e�����%R���5���)�&=�s��32qŭ�p�ܠ�G~"u��(�O,\�����*EgD�Ѿ<7�vcQ����&+�`�`ܡka0�ˁ)]K�!�-&�sg�?=��?K��^O|��)��*�(W�A�f>2�j���Z��|�c/���Qv��#�?ŉWC��*������ڏ�0����wͷ��d0!���-�����fZ�o��uS�rUw�1}���w�v��Y���i�'V�p��o��A�{W�GVԁ��Ӥb%߬��4H��D���b���RAx$u�s�8��H����,@�/{r���p�:EE8&U���:j��:X�3��!�G��V��i��u`�Bː��ӵz�p�k1Fζ�4L�K�� ʅe��oWKat�<��Ǵ���	 \�Z+���>{���p��������N͊`Ɵ$��p��պGgfU-���"JN'Շ��O�A�5��S26�Bs�y�z�9�B4&���_�OYv�D<{��d��=��l���i��.Cs�d'd�i	�~��|q	��/Y,Bq���6��d��sbل���'�q9���:�)5h��$^�����(����S��Ԟ��`ֿ����w����%��>
o����$��k�����K2N�_�����2,D�}�k��1ܥg'���r23U,����0�"���͎�+W1�'A��}mY�D�d;n�ߢ[h��'�B���q����8���{!Q�
�>�ս%n ��Ϙ�*9[�޻X�,��G
Q��,&�~l�E2���)nL�D���B���+���νK]Pv贈lGW��Q��O��y��[�W��r�$��p��[�H��X��b��<��=1���ЎM}�pmPi�>��T5�w@��})�<ڭ4���N�g�*1!Y0&U�G`0/�:U��KG��]'��J�2���Y��G�����گ�Wr��vz�Ƅ
�lzN������&��.���ʊj5�B^(��ET�!E�h�����M8��*�Ҵ�<[��S _���י����no���F]η��?�������-��j�f�k���e_���lK[���Ɵ���O�k� nN�}�����o;��mش�[���`���i���}�.���.MD��qY�X��/B;A	�	��}B���@Wnٚ���V�WD���l�{�;��%X��p��8iϓ�����pM��Oh�}R�d�Z9)��[�5�{=jX%HC�x��N¦m�|��=R���aKM�Z�D;�M�����'�hΙ�2�k�7��Eg����~�	�Ay��2s�e�N$������Y����r9�X]�zX��|c�a �8{oW���Ǟ�j
�oGchJ���,_������p�3Y���?��߮�g*ُ�j�O��(>�վ�>zy#�B��g�E����R,|����9�8�i�̲~���h<W����ȥҞ�Չ���/go"��憗T����ߍB�w�Zt�O������[ZN�~�a�o�" a&{���Tp��d�
40��]�c�l��eO���}(�yD (��fGH���=hg�~�ű���{(k҃ S>��S0����"8 O��ms-��S�[����f߉�麼��Pb����6Kv�[�E��� )w��Z���7��2){�m��ց���`�9i�+K+�5e�V�D����{'7wz^���3桿�k��J�8a%�w9�M|(0��e������0���Tz0%<ʗ�_a*.}5�"��(�QͲ_Bo?�Ь�=wפq�?X~�j��Tn�F�Ԍ��n]�#$C��ߨD[��vl� z�s�J�+��fD}�	�AdYPs��|X�NI��Tk��G�I�i��w��w�E5��j��?{�$A����YɅb(7�e��Q/,,Hh�=.}%��3�g�����d�iM�Z��H�ã�P�18!�0��V���n�b��e��	�Q�X�c��/�ȇ��գ<�!}?r��
�"��S�O-�d�8\1��i�U��'��h�j�Y���S�N�N��V؁�&�"J�w�ЊLzO��[�;�5F�	�'߂0�̦�{ U��q��.S�=�J	Dʍ�k�����Z��gbP����ۈL��0�O9Yj��]�Z���L�+=9yr`980PY����4�&��i�5ƭ�3f@Z������˚/s�bl*N����%�[�">B�S�.S��鬃ò��!ΐ��ټ�)^��X�V�P��!7����@���y��3NϞ��f=���v�-7���&��=l;'��BH�.
�4b�Y����Ph�����jH��QȔ�9�����0g�8T|����A	b���ަ�/7]�:���t�3�]����ގ��,�c !%�6(�������5:ի�e@�l�q�@��F��St�ڔ
n`5��	��u��'P�fJʁ11�3�� �S�;s�w:���I��P?z��*�1����z�{�#U�+7Wa*��=%�R=7����3e��M�8Q^��~�C������jCԭT�mo���^������,��@zbS�X���d��)�A�=����=�9-`1&4�k�h���E��L�7 Z�˞U�x��
[��94ѩ���Oc�����MUk�Th�6�C7c5��j���9��M��d���0%z������}{0á�����Z��,xg$CǱ+
��-�����k�|ܧ�=�k4�"h-~�F_χ>��x��Ϸg�˧����!�e����`�<�"a�6��a���ʒ�ϳ|�@�:
>h��]�X뵙��h�W�!�T��{_����>�U��Ьu��(s�r��e{���6����.d������s���M�#s1��Sa��^�Obة�AxtS*��j��vJ��dM�>�9B���Y��e�6�Y귈0��"g}�9��P�����ױk^����2�g��P�Zb%�K���87A�K�7[',hY��_ b����f���}aǖ֩��X�=�ݔ�bY���8��	�zLҫh+t6y��A����O�UqZH�_OK��>��unY�dMb'����o�NU���-d���ضf9���N7�'�du�A��Q���A~��u�q�d�2��ʷ��K:��FW��F��.�wQ�Kf�)�sE�_h
�#�0�/���d��������a�츏A����S���TP����p'z���(���ט�P����jr �82'�}VQ�G��$�7�մe�N2��U5��ֶ��a~Л���&���$s���t��Q�17�f>Si�HYy�=�V�GR�>�A뉚��@�ۍڿ.���h�J����J�v���pXf����$?%���"x��c�xS�d ��e¶����Q���n�0 ��ظnv�����߄���%��]E4M>0�����e������+�v����{�}�����҈���A�����n�sȝ�Ռփ����UI��*wH{��3���Q�n��Ϋ�ʡ�����n��"~�v�w��L��p��� :�
���V���I�҆�`ʩ���zW1֐�F>�U�0�t�OIZ]#���7�f����1׃"�K��Os�|l�n.���[��!�,hϬ[���sW]L_��A�؛��0�yT,ݵ��p� M�' ���mI�`x<�)�z���J�H@�E��H�'�w�9�ߡ!^T����T��|M�9ŷ�(9�J���g�
POL�bA�n��W��g'����#�S��^����B�53`1��IQ���׻L��/��j�l�V���8<��[X�\׍����F���U)�m�o،�:���k�]�r��|��<�f�!G�}�x8�j��(z���n�Ι�A�5��\��ןGL�S�@��Y��!�)Bi5�_�=�־�v�����d�Im�L�a����p�Di��+��'��T@�:j�]��[D��;-�p�m*�7����@(.u���B��3�#��5v�ޅ=��1����@�_83��'�]itS�7^ͻ�[έc#�2�.]��j �k�O,���HS�����k�G�_�'&m?��X%R�����M�ܚ���8�2;��ы��6Uu�}�o���()����ϯڗ�F�o(�)��`WWA���M��Lr-cΦ��������u��'�5�`(Y3cܰ���%������ͺ%Ҵ�T?��T�`�ɜȲ�v#
��5��U��ܱ���n{�.�Z�3}a��� �N�����b��
|@U���c�] <u���<� ����������D9�*��(6V�6�?v��SD���e�v�F��Qw}��J\0��@�>z��@5��u�kvjr�C�2��B��#w\��Z!�o��'����}k�D��<d%;�W%�N"S�ӡ ��������b×���C�"z��)����J.�5�nDr��ܾU��/�������/�� m·�v�N<�NgThW�v00C3��9����~%����o(1݌ Z��/��K6�����5O_��#@\*ò�l9�Ӎ�qK2��4-�`a�d%Ҟ`�� �F.��8 6I�Z�(��,�H�v9���T�\�x�sa�&��蒸waǁ�к�4�]�ǌ.�?k��y��Z�PB�]x2��n���;v�Wz9/�Q�>�j�'�w9	�w�Y(��l��s�i7��-^���HE��/��L�x���%�����&c�صC1Z�3[�B���B.�G��]P������$�m�r�xo4+��r5q�(�s]�Y��Hh䶁���VTgMӡG�3&-D��R�[t�ʵΉ"��ZS��vWhG�ܖo����(�~&�q܀E�o��	i9�1��Zv��O��pR�7�i���H�Z=*�k}B4�n:]��+��$\	�ǡb[>��'&�/*[s�\�9�������?_�;:�	`9���)�*�UNz�-�'���!J_)~�i_9>��K��}ΙE".:&��w���	�v�/�J���������v	�yo�"'�#h���d���j��Om%�n���xsɽ)VC��"׽�Q��݄�ܗ�������;v�[�`ƶ�t���VP% ��3[�|0�I�5<�^�eR���Ӟ�,b��d�L��mK�\U9FO5��Y/�a_!���ћ�� B&�l��H��L�YOgۖ)�_���^	��k>���)`hn�)��3�ScBd	���YP�RZ�T�f�{sP�f�ȼ�YoQ�T�.Qbx5���b5ޜ�r~"�r���qQƐl�Q�+_R�Vȡ�i����u�QQuki�����������Vi)�[B�c�@��������g-�8s����a3��Sp�׳6����(���f�٘�Mg�� ���9��2ʴ�kj,�����Ii��!�s�3=��-��fGYDᑈ�����TG4b��:��?D�l�d�����o�I4zJz��]X�J���Sh���lX��~1�2E���	����//
`�i��\�6�~�^�5�倾��ւt������%)��]�~��p�����a�I:�a����#���ޓ������q����J�U���2��^����s�׿[R�L�	�����ӯ��:�~ZWM|��-�zx�<����C�J�ڣ�?���D\��>�z�kl�S�J4|j��1C����i���@�ݽ�~��2��g�Bq�4"1�� Ϥ6·I�DH�Ԍ]���1! �yed�0�C9�1ů}��1E@Ԓ4�3�I�Qh*	Q6w�T1ʚCZ3���u���YglY��t>^�#�@Զ@\i�qlA�=�	>�$O'�Ԃ4�֣L%	�Ö�$+�9`�\��Qͤ[�<W�;�5cJyrC�Q���0y�F�]A�j�I�^��Ϸ��=�d����O�EM�"\ͫ��øA<��u�Ԓ��+�~�A�n@����~��)'�M��o#�UU�70��6Ԧ��ʐ�Ls�X�r0ݣ�A�.����w��R�D߿6uXv[d߅p���^s�e��S���[0���� �ʺ�ox�ä[����o5��NdJ7���X6�*�.B>"ݿ���w'�'f��W�L>�:C�W�_".�����C�Q�N�4$��;���.T6 �/�����'���ϡ���ۦQnXb0�?V�3/��4� Jc]���;̔�m(�;��-2R��-�I͐�ؒd�ϓ5J����j��{�c<5��(_�rK:ٞPpﻝ��oG�Y�I�uF�,���.[�A'�Eއ��s?t���D����([nC�������k�{�A��A��n���
n�C5����Su�ճ���8��h��)!�(�Uۇ~�]ɛa<�90�+�6�>���kĉt�����TT��A����:�%�����+n�
g��7iW�*����e�Z��deJ�F_��@��Ɇ�@X�q�s]��S�̔�ӏ~O�l�$EA���FF�72��oJΏP����`��\ V�k����a���~{�؎���h�]E߳fN�Nd,�>����k5��2�Tp����-�����'��,���A�P�B0	�0n���U�SC>�|ͦ'H�����;����-��z?pV�x�%���),qur���A|d��M(���e���a��E-%�Qq�oJ������}��o��`:�&3B��z�T�h�'r�?����I���OS����m a�K��}���q�} h�,i�$y��p�jh�TT��&�sL������+O)f���R�#v��sմQPu�4l���o))A��m�DU�>H�#�\�j��2��s;i�t
��s�ݴt�J��h56���N�!�x���l=e�;`쬥P*�ik�=b�a�QG� ^��� �0���v" ��J��xɱ��{!.�^:aݫ!�mn��UDvi�S~eA�7�:�hYK-�c>T��5��5U�ިx�=�e�L�D.l��?�����.<��͛����^(�a�ތm����R{�����EP�F��**bFďE����qi��7��(��Y}�B�gh�~7�#�C�Q�Z������� ��f�㗶�o��QR�A�����̆]0Σ?����"\Db$������g�;=����0�ժI�>5"���g��'��n��oo��\�]�A⽍�j[p��p��Sm��*=E��Z"%���}�mS�X>S�0��9�Q���cr��_!��1i��p�]��k|ʇGD�Zx��Q�#��2��2$��@ſ�k��_3h�嶴-ymO_>((e?i-x�_=pBZ��ي�4����lFp�@�l�0�Qi���{��z$��ED[ ơ� �`58�L966Nh	A)3�YOY4iϲ�o�>|y|&ֽ_���#
д�*f�Ra�;���-��w��ƭ�﷥��Ur��BG7^�wf4������'��	�2Dm��N��t	�6��3j�	w%�u7t����A���5��+�c�]��[��p0�zSy���wg1�+��%�66��:�D��%����{�^M���8� �T��I�7[p6Q��g��a��jKA(E¼x�ar��w��i��j��હ�n-�J-ޏ4s�%��3�$0�y��#S���_>�����@J�0z�$�bL|���)c,$�CI �ۺ�\ �����ŵ�G������ĳ�)��*��H�j	���~��وS�a�E�_��q�xCV�'ݔ�.t������74������1�VРJ����@����3��.L0Pf��Us��*����p���*���.���ْY{}�|$Չ�4�&p%�Ǜ(U�?�}¤��ɴې��a@96�3>�߰��E�8��L[p���ޑR]n�Z*��CW�Gwq_ӽ�޽\O�ƫwz��6��"�����F�ˀ^*�C����!������N:��H%Ѧ��vGd�C3-�JIj� �ˡ3�-�~�EHm%���F��Hs�4�P�_T6�(����ɱ�;Oi�������_��(��O�J�� yvj��&����j4O$��9��n�ãPO=<h����m�R�Z�W�7�"�Ւ��>+D�E��>ꄵ��;��ޚBl����砧�zTQ`���&:V�fi0���yzj�P���P���df?�{�i��Eݩ'��^� �C��}��;�)I�[ݔ����U���4��_��
�u�Q����������S9�B��R��w@�;k�	;RN�}b��HC�T�ʬ�P�t�}�O�z�8��j_cc�Vv��%���xk�0��A�Dp{�������7�F�CSA���B}�{���{�ڭ���;�ڭZ�X��Eu��G�k��g�Z�2x����V؏C��t�e�K����F�����І��%|��Ժ���a v\&���.��/����nb�}^t�$�̆����>Y��[�T�H�%wq¢'���3�k��d�i8�>��hFM��R�͂&/��l�R�'4��T��/P�[���T�����o������L�N����H8���G��գ
�d���y���.��@ogz�v���ڲW/�yWc�F]��:�a��I��"*�[5��bG��^	�h;������k�4	*%�Z�vL(C���Sԉq�(K�w�����5~�b����&���;���|~z_�M��s12�䬠N��J�ľY����^H�tn`�"gÂ�̃H�4\do���&����kod^�0�Y�C������Q~��^B�����X$�rw ���i� ��^�*H�M;��v��x�m�nn����O��ձ��
����{���w�-��B[���u�/j���H{Q�>���I<�v�#W^�A~�7@�����ኄxMв�Tsy2�������#:���`Oq��2�fB4��i�ߣ����f}n�2��f��ù�����I��%dm�ԋ�f��Tvx�� ˾�E�M��d���ʴwK�(�d�)��Y��Z�|ُ�Q�c��c�ԡ0ip����ט>�W�LZ�M�!�C��Y��`5-l�Z�k-B>n%�����F"�ö�Oܡ��t�����L`�򩒁�J]&�Y��<��	����ϊ���@-�Bd��8_>'Yn(=�0E+����m���'��9�ι�{�1b�6b��"U�Q�;�GYx�c��|�xW�G��9$ECObt���K{��b�q;k!	�w,��j�7���v��p����q�(ʲ�G��E[T���[�K�1�?!�-Қ��݈Xi�p��u��vg9v�(C�g�fq�l+/�41�c�O���JŖ�U�6!���Jy>��{	�_�]�T|%*^�z�B6]-�X�+ls��vȻ�X��O���5�.�-I���T��?�����J�t��(J%�;E��<;�/���l�y�qr��b!硫�$�,���j㴱���4o{;�*�B�wٺ�4��]��}�6�6��\���+i�Z
�k*6���g��L�Ȁd�~�f�z����n�"�(�lp��Pn3G��ޣ#v`�?�w>��Ԣ}]�Uj|����cJO*��{�J�C�~A�M��%s�s��C5�[<�A�	^�����o�\ގMw�cG��#>��t������� � ��*��÷�D�Y2�����ז��FAH&؞:�%�\���:�
R�&�o�~6H	V�������·��+�:;�=ϙ���2Iv�� .k��
y�h�B�Q��#���4swV�.*�m}����`�O�sA��G�ܼ�OEݺ`�7H���ɜK�h��ɨH����/x؃'��:�;Eu+����a��@e�r�I��p��{ݱj�A��{Q�K1���p�Z���.1x��6���f�0瑨
y�{�.���v��5
?5?�ɪ���#��򵛖��9��ϽR?)<}�v7�M�1<Զ��D>:�K���nV�q+w��>�\�α�*Ysx'55.�u���`�y�?���gW�n_6]g	"��v���;����	��]ѭ�������\�C���� �n|���.}璨�,ˇ7�<�����rҚ��̪_#3O�U�k�C���ɸ\�~��Ul���e�ZOP��v�a�P�g)�%����U��>gΗ}��{��%�7~˅v��i�2��ˮ��:|���J�,� �� �� �1�t�j��f/�҉s����y�g{����i$�w!���ֳ�p�%$/0'��';��6*�8 ��3��B�'�~.� <��{)Qpb9	�'$��ByQ�V�-����m&��1��t�&�
���=���-6��T^gK[Y��(c�Pw�u��s��l��Ώy�Y�>p
�Q�=��=0ƙ\�x���S: �Y������Y�(��l3<� W���W�I 7�І�tv4c����Q�����9�V��Xk�h����V7��F����⬧)�Z��w��W��ߚ��)vn�����݇p�L8�ui�Z�j�3�[,@6��o�,`�?-��v�҄uѫ�1�,���u�w;K�y�Z,d��i�-^�����v,���˚�0���4Ek��N!��f�>��56a���4�������Ɛj LU����d�G����ހ��1�T@F��dr9���?�uŔ��[s�m�����X�zr����7[C{�׈���IJ�1A�YmGߗ�+��0���BXq|�s�Q~�p�>1k�9��e�
��������9k2縉���sm9uNϋ�4���e���raR��)�GS�����y����A�`-F�%�tijf�� #'?:��타q[%�O������nt�-u���M�!s�f
�4��eݿՙ5��n/���b��j8R۹yQ�ډ�fj]�0����h7���|����ÍJd�9�0�;EUFi�PbYN�����a����̙O��6�`�=���A��_����:cT���#�A����t6���tj�����I�����g��L��5��d:�ٷ��d$������d��4�����%��ʕb%����E��M�W{2���;��.��W&G���X*�<X�Uk{��M~��CA�^s3�\d��B��$<��&��a���4�\�\�̦ Ȼ��`��",�ú�\t��Fx���`|��#I�uֆfi���`9�e�z�Ua�|�9_�s�2[ �8+�]K����|�~���-[�v:,v�<M<��#݊tʂ��^x���w\d��&��	4�k5�9�����6}m���u�8L��B��S-�g��EO�%�1�����L�Y��k�Q*m�O��
*|��v&�ōks]����G��nlqE���������y1;+qv�4_�+.w�AAj�!bǙ������U����:A�{1'��"JM0����G�������N=�����*�ZT��~��������jne�K��V��X����!�Bt�ȃ��.Z.d!Δ����mq�g�L��uA�i��kz����G@-⥹Ň�4Z��B-]���=�����;�¥���rL��M~��W�f��q:�����5�p�I[���m�>*k� _���f��.�m��N���kG�Z'�;�4�������8��c�ç?ȿ�դ0�NT������Wpm�0z�>�����/믿<P��Mt��
�<�:ADl��$|��/O�Ҝ-N��O��l�Vq�[��e�`�L�K�QÇ|Ɠɬ�}�V��O��ʄy�,��
�=��z���Ln�o�N}%2U�����Z �lؔD��mH��M��.�k�C9�����RKz��T*z�ST'S�q>�v��>u[ژ�(��q�et�,?���0ǭƧv^��$�nj�۹��r���^��
����C?���utc�kP�W?Y��BA-.�1��馤j~P�|e�s�l;�&+�K���.N>���,����Bn!L4�@3R�6n�5PjS�+��3e[�:�y%�}�!�y��\��w�פ�<�0��G�D�S��ǟR��ǐ��a�����
K]�� ����x�n�7E'�}�������u*3JG�	��ro3��2�]I��7.��}�'M�͞���s��
7Qz�V�E;�F�h����/��Vm� ��_�w���3^�u4�^5�߿�'\�AZ�OTE�*t,��JR���n�����?.y1��r��Wg��AJ�J��j�#X��6��M�鴐�?��XsP� ������0��|�PRӟ%3MT)���Yx<y�˟
�����9������Q��iP�RK���
�[����	m����7��1=�1�R�Y�[|7�L��p���/�֕������~_��c�������+�(i���O�
�Ud#';*d�!�Ze�fΠ&g�%�V瓿�[S��(͠tݮ=d����,���>�%�6�:�y2�M�-�ta�ߊ�(l��;A�V�ؤT�)ʝ�k���mSs���p~.͖G�&+�|"�E.�C̔ȍw�O9c��h���E�؏�(BJm��\~{͊2�<����|'w�xu�F)�C_�&̠�z=�:N�Ɍ���@"sWV�7n�������ȏ8P��F}�ڲ_�j�$����q�fC?�ƷI��}�(�ɻ��(��YY��x�%�b��6sIy����*Pfu� �2�1��H���� 0��L\X�:E���6�LoVn]c)|<����f9[�G���ʧ{v3J3�0�IWVV�vt�/We6�����mH�����b0���)��ZaiQ�Ty3t�F�	'��%%�vW��.�=�T�=oROzf������_w~�풅�5�<����H[-2��?/L�j���BAU'��B}WG��q�h�ܧ�6(;���|�����\xshߩt�s|T���iЇL9�׺�6g<��L^���[�h����:u��k�v��:��>��/����DN�<�G�(������n�<N����dO�q(&�F"�[��\m4���e��.��`�Lz�M�#�0����	�����ڏ�ìQvK'T�n+��Պ���}��§�9������2��f����]��Pr�W�Q�{I�3�N0�[()G�̫r7��u��Ց�6	�?�8ހJK��2�#t�y3pX�f	g�[Z��|�S��"�
(��$NL�41�.��3;�r1�ARlO�yr�����M�朻�������g�c	5L�ذ�9TM�-8f���M
�~0�<�q��\�sh��W���!Y̺{��dKϳKi��UD�У-.q$�Fq�J��獅��.a��R�!;[��Ե��ֺEA�I�ߡ.g���>�1Vr�YԶz�3n��e7��wq_[�A���W�����s��tx�ee����P]0QA������!_ ��� �mn��w�S�g[�ȠP��k�D^T��	fQ�0I!Or���L�3��#D���~������/v����O�H�������#�w��c����*�
�$k��͊6S7yE�t�d�#c�t>G�Rί��8��wb�>T;��-F��3p)�Q�7#x���/�i����h�H5?�j��>�Y����x�����}�d�<\/%�y.���W�2����BRYGo�����9���s��?��N�d�S�и�2	�T`������T�?�.���׫��VlT��W�O���u�Q"���K{�GO�g��  �[	/m����1���e��m}|/�	4ɋ�h���$f\�h:�-p&b���׃�M܉G1f�w[���cT�-��;�w=y��=0�ǍZ�q�#�J�K���>�9B�a=�L������Y�wRM��j�7�3��*�ڟ��)��K� ꌞ��gS�Q7��a�v�d,�ff�QO��k�r�o�T�	�}������� ���V�J��vn�A�V	9/4 u:�׆�t��{�3O�F��h�H�W6��/��9�:w�W�Ҋ���uw��C�O�t�,��볬h�/^��u�*C2el-2���`N���A��,ؠ�#;�&"����u�E�[�2��a��/(�S�X�^p�i�cw�	�3��K�
!����������LW��w�*K@Ǹ��|H�g:y�K�QسU�QѿW����a��e����,^��dM+"�w���!�1�w��WӒ�?�F����2~��v� �n؆5�������)M�C�m���S"MO���Z�����2�i���ǻ��@�������Ŷir�`���/l�����ZKc�!sl7���ˁ��S	n��ʧ]{��Gp��� ?$�e�<����:i��PvS� ���!5T��q�q[� L{�##��������湓!Z=M���Af�a�9�0[&�������і�����쿲,v�78��1��H|�K��|D�!�Av5�#�����Xù�Y�~ێ{�(.����|c�|�§�Oy��Ÿ��&j���`H�˗v�tw������(J���\� �@t�=hҕ�6���\��y��(Ke���D�w5V^t�=k֍�s ���m��o�����n3`�z�Ye��F�E��T9eG�87j����G��;��#�1�d��?��k�>��ҥ�Ω~p`���G�A����B�<�T�9Ĩ� 	���~�Z X��s��"�Nf^Ni.U7�q ᭧��!�lO^L[L�8���D���hsm&�]f��߸���ӯf<,\��	�?�k�����\�sw�
G����""���cGv��ϲ�.�;N�1��m;��7.AI��w��F��E� y�d�*MӺ��a�c���0�~4+�c�EA�����!O��x�Cǎc=���!��?̝�M>[l���ŞD����A��OA��c6ɮds�G)�h>Q$������ ��Wg�@L�EVx�)�2�̊ޭ�Bp3@���"������INg��?_]�a0���8?@�P�F���EeS4�ɋ��Y�����$���qC���_�;��A6��E"��xW�Z�~�{ʊ���(䪗<'8�GH�5��Wr��"!V��������)n������VN+c=�|�����^^��n8�z�����辎�
��iF�������66r�������5o��)w!�!)��n�%\O8��p�O��dďQ|�+���c$�H'�&H���=:�;Asuy1� |8��b�Z�q�_�O���L1��{F�.��]��=q Ѡ�cB�ߏE��v%�Ѝx��]"D��靵�7?G*��`EMO���*ݮ��6�6����#+�8��ea� ��l$D4"_����hj̉���ԫ����Ю��Mb���o��X|�ʒ��H#�˳��M~�-6�%fy	��aT��m�SSz����ĪI��|~��IEtP�u}�ovɍ��I�$l��G��(�d���Z蕇s��"D���vWg�Wl+{�1�=K؉��䈡��%4�h�ـ?5��xÄ��)j� 4��]��hIJw�����F���FH݁���N�������2��� �c��A2�l]�p�;C,~Q[�����]�H|[�(9?I��ʙ�E��l��e�(�[6j�e�J��NGv�R�1Ɂ���:��
��kB{[I���hP^#�&B�h&Y	�b�nJ1�rzfw��cߛ�n,�?��|b���,��9/v��%���To���h__��<�5u닡x��#p `��Vҕ���)h[�-�;�Kh��1Q��^$F�I�KYl��B}��OBX��.�=MX�+mP�Dw��m2^��m"X�	ڣ����2�<Lz����<�n���沛�r�	в�1`־�r�����\_�����
40&����,i� š	%T���*��ڃ�z�9�W��3�P����'�MZ�A��4��l��W𽞳�;j�^��l��$�BM� w�e��tAz`�U�w�h�ߵ|N�&򑎐B�E߹%��U��
�?��/��bIEV9��k�޶���Gw��f迮��e�3h>�U\�<�:�	x���$���O�Y����@|���!�3�䖵����ǖ����C�w�u��F�g ���uq�+��6&�%�H�V¹�F$�~��&�	���		6��b��w���Η}�@:>RZ���o��+�U]��<�YqH���Q��� 	�`hzG�\������H՚%KN賈�l E�)���.�c#��5,G*�k�n_g~hIr�@�@�@��,#�3�$u�C�M�i��R-D�t�:xR�}�7��*�&�R�5�a����h���0�����i�<��8[���3��-�jkڳa�N8Z���+q}m�b���A��]~�h >|�6<��4����>D4�%���K,�9�z�ex�a�G�H EE1����o�ZŎ%��zs���	�k���ˉͫ#�_��HAW��'�2����~��@��P��~b7w��v�O�F���t0F5t�kn���IZ�'2�NO1m���.�ͫ���ȥ�u�mp`k����n�w���?��)��~ޒ�{��1���ĕ*
C�>ʒs�����������Z�Ͻ�x���츠 :�/)��<��6f#k���a'>չ���a�9��r��'�����}k�w�b&--<����7���G�U�|�\�`5�*��M��b��d{�󰟽;G!E���<��n��:'�^���I,Fpjl�%��₳�m7��;�X�3��P��W���`v��m���Kk��qG���[+�tb�k�D�3��U��v�LU����F�l����������	���t�U<�{rV�@�� �aB[𥳜,S���~PҲB��ˍ�i��hO0��3?8)A笿"�+b<`P�ڣ-/i@�©��k��h���ڰju���&�)W���q��	���x���8�eB_ɍ1���݆/w?>���;����DU��?�g}DK����݉<�d>0��ǎ�3�5f>�9�ܪ�/U����L��D�M
�̴�7��_JH��m�Kt�C�;�{4�=i�=c�H]�~��L�$O)! ڒ������F�6~-�'Fk�Ќ��3m�D���z�#��f�۵c�i�%��N*-�6�Ox7#(z��N%�&*��Y�Z����8���λ \���Nw�T�l{��LJ~^�����4���UXL���A+�l6�<?�Fȑ����=��bm@uף��QZ�qx�<�@P.�Eq�k�?��Y�lU7dT0���4���E�����O=fG-��n�ћ��P+�y�����7������� >��榇�
�O���ݍM�n�#�A�g����џ�,e���o��M��=2��aZ��Z�P��j���3�������F�\�C瘾�|*'lo�8�گ]��(����9��/Ո-,�z:5�F�5��2u3ա�V�q_r�v�����/C�3��u&�=�Z���Y�����%Г~3�$|������I���6����������xa�ۓ��1�z�.�7��<���B�/�c)�o�� 6��w�{����4��o=0���k���&����CXd�0�-�=���u���\�D^pL�5s��-Q�C���lF�wS�l*"8ᴅƘ}�O0�� �1d?�y�����o��Y5R5�E��g���]��R*���M4���R��Z��(jZXuʣA�4��Uń�L���Ѱ9\�%x}�7�t[��f�������B�fdu8�7|�h�*�C�g��C�u1��
�4f��4/w����ˊo�CF�v�a�!�f&N�Sw�<8�G���$�}Q�џ|�����^�����������_m/���bX�-ʑ&O��3�G�sŠ�z��C�K(ɚ}m4�ǅF��k(�j~M"U���� *^`]!�cY�!���7�2!q�E1� �}I@ŖUxhOn^D-�߽8���\"�Q�l�tȱS�B���\\C$�i�C*�ˋ�)����)���O�����\�|��9;7�T�A��Ix���㎝�w0w�,��@��a�~����2��[$��,@��1"M�i|��N����Y����պ�Ė�7|&�A�B!�:��bVВ�&w���@o���<�4�)�D��b@6�g�e����>��&��/��Z�6b�;!T܈��=m���LF[���֓�e-�z�d���/:C{wj�z�'e���6l�c��&ȃߺ��.�]��[0��	�b�险v�=OLt!VX¿=
*�Y�ae�&6o�f}E��܀z5��QD÷�"t�(-��Sd��GS��Q��M�9����NB����uv�,a:�FiJ��f�c�ۼ䦌b��Bz,eG0��d�H�>PA�
���(Z&�ZH}evkw9D',�O��9������;s�.����>g�Q4k�pee%\%���2˸�!A{g@�S_ˍl�S�TY��r.���	��t�
K���~}q����c�M�����N�r���Fx�n%�������1ʁ�(Jֵe�l/��M���1|�u�^B.5�}��O��p8���q�N{������;]J
䛺	��$ 2B�ʡ��b�;'�&�+A��؂��C�����L�7�z�r�hn�ӗ=�6����Yrr��0ajC���}�+����<�"�Ӄ�?us5ټ��c$z[�}5�E�5>��?Rѭ��ڪ�kɡAt�?WB�j�z����n�ŧy���V*á�.��9W�����,~F�R�ؾ7�J�?��VQ�������6F�rL{#��K��������a[�ī�!A�F� //]�����Ɵ��T�0=�?23�x�����������T�(N��#����o3֓&�"�ZntM��s��OBY�Q���3}��x	�v�$�05��!�uNh��"0[<O��N]�fc���~x�'f'Bb�����S��O�]r��G�?N�}�-���+���$G+5�0��x'�����X}g��ٽ��h`���nG��a�Ri���)7
��Y��n����� /�k���C�aP�XE��y��l]����Lk�&̘6�1���]�۲}/��驌�fyr���'�PL��sWQg���]�"z^��g�D�%λ�Q�#�w�VK��~�]��h��%U���`���<��X�ޙ[���fJ�9�z6 2�I���a�Ziq�W�6*6 ���l��g�Ű9iM�4���AƢf����G�&�������>�}Z%Y��S�~�X(; �Ji�ѤH}�/R,�!�6^O��NAvNw�Me(���J���b��maKB���	��EC"���)��ʐ���5/������J`��Z@;P]��#s�87d��0H�@�0$ 
"m ����"��}v�A��m2�n�FѨ2_/5���w��]%iͽ���:�8Q�����3>�K\1(��������#�����KkR�VL��|xC��MG�Ĉ<����	�ew[���1��V�Yi�t'n�jɷ�}��$��e�b�q�W>�A	ʉt�<�r��}"��d�z��?��x¶X₶{Cn�
Q�uO;$Gჸ ���AZp�r�mU��p���K �!����h{�	n�&����fA�Ak�7��lspw�~���)&;�>5��=��������]N&ߒL�5��iI���]����+39��N�����(xp<$r����],_^Ř���3i�>���&�q���Z�t,fsC�Z�Yj["��>Q���t��W��>7i�P��Fr��ի�R�,�5��śx�,�8�eC?�G�If�0���c���a6ƣ�π��^6p���)y��u�`����f;�Y�j��'0��'���t"6�jG 96ې�d9��k��kd�Eqs3�j������5�'_�v�Y0O-n��68ݭo����>�tl���oʵ�z؞���2�&�m�&/���O�rP�⼵����'�r"�p�BΓ[0#�o����jf�b�r���e�)$$���7�H���d���1P@ �zf���icǿ!�|kz}k u�����(�*] ���a��T��9�k��=�~���c�J�LG�#$R�����Q��ԏ]T0�fF�h.2ޒ����?��P�b�nUJ���ɯR��	c=�M�����R�YF�o�ٖ:&�!�E>N�a~�;��P��{x�@
Q���R��O�E�CK��{2���-�ǡ��ab"!R�2Bʲpz�d�$\�'��-�m=�s|$e���"mm�A ��Fi�ъ9Ш0��'�v�����:h�%)��#|�T�7!����=�A�kT�Zd�U�;��7�Q���,���Փ!迄з��;�ڏ�N��VAX.���j0W��,fY�8��-~?ĬŢjPh&e�rwol$�j_���B-	�������%5�Z?�J������m�B��>���,�q+�p�(8��kҭ�#X�b)�f(�%c*0�Jf�Slnv*��\y�����2,Q�Xdi��0f�� X��-W�9�i#A�/�(bUր��.�.l���;�+�ZWg>���9v�G�'�x�����\x�i�����Y+c�V��9���8�P��0���.�&(%��5��&���-���od����^N�X�0�$�0*���m>U-���a���k��ܸ��ű�9�m��p�L*U,�nw����*H��F%A&��HB�7�!�Oz'B3��81ʝ���7,�mv���d�n}�9�H(sR.|VN*�7�[ �}�g�a��0����nc@)�f�����-|M/�!�jqz*�������;���#d�`z��K��� �ƿŗ�x3#���q= ��ߕ���|��7G܁����V`:@;��_���L[V�@����
�T���T�C�ϙm<�����O���vk����	�x��:b�+\�.	�t1��;�S��ʚ�'�~#h4�� ��[;���x_(��k�bT5�WrIT�=��1�@����B�k���F�h�(��*2}MԐ�]=�|S3&w;խmr��TE��l�C��k+�����s��N�<�����+ �9\�.t&���cgQ�6��XQ�`,Y����s�݃�f���$���`3�U�Ɂ�źS�ke����_t��7��]�d���0p���RֈmUWl%��/CO�6��ܠCy�QE��R��	O�#ԖC
$��C����fQ�g��&�� ��]��Z�C$�*I�� xp(ڴ$��q����ߗ��k��z�?˸�S���6W��U�����9p���N+_��),���ܥ�#�_X�m������Eu���Ko���V�=�n� �_�!�w(Ʀ ��i���+�˛�He�E�^n#��dz��Ŭ�9�����$V<�r��H[�,n��c�΁0o~r(õ]. �ؼ3���=�E�8�M;&�%��g/c�5o��k��7I�u�)��?ݛ�FSLMV��]���������Yf���ش��N8�d0�4t<�!�ɀ����{�?��*ڵ�qP����{L�Bl�7��4:��s0l#:��%_�>�]�CT����|�����{;�V�АG�g�,~!$vv��GRݬ?���V[�]}�u\�ЧTX���^8����`U�.�M'�F�~�$��G�>�=��zȵ��d�y!�}��n���C&����?z�S���#�F��^Y�DA�ܕL3&��[�f���'�`?�?�b{uN&V�1?6�}��`�}y~�]&�l"����Gf�2�b��T��۵�K��By9Y��+V��0lh�}�ܘ�H{v�b����������-����ނ���p�	�'����(��?>�yӁ�����'Oɮ��9���+�/�噢�>T$W!��ɜ�Go_��b?R������"rH�Ub��!�P��kX�q�\� ����Q��F
�\�Vy�}�x1��8k�U9�r����[5F�� ���R,�ˊO
�����[V�<֩����̮�n�x�`6H;�4��?��x�q|���������@!�����5H���!�w��w��=Xp�<�m>�����}����Xk��OU��>U5�k�k��߄�tb/���rKȵu�Vh,u�3H���U� ���FR�*\_�>�Ē����P��L���u�̪Z���ȄH�>�q'�`��M���H����Kh��t���T�M�W��cx�K
�Inw}���u�(\�J���t���@�r�"��nɣ��z�!願z��a[����"����Bf^���ċO�7���L�QZZ�����j���^�_�N�����<r�к�̋��ʼ�7���T&��}?��k�Ճ�K5�ʷn�=px�ѲY$���f�����w��	�&��ֻ�1>Qdܾj�I��u��`�'�7�H���Mܑ��c�[ú��6_/�.�_[��-��P+u���Z�O���Hu�a�x��i?�i֝��b����L���Kb�>��\�D7�i����W&�87���rd�]�c\�nl�F�p����5���ʼ�
��,6���Y�,~kc1ڭ��P���V(2_g�Pl�L1� �Ch�":�����sv��Y��Q���z0��^�_�������"�i�(ds>s��s�/�ֲ���nP��[��;�,{^wˣ�_C ̀�y�c��e��N9B�vx:��/��P0A|#I�v���R���ˉ*�4&��e�ݨ4GZ� zk}���������j��G�}̑�&����*��`���T_g��s�P�}i�	T���O��FL,�����9R���/|!~��5!�V.��]:��׎Y�P?B���M��CC��4�Y��ӷ�����:@0�̹����]�+Za�f���/�'.��1T�y�v1���J��{���&4� ЂZ�iږC�A���]Ǎh�m���F� ���DY�ۚ
�#��o�!^+�NݫT���-��}xQ�P�ӌ�42M����]Q���H� �p������9�|tmO?�K�v��QH��3Z^L<��Ǧ���&u\3u��p�թ���D�!͉�/��s�?sK���JWC7w���?��P�6� �H��y7�á�"������<P[��ˊ�o1��oa�#��I*Jn�V��٦�L$@^����:@�\��U�I�k� ����wJ�B=�]�3���r��#�{���b���[���=���1=gE���� L�*%���`8��2\��!è̏u��pE�dǌ)}�ឲnQd\H�� �[�k����w�J�4�,�{a�ܯ~r?�+�S
�yn�<�s[!�>����\�7N9�m�>Pw�{�r,v��d�"*ʺ��G��
$0ɳ�l���z0q=���!��XE����,\#@pjb�wߨv$��)ʜ��{�Rԯs&�3Ms"�2����5럟C>��N(�J�v�/xi
���K%N
$���NZ$�5��|o �@�T�(}��ڃK�'�L��3�G�C%a۳޴�ע� k����淎��ȸ�=���Ũ?W�'����**`�2���[w�]��8�pMwcBx�t\�w�~��f�F��7��e�����G����Z����:�ⶂɿ��J����,;�����8�'<�� ����7w�u}w��=�SH�����dv�_T�i�2V��wf���ӻ �i�_yżAh�h��R��B� �8	����lu���ְ�[�k�`Аw#='WG]+���ZJg�G�}��*��-�X:a��W���H1z_�3Ss�����"w�T\��}Bv�j�Gigl}�Q���V�q�����pst��!�6%E�u[���,ǿ�pE{iR�2U5���m��zzO-�� �<����n	����ܖ׫>uVu��8��r�$jy�xXD*��d�L��Df���\��vu<b�ٶ�ݡL�1�f��ͥ��7@�).����c9�p���U!��(�e���Ǿ���.�o���T�-��ɑz=T���橌櫌��VI�T���O"'���5��/d���WRx��.:/�^�x��4�F�WN����فj�i4��;��{��CJ����޾��}����O*O���p�3�Mk�M�)�S�9_�~�5��𜔝����F�ipI��h�/9;�V}�$�?c�(Ӹ����^���U�o{��.�#��2ZΧ�VP
I�)�u��q���>�_���1�pl���.
f��W`z���d]����I�I�Li��D�>��y����'�3^�n r*}��q_J�F+�U�|>�?v~��^���A�_M��p�-����u�N+�=PpKZ��N�e^<�ƣWΰ
���0�@4Ko�p>��˵xxr��)�es��^B7�E��-��
ę��ʶB?C�0�0��s kڗ��P2e!�ó���N�7h�ۋ&lJ\Z�7A�a�zф�L�_
�Ma��qkM�p�!H�\�HW���7B�Z��A�(9E��XN=���	����������W�l�V����	��󬺺�D���:�����5M/���D9ѝ�$#��N�&Xq���~��9¥e9\۝X�-
���ߝ�j�$�Q@dpx;��Z;��������ِ.`{�f��e�	����Jlp#�t�q�2cH���f�wv�B��������X��:���F��{�e�v��#o�Vx�=泟�M�;$�\Y<9�,R��dz�Y��c�[KU�S-P����H�;�b&�;@ �_p�K'(@�V�X��4�9��m����ȱp�;??��:���nug����>�>z�����~���y^�[oaet7-Эt���f|q̻8��N�	����_���+�=e��2�ͬк�Ѻ�}��n[��1�#���.�8���&>�����^>i���
�s��VÁ�Q��?�$S�`2F1ޢO�@��ot��`����(� ��Å���z���1�Oٙ�� %t�ٔpxڼ}��_"ݱ��Ģ9����+���=����t������=}?���_r�kj�8��@BjwSE��c����˻idG���C��a
����/.L����d��G�sg̲n++�mst�QȩːH`&J�-z�� .'u���[�Kҡ���M���+�<�U�,��Vu�\ƼNʮ��x��6�H����z n��4X<<�����e'}V]F(����:���p�����s8�8�d��#�X5,Ȏ�8�{�t.�/��ެ��<�	Nq�������U-6YGz�u�i�k�}1�eԾZ~����]���K�	�)Z�_��i�ҷ@>֙��E�$��H����}��E�G�)n;B $tX[��-(����zUi��I�Q�:Yݹ -NSn�mL�V�+Ix�_mȺ�s@��X��J��ag4|T��\L��(C?�.ȋ�G��f���QM��h�)��%"�� T����h6�7R�]]��ݎT)�2�?]�߇������N����= ��� �RE��?�����,��`���$��A����	d�Օ�� �hB��q���L�׵�0�#YR5ks��h6�}ͮ�_&�p�t�1k�?_���~�r9��N�[�kz��WC���W	k��)�p��A1	ӣ�p��q�5�����Y+{����S'�jv��o��Z���ds�S0K�v~��n���<ml,�9v��+P�蕜��94x�b��aҟ������
6��e����X����]�?��=&�.���=Է=)2Av<+v�i(�#>�l���k]+��Mo�[;�㧛(�d�BUq!�*�K���5/k�f>�L��}���}��Q��Zo�I�&��/F��ΚHʥ��}�0^G�����~�)�x\�����:�B�S�N�p!���+�z����I{����]���g��cT��V*+��VΚ���c�Aa�n�qZa|z>p;rf)D��;�4�rbu)��_F?&���#���椑�O�����>���1��m�nG�1iF�]�(���c�l���Ig���RY����8!i��
^rA��hG@<n�.�vƈv��z%�1�i4Z0[#��
� y�Ƹ����̺��]G2�4Oe,�./	Q�`�2d�SP�'	�f���괺u�&SMϒ9c��Og�ݳFǹq�p��yu�]knȸpb�4�-R�����x��2��p}��������S��#��GXs���^����H�F�i��r���Q�`K,4(H})D����v��%�8�g`�f��;/Mή�y$��A��J�`h@����f�0
 ��5]��
N��o)��D�vҙ1��=��;o��S���{�;֛�[�F~�u�w��zC����;�`��KO� �G"ۖ����}h���m�����/�G@�B�$]
L9�f�ŋ�iλ��Ox�`\��[�Bsx�$~㋭(P�b�ghDqJ�;��4	�o&��H��b
�O��<HN#�Hn�Y�;�r[��}� (<I����_^(v�*[��V��@�(LoRNϽ~��ӥ��-�@֨^�Pߑ��U8t����x�������2	x��M�`iJfg��c9e/#b�����:�o�[9�`�8�y~D��D��p�iq"~��hi���ER2j�{���(��'!<�
�ҡLj�����M���"d>�����$��/�q�.z43��
<0	b��� pT�2��Q�=L��O<�������O���l W�Iƒ妑D�`��f��&E���ģq�,�@Ņ�i�7�7<\q����
J,�1L�[ ��ZY��7C�o���x.n��Q	�F4Aw<d9��s�`����/Ә�NQp�Hڞ������}ĉ��?D�Z���}�h/z!_X�o4�0�J-�j�ذ	;�(%�1p#M�WO����d�9��V��]���W�j�Դ��R����t(�V�_����<���0O�2a�Y� ���mǧq���q8}��)L@:m���~���[��i�9L(`W�)����@}�&��*��8T�JS���m�z�"�d ��n�/d�x.D����;֏m���B�"P�Q$��3R�͇�� �ll(�Β��y�BN�=`ɱh:�ƧFŚ��Q��Í�J�d��D|����9�=>�z~"��|�9��Qf�s����:g�"���v_ZR2�uK�o9�d�#��䌧�w����ʸ��qp|�����Ö��T�A�6�����$����
�}����1$�����X|o�a��	or)!^?/6�����(|���F��?��>p���?�>F�������?+��?<��+ ���dXP�|��cq�3��X
���`Bû��5f���]�b�^ƫ�L��\�v�������!�66寣o.�>��P��g�J���(Z�OF�[I6U �����%�����%Dk+�g'�"@�����s|���F"Yr��9�,�,���������r�m��C�����cv?�*�T��SV�RV�U� !�3��d/�(�v$��7�?
R���н`4����p �)�mB�߀5r�<A��N��V����fL#&� qP�ݨnxM;��Myq)-٩���/��\u���wGE��������-:|/OEGߋ�\?��3�w�%x��K3�덣K��0��Ï�,�&I��V�N���W	�л5s�W����`�S8��^!�Čx�my87l_���@02~���L�Xп�/9\���w�>���e}���g](�~eI��Z��)��=��啌O�/���(�F����܃��T]�����R�����]❝[�j�c)�=b㚥e+�~��;{�����8+)/K\,��9�'SI��贴���y�h�})t���Ab���)���E�\�׮t#��ŹL�>R��;kTU	�#Il&~�v�~�U���b��j�-��tbτ�4øZ�	�2R1G2����Z\�0�M<;%m�7^�aC���H��� /g�ڑ�����؃wn��)�yE�D�5��0�M9�<4�0r�"BN�ce�U��
W�~�jN���8%�F��XM<TF�\a�����7h��c6�:d��[܍�pyG2�:�քS�����!�*%I�f���>8�`���u}���o���ճt�c/f�#�Pd��ë����=)��l�dK�S�I�h�$@�:K_����=�Hw���&�WC-{Tヂ	�'\��K@_�v�#A/>�9���B�/[�J�����X�X��h�L���)� iFO7�!j�_�V��":	&G�Sȇ��'�,��GRQ���j�B�A�y8ª�:����M'.)�05�E�b��ے�N�vm&y)�^O���|*���@?5�<�+���]_+嘣���)��$���>�| ��,Z�a� Vu<�L����o�uѤ(� ţ��G��?��30�"������� ����p����͕:��/�C���⨵�0�����m�>��ڪ�͔���b����q+����<���P�v�0�u�Q&���Z��?4�1�Y�*9vd C	J�ٕn6V��ɧu͛����a<X�	��ޤ}��)kߟ~������x��H��*�_rPz��<R#��m�pK���Qݸ�׶���Ӭa�a`����*�����>���5a�X����G�eV�-|�x���b��3m�*"@r�H;Af;�B�*~���P��R��)ۊ,W/tr�{��RD8�ş��xx�b3�0qE�+ح�'O�3ԯXS�#����^�\�]���}f&ij���
Q��#L0A1v����M�ą��6a�L�f�P^�4�+�$�Q�$�/rGQ�o��������@$��Λ"�r�G�����=��Q�\,��AYF��r¯��<Sk�XK�
P>�����Fl�#���l�?OO�X����Tz�"�w:t
-�^f������n������f.�_�|��Tb���;���)z����U�����8>�&�&/p���b7�p'�J��*	JV�J b�ܒ�\��,�}N�J��76 s	6��J��}0��ef!u��Y���<����_�7��nE^�Y���g��n�����iH���A�w�5��}�5Ko��0��������Q��A*��9j��,�q|�\���o��^���	��&�.�U��#��e�a�f�eT��-�HOJ9v�F�#e�d5&�sL�m<�΢#�{�
Q~���WRe��9Z�� �H���})�R@�����̏~�b2�"~�
0h-_����&���SL�L��9[]��{ё� 	4_������Z�At���$�!�T���CH_������Iv���]z���K��.23|��:�zq/��nX�S�2;ॕ���J$J��ry��͙���
��$ ��]��8�{�<[��6i��MF@� ����Ί1`� G�P�8�H5�L�^��QoR�
N�N�b f��s3P�D8����3�XF'��3���֒���{�WZ�V��H�o�z�X� �9��o���5�Q:���{;��u���LJr̓#T�z�n���v ���ԀA���k��h/��	1��|ݺ��l6�DXE܎�ЍdϞ'lB�Y�?)�J�*�h�0�AX��A��f�,��B�Ö��$�_�#T���x�$E_����W��zr��0z3#B+����h��ѐ���g�̉�k���XQ�s8a��;��
�����Q�#L�����)J���~�d/�э>e���a*��%@���]i�Ŋd�X���4o7j\6�y�E�^�ь'D�W<l�8�k/g>�����
��,[��ِ����
D�۰[O(Hٽ�VמsP97�,��[mt��;��s[�.�4j�y�+k��'<Ć:��~�Z�s4�!<�(�gc&p��T���G�%�����>�Z����Y���q���a0џ��fio,u����������ݦ�^���lrJ�ْߒ'Un���Q���7}Λ�/��A�6E����>����%T��ڪ�S�տ�w�p��eĈ�o��$������څ��W����<�)�7���[D'��:A,W���3^L�A��?�PL��U̯��$6���8(f%�*���oU�-�}�-w��t
40��(=k�:��j�m3-���K4���}��ܞ�����Q�Au�ԓ�A4Ӵ��s��t�u�ۘ>�r~r��� �:���a�Od�4�����u<�ɿ2ѣ�P�AJ5J�=LU�|Q�����}�zl��y��Zo���C�/��A��?�e��o[p ���"7�ہެ�ӷ����ђ�����߿ږI���*�����������ϓ�UP�5麟J+��g�Lu��;1~)���)1)<�d�}�Ċ���0��1�ųl��c��� W'�m����6C�F�ؘ����h��U�R�K徽�[G�/�)���qɘ�ePxS�l��_n�j�i�E�B�@��rp����WP���e�~h�]B;��D�����]���I��h�n.�6��?v�#nggk�_�H��laŨd7��-�|�� ����f��N�as=%J�.���A^!z��ߥ��i�z�����J�;�iS4 jb1k��9c��-p|���9Q�՗��=�.�߬����MÅ��CqC���)ɠ���b�3��RW	�l�-u��$�J������n��갳����b6M�e*�O!�?�N�S�m���$~�5�O�#W�%�t\+��E�z�5�c���R�À�� ���go�/�r޿O�&��E�8�Pk� 3�t-���k�����ߴ@�e��d����K��d�S����u�0..ʾ����i��$S?�ޕ�G�0K��נ�� ^�W�1a��ٺ'-R����&6��vw��V���"l���"$G�ll�1g��Fnd�6�gBì��j5���1��^�@�>WK$W�`2*s�؂ӿ��oi�t�x�u+fKz�-:��ۚJ����B� �=����f�Ju8�)��'.;�'b%���7�����0	b���(����s�'��y��u,�[���̧���
��p|]==�[#�kg2�Z�뺠n$� ��G��~;��ɾ�3�"^�� �yk]dO�Z��b�pW���`95�ߖI07��� -��D[�P�2��+-�n���%�:��0��� x=
ۖ�����cQT$�{�2͋�K,n!���3E��pd9F?��M}(�O�r6��i]�J<��d>�wS��;|r���q��Lh���{D0� �αP�%R���峯l�O+��jp����:B6D�B��	KL��q��\vT�o�cY=,�6����\�$tW��L ���y����h�V�.�VWr�dt��J����̽K��W�#��Ih/�TJ�U:������#%�� �y����j����ט|P?��1��~8_��!��-������.���׃����C�T�acI
�n����%�o�E��@B��w����y�U ]���ha��F�V���G �g��g��{�^aUS�����w�+m��͌�X�����v��ycVA�?[��*��4\^�h�U	] ��7��X�d�X��`�#��)p�#�K����x�J�����9����x�F�l}г���$Fک�z������y�6��c���}�B�����w�E]�I	��~�
�Ѹ���[����s�ۖ�7��o_��U I��bDB��Q��1@3��Z�W�z���>���hC �҇�|��� G��!,�ioB�(�hB�D�`ŷ�G����>����ճպ�̔�5�$���E���$b�\aR�3�F�O�c�k��:i(��./7!j��'�X`q�ɸbz���x}�L�j$5�� r��x0�%�7��PMdpŰp?F0��T�#؁�q<mod	�j�L_���Gn0'�&~�%nZsa�^>�Ά�.#���f2�?�}'��C� f09�<T�����6�>L�dz�Ĺ���k�$��L����|��dAX��o'[�y���aʃ45�<����Y{y���K0\tpS^�����d�&A��o�f���Z�?������=��V1��e~�!��x���>K��d��]��s�C�?�������[?FD�D,��>���QsN����bT�ɵ@�R�-���aaN%@���dS�h k߷({K�g�\���,Dß�1o�=.~I��qf��D�a�h�����"����9,r�3���@�P�"T%cv�B�<���M[��2l�`I�I�5�٦r,Ћ���2�p|�Z|0���
�w������D =E�U���-*\�k��������4���eQ����;������+��1� ��c�,��m�����*?��gEtm��,�����Vpxܵ�ؾ�$���:f+_�C�˾��g��m���%N��>�)����4Nc�0�x�����*T:}oC�4�UcE�S�	.^�fRl&�ܻ�&3�Ʌ#i�l�^��
lg�#�$�/~ob�u�;���q�)_d��&݂���EJ��>��lh
��v�����v��LRuQ��z�bV5m���/O�Тҡ����=�2z</�|D���#ӱk.��8���*
V�i�kд05=�T��WJIF�)��1����rLj�6�|��pL\BǮt�//� yв�2� �`��ݩ��V��~c�|�t�D-5���[�!��8����d��S�\(-����*b��_�m�l(Y2��5�oF�"Wq͊>�w��x�=�ݤ4e�e���wp�m0TP�p�[��hBfk���^ʥx��&7	���~�M��ۨ������d�K���6y��wV�Me*v�2���u���9���S�����"���"��כ�9�;��X	��
��F̘7�U���8��<g���$�5O����:�����UD�YN�HM�ԿT$����~����,�m����"c�y`i ����GI<mz��H :e��w��+���ݮ��t�����mF���n�� $�ͼ���\V6�1ڧ�ñ�йGW�����F� {m��>"U����� ���A�ăK���qNGE�L�3�Mzs5~��ts�QѰMFe�"�D�L��@ rdsX��x]��׉��[���g�z��O"��@�Pi���4G�j�)r_tq�|o �0�r�6�	�%?}[�58�ڎ�U��V׺�݈���>r����C���C����u�(kU��SL�Ant{�`a6� .e vZ<v�6��#�~� �f�K�A6���E,x0FXD��7i��g�3ef-�\�'�1f����j�w�q�w�J�Y,~��1*k���O`�L�������7{��I��̿K����M���W��Q��$u����&I#"��+ʿH��"q^A֍U߉��qӤ�p�C�:����m�20����S���K�Y�|���c��}\V������y�Ғ1R"qЧB�?�<�����7�=�Q�4vJrUw�Q�CE�Z���ˣQ��.5X�q{,̤Og|�Ń4?q�*-��sE�5�������������� ���TW �l�=����M'�'�Yteؚ��D�[���:� .�[����E/��x��~]���u\�6��BB,���$㚡��`��BM�w�y����t��D�ж���6b$:vL���wk}��_ ��2dMXVI�Ub�[����vv��+�D,�$h�Z0=����v��O��PP�~�O'��5��O���Kq�Ѝ:?�@TY�[8-E����$��K�j,��W��;�i�-�Gco��� e�e ]��-�6�_bCѵ� ۼ������DC�sYKⳒO�?��i����)��p�q�0�P��������bb�}ӓz9���=�sqW_X�dbO���
�=,�L��Ud/����|�`����o��b�7g�;k��� N���C\ß�k��rQE�y3li�!@&���}*��IZ�<OC�tǟ/�Q?V����0a5P���|m_�����e4�^���'s0�؋Mg�z�E��g������&+�F��rHrW��<l�@��:�J�sI��z�>x}/\'��+T����2���I����^|@a��L�e���4H�Ȇl����uo���̗�~�����?_($O� 5�UM���:|��O�q�'�
�l2�o\�B`֙ }��q����pl*w�u�[��}���&^���i�jv��L�v6 !_�<r#V��ݥ�*B{�F\Sgh{.
�І�.&]u�����:A�/ե��K;_'��x����k#�\�]_33K_��|�rnA&\�t� @�.T���]C����&����H�tR'�B��u�cÝ������
��K)ꯧ�A�����)�[��U�A��Ơ�{��O��S��jq�{�
�«�d�O��:x��]T�}�^�����i��S;��>_����~Eۨ�Py����<�l�$�Q����b	@o���b�!��@�.�]��kv�MHH��s��a\%swOw�sg����.�X��v�1����	���F���V >0�D]D��T-���\�X#�Fsx�?Ӌ7���*��hYB��־��+ot�$����:�7���a
:�D^�6sK�e�kP��X13z����0e�$��z圵$p��?N�� `��F�iJ�O�*�兡�LAg���91��B�������4h��-��t��&�Y~J=R�i7��jN~�z�׌%��Kk�ժ^�,�@��u�S[!�̘O]#��y.�ܨZa���=H���z�RM�&f�`���H�T7�m�櫸-�/��K�����1y�m��㰪�;b��.�"
>�y��J�C����;��]�B���O�3��H�C��F]n�����\�Jʜ{9"ཏ�D׈6�[�otz�_����(�����g���- �s�D�l���m��2  �n����@��s$&���)�[鳒��\��'��s57���9��ϛ>�(��A�����Į4�⍿_�i%Z�>��I m���~Q��C���#��&����|����)���i`�o�Ӝ	���u!0p�&)�o�����n=[���j.�kx&b%D���� �ܦ�Ar%ji��=�:3�0��ǃ9cش�,�U6>���ZaE*RJ�����D��r�Y,��ҝ*��2�y�I��X���!��7\�`\n\1B�փ}�0$h���#Y	�7�J��n�<�43?ގ�{φ�����z�<��S�i�K�#i�W�n�W�ꉉsu=�4]����Yf�U��Zb��!�/t�Q�*�,q�1� \Px��jJS���;DJ��;�xH)y���~��ZW	4D�����8h�p�^t`<���?�%�z+� j1�8��e=	�?\%L˾��o��� g�V��WV���v�{�"#j�`�H&,�R���p��Ӡۍk�u�����>{=��Ɍ)��ixovZ��P��)�-��ۏ?�%���;�@�&�(��������0D>�������܇�kY;Ў�O��s?�c_�����m�<޼p_�w) ��̘��B�*]���M�Vܤ�a��f���b��U�y�����L��O�;w ��G��!l�(�
<�4=��j~��?d1��X���	8��ĵ�}[fY�U_���n˚��l�_��Ddߙ,B��r����������L�d��m�T�u�w�q�v}�myy�j8G׃O�<l�D%ms8$ݙN��n;��vɗ�Z���Lآl��:`�F�`���{�Y~2�u�7��q�m|yOKt���|F���RWc�_��yv�$jkph�X����Y�٨	n�o�gu�)�
k�.����m��*p�������Ϣm��dF9K@��֎��C���:r�~!�3�}ׂ���A��3l��H1���ml���1p@6�".�����[zq�`�W������ޥD�n���}L�8��[㘫)}N��!J�^���f�&@}?O�$p(�.Ɯ�vg��>ǵt���T�w�~&��K�|�
��{�w�u��8ھ���^��oI7�l�
>�i�+\���{�L;�y8��~q��Y띯���X�����5g�� \�@��M�6:�=��Θ��v�7��h�l�����x�E�·ނn3OZ��Zv��2�4*4N��m��n�~�m��R�w�o�hT�M-?	��?�#י��;۩�>�!����=�u��z�r1դ���F$����ș�:%-Y2vX����1��\�ҒzW��9C'^0�*�M��3k7�9NQOD�}Q~ߺ�_���֏U<����"˪��6����G����B,`��ژ�H�ݑ��
�~� `Ly��~��.[��3�p3�:�����C����Ԃyx�1����f��T
��k�J�,��������O��]߰����ECHeͼd�HQ�^D7߭�qO.4�����"��W����*IW�'r�9�;�9붸��Ҟ��<�S5q)�����������-����Y�(�LwZU���� 4�?�x�"R�NV��~���	����b-$,2oqW<�i6��`�T�b�;�^����:�]�]ՋC�z� ��희X��!»?��m����{l�PQ!�752h8�&ܲ�C�wm���F���	��F�B�_2��]+�Y��T��l��D�4�S�b���o�����Ffg2cP��t_�����KD,z��$�8�������q�;<��.��J��+��X������:=2>��Ct����n�`<��^���]r�������σ��r>�m>O���"#�D{��"0��׭����Z��d#�����ؽ���w��
��f��d�@Oc��s��A�x�F-P�ۯ|�:�8?\�X8`s6m�$i�Af|���>�����I�}�����\��ϐ08�k_��Ә�O��!�AA�*kp�B�N%{W�<z���
j-�L��@No!�6�u���LW�?����T���&%�,2��y��y�Yk�r8���x6_�zp�`z��4�fǇ�w�=t�Ԉ�b��gW� %p<^�y'�p�VE�t�W��-��
�{ς��5h�6#�"8(��Zk{��O�6�I��"H�zNt��G��z���h�����6Dq3��A���9`�#��{Qq�Թ�ޠU�H��o�Nc�
�6��&6�	�z���Ϡo-+ϞS�?I��i;n���fS˯�v3�YQ�6�z����K�A.l�s�\_f������f/�S�,��l�0�?O[i�"��ʜ��9�	�g�!Mw��Qi�(☉���נ%�,ݝ��}F�k=N`:ZԘ����ѹ�պt�ڠ�����'vҺ��U�|���
�Z��D%�;��@���/��^���=.�.w����ɞ�7E���[�{�uFuSjx+�j�n�(`6�	�dI�f���ʷ&�E��*q��H���FیҗG�%���YJߕ�?|�7JF�'��arE��&��<Y�	gk��M�\��w�1?�F^��ϑ�����N�sme$�1����e���=/��1��F��}p�s�q����h�;j�z��+�:���X��O����@%�Ҟ�O�ܳ,WJS挸��sg�x�=�{���ځ΁�3d�@R-�����{�V�5B�Ϣ���~���]�h�B��K23�\fj.����k����'�!@M�����{ҳkf���\s"�g����u��l÷e@�/�V�i�K+�Z���],/9�SK���^��>��5{S�<>��=OcKyѣ{�.�LP,�2�F�ᒥ��
�R��*7��{GA��?��`di����ʍ,xm���ا�ɣ�ѷ����4� �����|��u?G�{a��.�I��p���dݵd�W��f�x��4�^ 3n�1�(�\��覴�O�s�����-'���q��y�*d̵�,ዣ7���
��;�M��_�!�C�@��";�߻��U���.���;��ד٤�ϻs����8cv�;C�ί[}7�0 ��{;=�_V��K���_��8+kQ��t?xI��trf��������7}����O��9��k���"E��M�xV���R��w��BfT(/iq�0��	�|}����v�T��P�ּ:VJ�NS;�DbwzI7N�H!�ɽ�;Z����:�)���7y{Fi6�f��rxU�~x�j�\��@�g���b�tT%�&��nw<�E�ܧ	��=�P�XcG�Tl�(̳g���|]�N��ո���+���,�9q��6{�����n���K-�l��.��9����%[�����`�C�v����g|v6xﬆ�]�`ƺڿ �1<�a�p*N��:��w��;����qq�.'�e�G�mFr@�{�תL�Qm�n��H��m���fV�KP��'�-���5���eM��u�~�|@���m/nsf?ڳJe�:S7�e�~� 8(�X�] �#��w���v� d{?tk����y`\2�!*:������0�)�ݒ{��O����n�ʾ���	ܢ��z�2>݋�N����O�a�1g�)�W�O1_��4O�;�D���"�;��E;�\u��ն`��f�%3�D�~S�]N���`����>�}k�!6a༚�U�8�ir�%;�qˈ$Eh�r�"bo�h)^�*k����'�v$��{�5��xC��r�ɇ�O��>�@��LLuv�)�-��nve�����k�o��A���TĦ�o�s��;i�����H�� }R���5�Wn���6��ɀYO���:�������pj��C)��Bq-w�`-Z��w��K�R(.-������w	������y�����2a�${���={��:�w"ʭ��� �w��?�tL�N6�~hU�t]]�1��L�3n�9� m���d9�v��.|��+\�⋎׫�W��qDa7<� �n�,�m�b�}Q�#��V�]=9/�R���΋W�Ϭ�_��;m����3�rS�8���E\��/L��|��'fهtna=a;�ʪԭ2W�=a"o>1�aF|^12�!bZ�J-^u\�h� K����Ѿې��D�2DƳ0��5YcH��%!�=1A ])ĚNϥ�L_���F-�(E@�g7����94�W�y�3��q�T/�>4��dazI����D�U ��3��B�~����ƕ�Ʃ$z}K!�{Z�0]|��r��M�h}�z��]���1��!i^↹F0M��(�9�ǘ{]�pU�&��gWС�E4@�=|늵ݱ&n�t�P��ۈ���C��&z_�1�8�}.��d\򆀭�� �	g�i�/�J��=̬��j��8�� �<��+��f��r_z>�ʸ�g�V�̺�ş�79?[�D$Q��_�G��gM�D%�&��y���Y���oK-V�'�z��6��w�z^Es�n�]�ҩ��}?=��H���FF:<ig��̡���%~9�m� "�l(J�a88�*���喗#r�}�	�?�	�.|���	�� � ��q��Is�cXLIŮ��($,�f�|�L)��-�K?���1��Șc�ZߩM����ݝ_����j�iH�1��z	��ٓ���r��W�k����Os����$���;�)ෂT�F;��c	�s���12�>�*mk[�>f�\b�YX�|���+2�ƑO�.��x&��o̊�hC�+�w�E}+d�[���:�ڍ� ��WҔz�iߓK�g���\~w<��C$�Lg��g8���f9YK�|S�\�Uy�$8�e�:Û�|x[����/pҿ�ּK.8�s�ؓ9\0�����Ȭ�~�;���AEU�ʡ�
������:k��GԒ#ⰲ���A�[���j��/��b͒��o[��ل4�qx�����Y���B�|T^gON����^�Н&[V�ʞ�n%Uw���{�����˝�v��Yfѧ7��,0��Z؝'"�-b����8���&}H��%Pywl�B4�9-�U��]�����Ϸd��5�Y?/jJ.Z��2jf��Z,�\����a�gw+����� �?����8#��1�����|��C��L���V}�1�O>Ű�g�e�	���;�̿э�ONyf���-�\��P�\�ڀ�@�%���v˯�yjݱd[�_�?�a�W����s�ڨ�>3�i�`�{�&���XSBs2�)N��A��y�W��;����m
K�E�I��+#�l(����U�5g�r,�f�Ӂ�	��i��d7
����v�عj3*�����I|��I�m+��N��W0fJ6��65V�H֐z�N�T�	�f�͓��q��諒�PTw��P��4Rm���B L��G"��e�]�:w�P��9��h�>������Щ
��8QK̴��Ѹ�5m�P�I6��%N<�\���%���V��xo�D �S6���P�_�de�]u.U�&��c���/��7�4 �T�)���3��]�3�j$u����ﰎ�Q)�T�8�93��н�k�����,���
��>N��'G�+�J4nx��e���R�6�/�"b�\��~����8��X����Mm}�Du�E;�L�[�?!C����`���Ԙ(��Ŭ�������������#`?� %�����k��0���Y���Qb����QN�d��9�xe�+&���b�7q�]��9Jw�wAf{n�(�B/m@lC��%���Bȋ�û��-����ͱ�y��(�H}<Z�x�k�u!�%70��!hY��U��W继�5NS��i��3�ʅ�e����Nx7i���.�ἦͮW�����D��O⣮����c�%&�����w4챕]�9� oe$d:�����������q4c8���ʜ:� �o�+BK3���n���U�
ab���+߬�$�\��A�g�T>�#h�'��<&� ���g���Z��}`l�~�����n�V5�`���>C3z~p��P)X#���x�;�jr�d����=�^���g�oR��:4�%�P�ڜ�Kqܬ�O�iS�s���7��e�r�j:�z}�[�c����[�n�d�^�a��z3����QW@H��2��g�f�d?����[=���1�>���[���l�- C��_���r�Y:͕o�\S���|��-�2� ��2F�?M;��m2f���������NԈL��
I�Z �������sR�y����r�$%*�˴���@,�,³�+��6�,���Z`.�x�yH��7�À�Zb^Ҫ9䄗���#��Ԩ�S�V2uQʭA���vm՝)��)�v8I(O�s��O�&�)�f]�v�ˁ�(t�E��ف���eK;�bԕ����y2�(5������ܿN�t�q��P�Ys����t�a�T�����F!��n����Y?�2\M����{�]��Dk���Yx<��8[�d�2��V�mmq���|�?�Uc ���2��"���w��=�X��X�����ӑ^Gׅ�:�>e���-�iU���:X?d��K@l烞fOu�v�ޓ�}��S��d]��9�����!�،���	ø=,���y7ţ=�#R�t���9x�0����%=��H��0~��\6<�үYo�K+�u&�):++���s�Z�U_i�6���, \����t��DW]���~�r�:2+d�(�H��7�!<�m�6SŶ�z�D�"{!�0\*c�Ͳ�'��I��Ue�vW�Ƌ�����Ե�Z�p��*�)���̢)�����g�n��C;(�&
w�U����&�A�r$�k�Y�Ut��~ܝ�胠��E�/�Ҥ�'�qB$���oJ:\(���i��v-�y���D�k�����պ��t������v�1>��:�{�/�����G����L����w��oWv�?z]�	ޓ�ZVO��}W��؎|�d��+�����3����Gir���Tٙr$�����f�r�ny#*$�M����!�%[�[��X/G��^�R���Bpv�¹��� 0i��}�P��C�a��Iّ�v���X �Ii/;B�!:ё��K�������}��cɡ��ֽp�9��7N�W^�M�������Y��4�����z�)�wYs��
 ��|�9gϑ��̈��⥂j?�,-r���]5z�����		�����	����H�m��T,]a���7��{kQ��PI�.j�`y-�K7���T�+B+nr��xM�v�-"�/&،���?�c1�^˹X�vj�RP�9s�b$`��N�M�3G���#��dq�x���s�|p���t�����R�"��,�J@ʅ�:Ҳ�$�PP��҇�j�.J6b533g���x/
��9ip�V,�R���^���;!�Y��&�%�h��n�A��&�|���*{ɨ��,�����ѓ���e��b?���5[�xa�\f��[<� 7��BNSf�R�sr�q�'0�������s^�����*k$7w:Q����;��?�i���]�\| 5(4�R1h�`�cd���TD����3�T�}w~w��3�1_���$e�=��:_(K�����]�NH+�0y���M���ܷ-`�[����E��O��˭W�G� �&z=��9�G\�&��,^�0W%8<ĝq� ����s��l��qq<C?ю������z�:��1�Ug��Ӱ�;��L��G�_v6���آ����e�h���K�gC���4����$���1F7l�m�xA��u���݀���r�MK�@f$Q��O�W" ��g���N���ȱ�I���JlbeN_(*��ITMV�����iW�|�D���dV.����붭.�AZ!��Ț��� ^�j��k���)���$נ�ED釻�~����¸P��� e˗~W��>��\mk"݀�}�3���^WT�i���f�{rDbX u��n���MW�.�2������%���L��[���� ׭�\�d=<=a�7Z�&��mv��(�m�?+�'�1#ϥ(nL�ǲ��,X�Ҟ���t;�*s��iV��JNr�)�hvb�����m��j	y��4	�l�2�S��A�ŋ��v+;�q_��)����r[TƵЧ���;#��ܞ4諭�c�`&?�A�m�!���J���{����V¼�v��0g�Q[���� ��ݤb%����uXIn���A�W/mlpxp��X�?�~i��R��������Ŀm���t�#��Ǵ�ZW}�J���b�l+d����@x�
Cs�k��j��D��Fc����!j�9ŮݷQ���lM^�&�۱�<�3����^��)�^6�$��]�s��(��ƶ�����{��A�h���fnO���X7�D�]���U�$�Ճx!���w"����ކ�:�q�K*��{�CQG��M/:�a��vʖnޣ԰�'\���C\E�u}0�)�l_N�s�#����z�m0�t$����w��><�hq�)[Rdm���Rn[��W;K��/:���#|>�x)�4j<Oz��[/�+��A!Z���~^�~�B˚;��Zj�!(�<0F7<S�s��,�H����3�)TM�I�I壘�;Y �>��N����0�wi��*�ʊj�2��)д�w~+�R�~�9��D��>׸mؒ=ƈKj�R�mUTC@ou��L���H�5�\������E�b��(���5'�ޮX�������R���z����jLU����m䨞�����e�qoJ��.VQ��Ǽ�j��[�_�|�����8��dx���zV�7�/B>=.�����pw`�
�� !d����57@�� ���&���Alr�ݣ�O���f��4�Q��d�5g�+��k����a#��o�%�؀���0�k��y�Ń:��`��'zm��׽���/D}jDV��$_+�"���~9��	��E3ק_j���&DĿ��\/s���?fQy��3a �l�x���-O�3z)غ4��]ĲX���zl��K�#H~���!֧��̈́b�b�����]u��R�Y�(�����$��8J���E2gU�1��u7cJ��¼��@+{ ��Ғ�Q2=�	�j��f��pB�s�D�^=,)��R�ǃW�9�,��
*�Ȝ<^J���[L�7�ҧ紬��W���p!�v ���I�!�ø�Kw R�zU����/�F4�p��|�A��e-�kJD��M޾��	�}�e/_pc�r�o`-:����p���;-�ۤ�c��0*����)��2�1�A���UG+ͅ���׍�r3��[��M�`��˾V<���&��@��k�V�[��
%��3F`S �C��C;�UہLr�m�g���b�{Kj�!&�SSU��!� �F�6F_J��L��Ʃsl3"y�
}�z���"c��x��R�':�3>:�a��?==-�<�;r�\��R�]wSъ!Z�5f��os'1�z�p�Pk��Ұ'�s�:��ĩ  M�!�5|q�3��Sj�ɦ�w|�_V?kr�oyo):��U�ٮ���ؿ-	v\-ז���٫����9qէ%Er���a���0m"�öl�I������@�eMs���~0$��Aʮ�� ~]
L����?�Jl�ȭ�S�a��D��j3�zܴT�u:l�"\N�4-���t���%��u����}��l�~�m-	��}�h��{d�9v(����Z�Z�O�uDp���1�ƽ�KE���]�'�^�	8Q�0�����o��w'����_	D�u�DA�_���~���0����|k�����X��3�,��A%+Kz�+��x [��~�Sv^C�D�@��8�������cK�1����R�ﲬw@�A������m%��o�֞pk��c��r�ڮ�KiяW��fi;�����9m'�9�];�{�fS-�.7,^�����RwQ�-��j�r�xL�X�4�ܲ1�cU8�Ȥӎ�'���lCx�|�ϐws�W8W��#���c�FB� >2���*K����m��2}����;rH8T,x�.�n�~36Q����1��p�<�Д�e_��	�ީ#�	Yu�>3�K.��.	�+�q�1{�A��+�����2�?�``��#�N��l���������A"��n�8x�Kür��f�1f�΀t���´%\�:�:e��2'��$����-X[��j<����k�uD��lJ���%�u��W�Cև-�v�����f���r�(�����p0k�RWsH+�װ����9]H����R�3N}����d�i1�}ǜ����qڕ�R��_g��X}�J,���ν+�c<Zb̹�,���:/�S�޳K�U�S9r�J��;qzoլ�8�z��@ �>�����'�o��L�'�T�G�l��o�>R�}�>9���w��&��)+��[����c����r�l����9�����lP𫯭�#�g�m�|�)�:5���ou�r<,e�`\������7�~"�F�-��)Ϧ��	���P���֝]�9�-L{����E�%����*��B�XS��Ȩ��F����y��.Z�m��EgS~�\�y3��vD��g[��SN�H�ee�	!�J�ⳬe��oz	,�
�]W:�01_�8���m�q������YJƏ����8�
���=�?������u�(����ǡ��:��N:
���g��4�m��@J
���6��PGJ+�x��d�·8IۙHWϲrt|;�a���ώ��(.��r�s��(��T|�X�\*}<�����w��fg�p������q��M�X�ִ��$�s�"�w�����_��N��tt�ߗ\��+�;ʀٳ�4��j��V�+�+)H2!n��Vl=a�^w�l�&&��/�JIa�g�>L�to����Q_�a���\u����eN`ɣ��#4�"�,T@�s�FE;�?O�6��@MJ�΄���w#ˊD������G�d�t+�~�?�j�+�!�D�^cc
�f�އ�f����v�D?�($���H��f"�_�tWH���HG��
��*L&!�B �]r�Kc�AlS�K�uU�_)IE���W� �/h�&/ڣ�sl	v�ah9Q��X�����dr��Є��d�o�>o*��Sr�>�٘�Ѡ��q����q̅�CB�Y��2�ǖl4c�PK� ��t9Ǿ0��꧙�Q��n^�U��Ô�Z_�YQ��ip�ؚ^����o3I��M'��;Σ0?�3��f� �t����kS��_t�ў�^H�u.ƧB�.7�\@ZC7��r;�D�싼*<B�}�;Vz�� >߷��ΰ���K���w`�s���8�̷�=�z���%�W�Y�"�\�ǃ\�=K�9����~��z�C�d��-b~��G�e�F�|q
�O�IF��'��w{��ss^S�������v�3D�,k���u�6Z�9y�*)*A27�D�}*�jV�ǁ��0���������q�;r.�����̹I��jf���,�{��O81/-~�������Q�޿L��	H��K�kOUT���[�=f�D���G߈ʿ��J,����a�����L�	�jW'�P+�8����ˌ�~��_s5����@�~ߜ��4�p>���Vj�A/���ʸ7� ߂M�K��uN�:�Ƙs<7 A����O�R�ez��{��"{s��$�q��2DN�r��*"�8��Y����WJ�F��ԛqi\���d�<3^j
c���~�u�$Z�J�H�5�n�f�/�
+�v��V�-^9�F��3�Gm��E�F��Q��ߖ�9��W��u�m�����[�߁�'���"�ȄeΠ�v���ed@�*C�K	�}"�P�ř��Dv�7$�h{rx�׮�r�;�.�eh,W�@�2^�k/�;��"���iE��[����L��B��+���0 ���1�_�i�J�b{���LW[��bC�U;�{���&��ŭl���O��783aB�KݶU9��#��逸H ]����[�Pr�s��e�Nb��C�E!���������?�wx�pJ�Eat�a�?N�*��s}�vֳ�9k
�W�q�H�R�-�5I�0BǬcp��-����w����9��U� �}��6�J�s؎�>����_�voh��c��~{�����uBt{�DC%N*s!�|���l�zKm��E⾇�M� ��O��tsH��Ng�V7ˏQl��=#�7�|�����9հ�؎gbS뽗2Бzc7��U�p'�PV�;�A�Zj���(� �*"��n��xY�(�0f/v��o�!K�����89�[h+-i�9���ۏa*��Z%.�L8kcv��k;kG.�"����H��Ը[���s�������NC�;���d�vzT��z���m���u�T"	�T�x�Ѿ�x�ūD�0�,�W����z�P��"�A=�+�&���Os�3�K{�uL��wU�C^=�hg$��H���L�<�J*OA4�=��5��u{�` F���1�x>��������4����,� � ��p٦�]vff�F�K«װ����d 6�5/��ۮ�|7��\���K�f~��ץ=���t�,�yc[)��Ln
��q[ڷ��"����})q#	O��{I�gB��
)4[�6Î>*+�vC\�8��?�.�+l�lQ�������!���n�>0���Y���r:Ż]� ��x�~��U_���cҭw��8Qȣ�kS�>Vq�C��i��_,l{y��]2�n�~� Eh���a����O��+O�L�B�a�<���nіw�pt�=
���^�p�V/ݍ��D���GJ���:x����8�L�颩�s��2��No��v���k�j:�Y���}�ʚ�����E5����������Je��ѷ��U�|}����c+نQ��`��)�I���CO���ݢ�|zE�X	s��J#%v�?L4�`�
��|'��ݨn+v�%�l�a��0x� ���up�D�ͅyˬ�o�͗O���9fO�?z6W�Di���yJw�іo|cz��}Vh��w~wkp��CA��h�W�d���F��^�`���K�	�����n>��{�+$�k�t��g����m�6�7�ǂ>����5�4^]��{3v�9m+@3=��y�<�K��tF�:�����`1EI������S��?�f]���iG������?���\6܉Sfd�X��s`�:��m�N�_���a�=��MEt]M�e��*J�T��>9�OuRMY��j M�Tj��	�,]G���,�3�21.<b�ǬWK�#�ɨ��4R^
>V�5k���J�JiN"���}�܋�Ƙ
�[�ƍu�d-�ΘӰPW��#5aF��G�Ht*_fT�iT�68q"V������`>j�'P�M���[��#��zW�7�--0���W͝}?�
���ϟJ�w33)�	.�����e�p�ܫ�{��|��&so-t��Z��c�=���z)�����jR��g�����u�XՓ��.����D�[_9"'��������)��=�Ic�jX�ci�	w�wr@>���ߘ#M&���L)R�tY��h�+1�6t�d��y��"�5� �o'�y�	Si���ƷH��jk%�ğ�����*��2v����%���E�-C��t�7�Axe���b;�j�*8��^�~<�����9rͭ��.F���Ʃg�6Wbw����%���_��rRiLnK?.��AV��}�o��� A�)��Dт$?Y�Jy}$�q8~�q��wum�d��]�F�֩|U�������8^���^�Q�F�FՃs���(����F5;��fр+��ǫA�,s�UEl���״|!N��1Y�������
VU��t�7~���G*�9��y�!?�u���"Y���A����7����n��Jl��u�pV���B�B�-�`v9�3^2,���+b)�?��H���A����<���w�*5��ݫ;���Qb��?���b�1��#�>���3�2�x� ����F9W.4��ȕG��:oer)T�{�*���'ض|sڟ�ghvj���R��P�E�~Ex��K�W�[!׎?a-a
5E"�@�
_�48��E��Ru����[k�a>�L�@,����\ƙ��E��:��`ZE����(ل�?�%��o�m��[�K���5���������+����Ge�����r%R X�zk�hf+i�/^x�;��cm�璠��c� ��W�_f P����r��#%`N)jR�-$dǪ7��%:8�s0�+�o�}VI伆rܝ-�V�	ˠ��/a;��F<֕`�T��T���n�]�O[e�_�k��Nt�]$So�Զ���ɮp��tE��A"\��v��E�^��	��y|��j�]3g'D�K"�mX�ɖ��
����Y����CU��:*��tW�WP>E�G���ɵEc��L)��V�~s��}p��˫�(׈"��	c���X��
��x�	ޡ��Xb�7u�1�R(p�N�^���yv-��N��{,��T+�{J��]��� t�j�l��m���u��(_p���8�-~��@�����+�u��Xr�v�}xW|K������K��e����Vr�:q!d��%�wyi��d�͎���̽{2����K
g^P�~o�>w=�5�B�9�ư�!��7��,g�A�ޖ�MmͶ��o�g<n�������o�f�z���~�� �0=m���F��E�� ȡdjiQ�������"Y��d=�Ƿu�י���H�X�y�LMy�@hO�� 2�dH{*�]I�!���vwȮ�>i��ܖ�I� p��֡oa��'d�A����+%=�o�����n���̾5���b�k:�H�lq�補�G�D�G��=���i�WcAW���6@H�}��!��~�N\�WQ����,d�*\P��uq�P�:����w��x?��4�\�:G�M���>��ֿ��'��!Q�t�<y�m<b�pz*5�d�l6�� �H���+7�~u]����9�N���Y �}�4p�%��G�]F��|�G`�����š�a�;O-\\����9������獫�Ex��ٓ�Z ���R���Ge(�p(5:��n��coN�����sg���G�tHk��2_Q�|���m�)����`�I��q�ZI�o/�C:���K���0�)�0���Q {��FBJ��K�Jo2�����'�÷}��'B�W�q��&��F_� ��(Ͽm�_t�P��T��!���~�������Y�s�E��2�,[��1i���}mx�՛xI 01��0>�;���ε�b������6���>����e���*����Μ�bN�=� P�.�s���~�͍br�I��׽�E~>쩾��ڧ���1���,f�
��$���-�u~�W�/��Z2p���	|-Ad��g:�ؐ�/��hX�x��V}�U)pBK1�����$|]|�]�۪�b�j��TYe�,��-�,��=∅J�Z�o���o��gRA<�8\����8f�Uh�g)Q�:3�[����a��ꕅr�^���)�v��i:�Sgi��r�	�/�'���!�ػݡa�X]ɲ��R�*�}֛b�Τ����Ok�+�J��&�wnU�k4T2��ԟaFAYٛ.63O��1d�CTCp�0k���R��g�w�A
�B 7P�4�M���^P袧e�l��hy��O�
��nN !���$��R� ���������S7"����-$���Jq��l3u�:^J��k�֚�;;�y�yE��0?8B5�?�dː�����sWr���ڐ0޹�o�tWl�l*�\ ���xy�$:�W��[�xYh1��E�Z	I�����a�����\�����|�2eY��*ںT'�O��ͯs!&�p1���yb@qzfC�Ͻ6]l�����:���`i<�x[�<����$�FA�	I�'%�w�r���C
7:y�b)*˥]�Z�,���s�Jkt��rFR�~�4~:#�9��/@�j7.�`�,��f��l��L��JIУ~�00_6�!����h��t%��v�	���/�W��X��J5j|w7�NC�J��j3�˰K��Dm0����iZ��y��&
U�6��E�3h�V�E J���(�MJL��?X�gβ����{�N��D;��x���Rc	���$����>�~��tA����s�u��Q�g?G� �xfu�V#Ӎ�~�Aǘ������Oi�Z��~;�N�x~��I��A�c^�LJ�r�=��P��q1��̹Y���F���A�w�AE&�C����:�z�e���y��p>lp��ҩ�@�;���g+��G�H�h��ΰ�M<{��@�ܛ�ÎT
K�����S�u�R^��h~.��1�<�;���p���uKh�!�k���[���/`�3t3o���k�><s���|���O SB���Vj'����a��@�dX���Xl�e�G��N�vN�
��/����xG�Ĵ@i�ͷ�r�m��9Γ��p/� w�D@IF�A�u�J��УD�׆G�p.픎L񉹢Sz���i��α�,�h\�']�#_�"�[�eBu%e̿,_omk�/�^n�X��)���Wϛ{���۞+�����WQ�Q�VA�ѓ$��Ϭ���$C����|����FݡE�N��'.�0�Sn����/��7��$�I=G�ta�o����2�t!(��*{.}f����ʺ,���+N_%t�����TBzt'']��2M�)�\4�T�AJ�ٞ8a��\*�w����Y�Ak�����Rrْ�uH<Z�0_�-B�8&�q�P`:�^ib��u�[��jq�J�Jl<�	��ǭ��Þ�E��t��UK2a�bi�Ͼޔ�N�`�j�#X�,Ĕ�D0��R{Қ1"?���G=-»^�pn{%��9n����;jZ<�]�3�������<!��OnNA��g&w�������0����-`�a'6^�"��i[��Dz���K����@LA���W�)�D��q!�`��n�2�O+o_�T��Z�N;l�	�6��H��suOuu�w�}苓
=a��1�S�N��)���=�t :V@�%�7����M�pm��t��o�B���(S���c��[��Kۡ��;�S"�N�^D6_��-�&����������5g�z\Z�s�ot���{���p�I)5�D0��y�v�=�P �]�����
����-8����$o u���,~j��M���-8��"/4�>u�[sS2S*:/��k������Fꬓ�,��"w�%۶��ڃ���b�YK��y�Gg<�1��J��$�
��7hWہ0�p�v؈����7KQ��1\a������0j�y��8{�&!�'�n"�t��0|6�	��uO����E� ���K�	{��\U�R\M�xX�ݳ�_�} A)�����S'���p�VhHXx=���Dǌ�;�'gO�qH*�%ȃz�'Xm��d$ >n��:�b��-�e���+s���r�;�	V���_X�<IoP�F��{Sr�7���+�����I6��|��3E�%0ì���R���3K��/����!2�xJc�?#q%�������x��H��ۨP�� G�41�a��*���9An���P?L��f���GS��L��V������ �1�Xcvbjj"<�q'ؐ	@�B!�_ 3�2r�$���D�/8
͖�'X+�@�󉵰�E�%��#�9�=V�[w�xDyfs!�\�
_"6V���M��0XA�)JE�ij�����3��
��x�����e�Ҩ�w<��W�=����.�g��lњ"ߑW;2-��4u��8aXa���_���_�Ã���0���Y$�!?�
#v�\e��g�@O9�K�
l�$�{X����}g�D4Zo�����Tܖa�$�2ێݞ��t��U������'^ �3M�U�z�jN3�Y�2)�tYe��Ӟ �s�90��0{���ݹo�sbx4��k�r�xK�B� �1	��)�B�39%��	��be�����j����K.�|?��S\�/�}��Q���f{�f��C#��s��KU[mK���������˽cPԜ�9���7��TT�'������y���3�i��3,܇�7&}���*�h^��ؼ���Ѐ�%����_��.�ͤX�7��H�ٌ�����f���on((��3�e��Dϡ��<���ԗ^8� ��j���S\P~�sCpp���%�k���_z��^>[]r).�a�=I���|�G�ƥ��ؐr�
ǟ����D� W�t�҆y�ߥC�D�k�e5%O���{�	tt������᝶�h)JX���%��)�W�95[�{����{�t����J�ߥ�c�z��/sJ��mw�|�.n�B�/e�=��fN��+"&�w��^��-��Td�i����}#1K.ɽ��>��}s�IH��Hif��8ϣC�] ݷo�v�����?�ݒ���D:�,����,Y�����Q���8���˜]\	D]���������`���2����nv��u��3�<rw6n�6���������L8�[�(W#5��}�T�|h0��|��K\�4K[RX&���&	��I�	r7_6�ǜ������2C2 uAHr�Kf�)����b,� �Z�t�j1��]��o�X'��ߪ]E@u�޳���tC����v��/������0`O�]M<L�O�E� A���B�$��Q�[jʭ�;Y\}0�^��C?���[o��ᤃ̻�	ѩ_`N�����?u-���ᙕC3���8�θ�^�~� r46IL#U^bT���Ԥ�[AF/S�7�<����,���hG���h�Oe�m6\!T��d��=PΏi����<ǃH���Qz�4v�K��#�%�Fn�xg<��d��(f��[�d��xqs~TP,`��Ζ�׌? ځF��q%2��F�DU��]Jp��X��X�R�����v�U���(�gݠ��OZ�뀐f���@�I�Bx�����3���B�b�<:�I�&��w'y�r����AC����'�O�Ǧ�0;��JL�t�r��i�Z�����%�^�hR̳�"�}CŢ-7�D�)M�'Rp|o�>�!>����U��N�i� ��Aw!��8p<��w𹟩O_�O_�6�Q�Kz�Oi�O	���Xk��:�J��ެ�Цƒw�|�SR���0]��@Z� -ka�Ұ|&[��*K���W�����r��^��$�%��ܗ�j�W�W?+,������!@$�I�6L�&�{M(D"Z �m�����e ��]����t�}������/��V��x���L��ᨡX6bx�i5K�/E>��L��v|8��w�	q�Ϟ�ӆ������9  ���܌Mt�&hY0�-��X��q�1������vGT=5�ک�pX;�\\� ��/����k��+��s2�r�q�A�:J���rSP�����HI!��.�[��ځF��sNp�#����|�EE����Dttt�

?���҅jq�/��}�W��Ww�g7�<�V�� �a�sg�����[Z/���/
��D�� ���,�����z�Y�a}e�:�u�P-6[�%�������s��� �c_z����a�Vwh��q��Dh����s!�^ؤ�*Bg����`�G�Ou�b�
N��6�������%�^��n��o����!�B{�; �7h���⟸j-..����� �`�`���o)i���}�H�_��Dh�0k�v[��R�:^ |�=�ذѫT̏FDB�~�r��]EQ�<n��Ћ��JZ����jEFA�� �({��v�5��C��C�_?ɫ���W�{�k��S�nVF��JE�1��1������� ���I�+�>MWa]=Ud�Q��noo���Z����~�Pإ�
u��b?SLNLd>>z�������ܸ���l=����-�a=����~�|��/�t�EgK�Y��%Ã%͋܈%Ė�Ŗ��|K/ʓ�����>#E0�wt��?e3.�w^�)Z?^ ��ZK(�,���C���)�:}�Þ��狂�~0%qp˥�!��*⽐�)l&���0�e}
�ϻ�R�b�,s�Ϝ-��`8���b�%,�s�=���2��O���/=aax��fwm�����Sn��P��q��;I(���*�1�%v�6�'�i���8�-��_:/����dEV������Z\�.������gs�]ꖣ�	$�	��5�T��U>2-q�lu��l�W1��rV���9�G"U�Xȁ��d�d$^�$�Z; htt�f��_�/���Ҩp���4��5t�[~+_x?y�W����l����- n���~��uu��V�R��-�P���-�#*�,@�P�!�ω�-��*/�����o�����GD}�E�	�✔]��,��v��P�FI�h�Xk���/Y�ѣ%�gzd������38r-#nå��_���gm��z^�h ���	u����Ֆ���ЩW����Wn�Z����abx@�ɞ�'b%Hλ}<.bQk+6-��f|��֘\(_�;�:�?��0�7��`cBA���������pU�At�>��'a�j���l3�$l�|��Z��?D�u\T��=��((��(-�1�JKw�tw��!!�)�3 ���H3�934������~���{�9{��Z���TMV��M�{Ь�:���&�F�yݏ��iY��]R'���B�l9�H�rt�(N�vz��#n|�_l� �8d�a,�"�$�|�ւ�������j5z�!k���D>���3+ɸ�H�]&r�V�נ�`�M�[��HX�,�YU(�}�ڈ~�<Y�����v����^�^aE��?��ٹ����hŕ�[=�S���՗Sa%�Y��Lɍ�5w���p>$F�(���v��`� �
����f�������Κ��<s� ��xX��*A��t�?�K� K��-�|%�Q�[���'>�w{���� >Vd4%>o��J��JE#��M�]�:C�F�쿉/J�PL/�5VnT�.�O�/���|彏ߘ:�j�k�\�J$f޼�rs������� �Y��U���ͷ-[t<7�������JՓ�͸t1���|jl��>*ITؾ9y�	�b��P��ۭ�Bb- ��	���Y�ٍ�m� r����ӊ�N���~@���*�,��).0k�q�Yկ�$o+s;L܋�d"FT�γd���Re��e;��Z�ҿ��K�Є]G\n��D�S����]=�δ�L8���|).�4~��I�m�mh�ȸ1Hq6�)eә�l�[��N!�(8@K�PH�X)0r��U�M=dF���ɭĥ�Sz�G?T��� N��Wc�ߛ�g�����`�3,���������r��N�|�v��������.���<��Wv$��n\��&���'��͈��0]�+*o!bR0t��r�g� 0�;̴?��R�AAS"���Z:�Џ��y�}��m���F�`g��v�䱀{1�r���=;jY*���u�}�5���/M���9kg=%���B�al��)Z���Z�0��
$��ԩ�G_^�hhh�'�ؤ�ch_]�����璳�F��sW[�gd:�)>��$\�u�����$��:;��[�g$ː(�p��](Ჺ�oo�LqJ�d6a�c�
���&;Kv~�� �aG`�%9��)�c�5�?�<�� 	&����d����Z���C�M=B�̱��ͱ:r����&��p��}�����`#a9���b�T!ƿ�W��|vK�&���+�E;��:���+w�~��W��_elS*�U�"k�������U�[c�bb�~݆f� 9]A�h7�8]�fe�gWeW���t�� Q����q}E����O'��ލ��/.L
,d<t�}�k���F$T��Aa�)�>V��-��g����_7HD����}�����y����9]�O�8v�M��A���*ү�Ƹ�=b����TC���	���־��{#���c4\�o���E�~02j0d�t#� м���7��d��`-<���C�M�)Ig:z���ɉ�S��6Ak���w���B��ԁ���wzoI�w��<z�c��������eqR�n7����@��*�W�/��;wo;s�?��fSG���������4����d/_���&%��j!
�rY�(���~l!8�������e����E�&?���.╵�}�:X�{٢��H�~�ᅇ�N�'�O;���yM��*`"���ߔs��u i=��K���$[5ړ��8 �)N�O[�pp�q�����%���{��>�ˬ/l38���Z��F���х/���ZZ:U�S�%?.S��������/��nZ$�h�$[x0�c_f9��7�{��`� �2p��^�t�
s��K��&��y�֩�X���(�s��]��vK��Q&�Y��}ג��}��[�!3�uA��u�]��ϧ�YSo��jɏR�_��YV[��^��_�_���/��IMq�js����%y����FU����w6/;���@�r�{����'��n�u>~1�9u2=OqlM�k�����e�#U;V]�e(���l�R�t��5Y�����G�����r2�%_f/����6<��Y��N�WY��lE� {.\�����p*��ӌ��4����D�s�R����/P�xs��9#�Mp�~�|w�н����8!��w�5Qo``ځ:;��O�w�}���x��j��֞�����%CY!ZfX,�:.�s���u�{�}�曵y�̨Dc�FTȳ>�q�jJE��2���u�=k�hL+<>dja^�����]�
�7=����6��ѥ��rA�rZ�����2���q�yn+;\�?0*��i���� s��Sgh��j����<�K���ܭ�+[�S9��e�N�]N�f�Q�Y?D���8�?�&�7�&���6W���� M�3�mIn���n[�p�%ՌN�/:@�&l�v��[�}Z�e�~���3��)��|u�5B�Ũ��@��ⶋ��|�����LE��TgB��%��7�X\�
����{��Q����̱P�k*+r��c�� HrC���6*����7��`!��/$�lm�d�m��M�h9���=�v�Z+�b�}���ǥ�I����Fv�sESo�������/��!vՕ�Y��PJ	�2l���!��e�OK�l^��m���`Lw�g��r�i_���'�U��!�� �w��C�C0��5��07�. �o7�cG��:3�Xeۯ��g$wx)�֠�UǶ��E=�-�S Gy�a��ۯcnUͪ��w7�=�bp�M�ZƘg���v}��h������������N��� ���+S[� '.�{H���H�m(��e&t/�*/�[��� Q'�o#�=k?����|L����'Y��S�q <Vk]�XSټΌ^u:�,����5D� n��8����X�=��&n5�i����0����V��TbefE�z�t.�dM���&CG˲3��H-?�!�]���_���z�����+kr彯��b�����?�W@��m��Fp��2�<d.�"��%C�~Ut�s�A�2d�F�.`S-�	�?@��7��&�nm:yO*�-�8X l޽<u�s=]�f�l�8��\ˌ�g8��Ѻu���|v�{p��+�e�v�z��';C�K�hj� ���F�J)�d���(�/E��>V�"��UTin�Ǐxa��hkQ^O�ٗ�@����ٗ�FH�x��i)���ش��$��ֲ�������}������7��� S��x���рL��8o{Q+��/+�ܮ�v��a�-^CU1Q6���<+3�+�t3Ŧ?~�������;Qw3�Z�D��ۇY3�� 7p�U�����������j��:�A��J\.��u��tV��<��(x)L��T9�m޸�כ^�7��-�8jl��9���a��.�������ݴ��S��R����v�!(13}�x/S7y��E�8X�8�?�O�w��/�Xz�Z�m�懀C��"��]s�.�_��:� P�
�j=��6
�� MqJ��:���a���OH��G��-+xޜE�*X�6_���p�
��"p����� �-��ac`�`#��?��8�ܘ0������PqT�����0�u����Ğnv�7����Fvfp���e����t��pP:�uE(L��c����)ۂ�W���r�
�֥-�!����������gz�/�iJ�t��&�aHաfD�m���%)3���Z����ٜ�m���e���S?�K���2�d!��y���K�rr��/��:@��z�X?|�-Lٺ�0��v�`�y��S#-��T��g�Go[�r���@6CSАv�U�P������Sd%�O���L��	1P���dDsRr�����6D`��+��j���DS��WC�)vss�|%t�p�F�J�>�����+U����M��ll����7�Q�
��r]$>E�^��S�����E�Ӊs���7?�ӄ��Z ��^���>*Nѣ�?#g/Z�x��/y]}Xe�D��6z�gs�j��Ͼ�/��m��D�TNX�=0ކu�NNS��6+i_Ŭ�Bh�)[��V!�<k��&���"GC���D�"�Z�����������WC�KR�LXB>�7XKa~M_�K�㦪����@s)��2��ub�ozt����'�)4���˘ꛏ �M;�;P�N��'>��"_��;#�M�5�0q�8�g/(�M�:G��
^*
G�bȔҪ�|nF�����&x79[@��sq�lʒ1l�H7���e6d}5A��*�N�'4�Unw�6�M.�ݠ�����J�
�Ta��?�8����S�o����"+� ~�uZe��OYL���mu��5m����4�s�qR�fV����(��?�O 7޷k6��t�������ޠژ�<��:����~��z[����)�?z�r��1U���B����:�n��:=|G��ߨ-�=��}�M�������#K��؊�t�����E�z�G�f��"����+0Anw����:�d۫�!�Y��G�9��+��v��/N�.|�6]e)9��Vmm���$5����1ޚ~���0p�(�"b��c��BQ�[�-�.z��߄�;�O����+���p�a��|��Í~y�����F{.^*F����3����w��h�d�/����г�c .�Q�&��Ŧf���M�gt���F�D��W����j59\@���&��M�6�s�@]@�U��m��ss��P#��Z���6;����R���)��X�f�P�շ�-N,}�vz��6>YJD��L��M�y��:����㤇k��m=˯&WP?L��b\0��3� �W�
����휦�O9����5~�Ey�_�M�~��z��͍s�ٻ��0>Dׇ�~�lT.u�+�ƿەBj�2&�Zh�j�^Ò��;�,����%
M9%���{x�9x���3�u���Շe�c��?r�Z �`p�Ip�kp�~�Hs1�ş��3W����W���߅�� u�9�
M���+@�ʊ]�@-�P�>��K>n��1Y��4�51�SLU����(��Np$������X����1M��En]ˇ��i�S&�� ��u�S���b9߅O>_���*w�<m-��:�'�\~E_���R�k��G� %y{��)��Y?n�g��~��O�< e��F�a�|\h;�v-ɤ5��\�Xg<��pi����{1����%����x�_���*}��:�qK(&������2'{e�R����~ee�M�T���,�q�jj(����M�خ���s��z�v_I�<�r�X��W�)9=M��(����w���"4
M�����:�E��i��������f�δ�/��0�����.��b����A����5Y��7q�l��l�j4[�1n���=�B��5Pr9��nO>�!鸁�x�_y���G���1���d4d,�3�h1�;��~ꋨ޾�%T3Q�Ħȼ>�U�%�W�u�y�چ-�t�~/ڴl�#A6h�X���[�P��ç�аՕ��.���*��Xs�3��O��\��r�p��4Uu^�������dy����B�M�M�'���^]ͦC�����9�h��֯Sr�§�j���^͒M�?����s���13����"FH�(��-J-|=<���؊ׄ����ZY�LV�����D !��"�d{.�?R���輋!�H*"i>�߁T��/v�[H驨�$I�����`����gp�ݻ����@�B���&���r���	+uJ���G]�8�o.����R�.9�����U��7�ܮg����N�p]���<T>̓�b��rdڗD+�*�iu����Z��ѕ;�Fhf��b�wu��(��S�ʛ�#�D�~��#��tU�m[gW�^9���!�Wc�:�����s�N�rw�*�(E�J�=��P���U��.c*:;K�v�RةĂG���k� �Á����IH�e����{�-�=^8����
�@�s_˟�n'k�Ay�����G�����}�g����L���=��ꄕ�~l��:˫o�h=��1�f�˓ N���a�z�ì5����*�H�̽��7$�2������Pr�ũo�e_X�u�J��X���PSܟ	�(np�l��Ottb�M�98������֐Z���@{8��^57��,��������nU�R1O�)�����n'#�	���Q�b	ƶ�z�#�*jY<{3f�6���V�9�wRV/B�_Jn�77.�]N�5�Y�m�a`�լ���}4�(ؘ�yA,����A�7_߃VC�¡��}���,����,��-��I��2"�?�8�����3��CNNyJ�Oݶ��\[b9�����B�Ζ�����Fζb�
�4;������-�Ҵ���������-����IH|�����Vb��./�#T��mzJ+��:���f_��W����:Z��đ�$'����[�^�"��vq���-|��J�I�g����%��'��9r�v��[�u�VMF{xݢ]�����H�ň�K�{��\���$5���~v
s��eH�+����f���7�8َ�����59�ǼT U��GC6n��%�Qϒ̮i�B�v��r�~�q���a��Z3���A�w�Dt�l�7ަ��m��\BHH���`8~_��ֱ�n\�b0-�5	\H��h]��9�B+̊��)x�I�>�s�L�: ���&�k�V{9*X��WY0��֎��E�v���@�M7�QZ�~ko��,`�'��a;��0f� Q��?��Ns�[��^R#���4�t�|�u�N��B�{�L�>����ؘޯ��w7�
��TgG�Xh����'t<�#�_+0=WdL��D�o����W�{��Tx,�H�T솰����"[���>P5��-(��}���︍�g����fd��/���	q4-��o�؆�J�Z�hJd稊=t����N���r��֛RwQT�y���L?���/�_۰JF��� �{}3$��o�����q���Zu&~��y��*�#Vء���/����Ymoh|�)�a����(��F�@�}��Y�K��4�V���at̸�ۯ����V��V�O�Ğ1�Yeq������`�A��Iw��K��68YL' ��Y�Ĩ��7�D@�ыj܅�����e��?���a��M��-2sD��c.�x*S܄�m��tk_)�OLΛ_��Խ��RA͠�&�;/��Rg;�,5�7�t�@������0���_x�O'�S�����i	!����s��g�r�d�
i����_����<ק�E���;�.֖i.]�M��[NBh�_�Ӟ���!7/;�ꕄ҃?��ا���1M�+��dP���Efr�u;/�+o�s��[o�wM��;�ƣ��t]r5�#%���7���&ڂ��n�c`�º:����\`�?�2�7� (�.����F`׏�йU9$=/ؘ>�WO�50l��۵+ ��S������+(�n�9�,}]�-�!Ӧ�c�,�B;1�`yR"�
7��1ϞH��O�M�ݵIĩ�7�� ���,�A��7n��tN��y{��΀J��Zo#؟֭�}t
�E���ePS4ک�hX�+f�#;e�������VO?tϵ����1�p�}+�D>�=�T�)}���h�[}6g���o�_�lJk,5?q;��jC�껷��8���|���M��]�ɣ��;��-��]��I���x�!�,���f��yѭ��6U2�Y�>��oED�NϑM�0/Juܮ%]����2����j�djCY:���-���*��o����R��� bD��:y��՛.A'14���R�ܠ՚���uw1�Zr�����B��FS�~m����x�Ӄ���%�6�щ;6����\]ÐsN,�C����6O��g�4�ewcPǜ�걜���KRd���3��n�Qf	���V8��9xm����ӧ�8��T�����D�%�?��c�b+1��;��P�+�ݴ7�B����1��۫*�p�N)�v6���;��1��DgYC�tr��|?�:7y{�|��Z�#�	g!4�]dm�J+n0yڏ�[�IG&��ͤ��{kC<2�mk_n����0D�$?k@�jUMM�e����"�Eӏ%O�r�0�ޮ���-�Ŗ.�{,���'�DBK��+Y�Mɴ�B븄���ȹ���<MXȟz������(E���	��B�S1"�lO��w��*��(�� �"wOnK��l<�B��͑uZ�h,�ct9ѽ0E��7�`����i'�i_���][(��dp�o`ͼH�~��
B��@BA��� �O�sv�Y$,���'mF�������H��A�>�w�=��q�&���.���a���g�����l��v�E�z֚�x�k�;PA�vފ��T��ԟb����ߝ�$���$�����<4��-�#��2��ql�����Hm��6�eN�f����7���^��gu�ID��R���gӹ67�b�Z��Wq�����壆�q����S��O����|�õi�BV��v�3���Sw桄����|���S���3#q��Z��?g�;jk�>d.�4 �e��i\ $�>CJ����z����r(�����lq�d��q���Ŷ��Kr;ĺ��=!y�l���fX?;���R{b��p6cm�0��m�۬�mp�=�|FX�6��4�3�Z�
O�=�=�性��O��6j07�cm*��p���`��������
|�	�;Q��b��aI�̧�
�����x���ʸ��ckDO6~F2����u+6,����5�R���b>��G�߬yy�5�v�4&���APb;��c�;y8h��e6�L���Þ:����=9
N�q���Y�*���q{\,�#�b|��z,c�7��3�$��n���TE��'�du���Jl,w5,�:��Edy?�B �|�O��b\n�qnPb�PZ���\��}���v����93��#��?3P*b��i�R��Mkj�^O�1�@�}�Jiq�+��Qh�j%"�|�S0�~��en|��]�.T@Q>��*������7�׬ľ��x�׍9�KDE9w�E)��V�}}��'����e�׊��3b���w�U���p��p	T�x�8<�����2cBX��S`���x�sT�^������+�9����r>�<�*��u_P�	lk��n"��Fa�Mzo���r4;i�(�u�-�n��F�"��f��[�w�!nQڣ?I�x��?����>��{y��u���Z��:�A�C�ڹ|�?+Z!bw[G����t�LwIWG`E��k/�?��!��X�E�7�^ ���.l�#~Ͼ=���C�]��yV��x�0Y����e�|'k1	�n��U�N^����unk��x�j:���nW�[�y�!�\��۾�N���=���5tS���u�$ÿ�����Kt�E���P^^���JK5s_1.�N�]P�#���\��Ɖ����V6�XZZ��	 &���_�����e||�!Ce+������3N��0��T-�n��Da�V���0�o���	�I;^��T�T�@�y��ł}��T*�Ϧ{H�"� ��%R�c��%�#<��Q-����ؙ��놤<3�5_M���6��N�T�	tsS��W� %l�r7�N<�^H�hn�r�6/�\����HC�!��/%�S	N�kjYL������w�&�N�I{|�fЇ�٨P;<mG5;�s�y�Ch�_)0�M�m��lۅ=�=����)�G�{d�=5�&q�o�|�fq�:P8q�׫RqhH3���\�/���+�KE��-BM�6\��<�_�d\��InP��t�ګ�+gF�1�,��ڻ�-/δ�roN n��G� -a���2�0�wvH���sCY��v��f��g���Y���L[Fؿ�����ڀz��+�đ��Ao��8+@g�x�)΁Uz�	���軻�eO����G�K���4��<}z�:�3��v�6���OY����*?�W{��~�lc��ďt���C�V]\�o?�Rm+&�r�:�s\Q���9!IB��+;��}���9�{IFe��V�a�dA� ="�}�q���9�`������Ȇ�0w�?����8������@��@;JL[�-�EA^�����^Ǔ���ot�ل����<:����J{�'+��?R�_�S;ˢ�p%�m���)JH�8�˚6r�S����BpY�t1D�_x�s��#��w�<�6��DĖ�ەW�Ȫ�&ݫ�"K���_�`���gIxMoV��j�E���k������~=�@8Paz
���|���֪:^6�[{D�?���Z�Hc���;�t}.'���'w4F��큁���Nm~5�>��,~^Yd�͌�JK�V	�X�"	ē�ܭM�m>��(���k�[ᛷ?�Ɏ������D���0� l���y��?%��W�3�4��<������g���7�$y��<�F �\Oj<�?iP,.ږ)��?����x��HIˈ�����?����
�M�n��-����Ňz�.��W�.F��f�4w� ,2Sg�H��-�}�l�զ��I�4�8R|bX����W_��[�
�:BɷbbF�w\��v�V�����3�VbW�K
-\;`v�e���>6x�B֔t`�
����(R��#j!w��2��u�s��uj}5֮�?/!��C�h��E�MRe�b�
j(J����fJ
MaWte�.��2�+T�4�1gK���8�~o�Q���x�l�<C��D��b������j-z:!����\�pj���@��T\Du�T�]x.4"��\��$��A׶Q^8��e;U[��y�6Bw�S� �v<n.xc����LD��8�?��N��I�q`��T�W�O'ӆ�guPe�,6��G� ��?�˘	C@dp;H*���0�`��Ҹ�2�j�ؚ�dZ_R�r+Q�|�)O�f��qХ�!CL�&���ytZB�@�5��[�}���Ӳ�Oxc�H�)�*� <�1ɯCeAd�Q�s�V4J�P��%	�m��Z̉�6�ƼI��kT)�3n'����a�D"X*�i�I1IƓ�|1�m�!��>�u-3��������(���aY�c,�.��D������9��Wן���҄�I���ф)z��"�Ŏ���C�]��5�1�X2������K:�3H}��D�N�L�Z��T��uM�?�� �B��y�4Q>��T�N����L?��,[�nD<M��ï��5���&�_x�`��Н��菇��*ZوQ��w�����u�k����}�_��$��ŏ%�S�w5�R4RpV�u�){+w��a�X�P��0lZ���B/b~��%����f��߹��9tv�򌲼����ؠJ�F�p��!��Q�� ���i�'�K��d������3~���_���3����������%/�W}�R�����ׁ͝m����W聈H�4�-�O��J�����z��z~kvE,���%x�Uʨj=*�ש�7�0�����ްx���3/GY�ߕ���~��P-�g^#��'[x�B���l9B��Y|������v��A�.� ���BPA�$$�m�t���Q�K��M��4��wޑ��H�)=!;��=x�z��"m�p�@b��}d�ß�Ɂ�<J�[�m�f����恗G�愘˾�W�o�@���Z��$	��(߲I[�E4s�6�x��{S^���`�p.��V`������NNi=c�J���w�.�F��������]z���İ��<^P��`�����y���y��j�l5�����5�	/Oq^��?���
��tWA�C�ه{�b�J׿4?�I���/��̳�=���|(0+��'>q���P���/3��:�T ���|�Yt&C�Q���Jl�#����˭Ɋ�HovnIb?�KYv��n�����Po�Mᱳ�q����v)n�����H3��^���h��EB�M@̄�oN�d��Rq�aA��ڝ��|�N���U`)�$(V��Xb&�faL/���.!%�GbD#��8Fu�����@W)�,n���Q+N�/r��&�a�:�iQn��������'M$z��C+'!��p"�n��w�]H��R%h�cE�o�9���%S�E��/6�-�S�a��G���d�k EX�����0��7�T�/ʢ�(��{FNCקe��a���XzW"�u�[����;��#;oa�W	#��[�S[ۂ��:-�R ��;-"tc�bQ'����9��O��.l 9p`��Wn:(����2t� �<����z�oD�I�ס����sO���ߡ��{��x
u�m'q���l�q��;)��]�E;U��я�w���oŌ������p{�m��L&����I.XϷ5wa�o(����vfde���"����ȑM�n��K[����E@�{��1�cعQB>���_���b��nlЎ�ܵi��s�I�4��>?Yk��ķ�9hr�'�������n�eyi��ӋG@Y���a���@U�{v�P��om�r�]s����-���*�H�ڳ=���I)Q��ܵ';C+ϱ��.��rO+X-�dF�IL�8�}�_{e�3��]f���D[/n]G���WȰPF� �h�t*��K���;�f�%��p��SO�ۊ��w�Ӌ�r2x��g��rs�Ko+�w��\]�\LZ2��9��������OX�	����%BX9 &�R11���]t@�?:�.�G��ب��k�SS��ӻyʉ���<�@� �����p ~ی���M����I&7r�\�}0���d���_S+>�� �2%D6��h1_��P��f�]�T��!�[S_Ac����Q�~�ջw����Ta�1��0�c�[y�?9&z�1o+��c3&o��^4yN��zZ�ϣ����^{b~�������ҳ�J/	��{��~A�k�2߱�z�!K�6����?�Q ��~���V��%'h
{�h�����b�i�tg��w��T��Ŗw�XĄ7�Y� �+h����9���WSG)����`u~�	r�f��}�m�t�.���<��I��̦�am��H�7C�Bn��)�V�5"�������ί��ҐB��М����u���W��zQ�t�k�X������m����ѷso��y<��S�}��q�b��s�N�D�Ab�r��@�5c�2�9BP�(�P8RF��]ý��-��b�a{mN+�N��b����)c��q��s��ّ=�9�����ӟN��l�)�k6�"��m��h�W;h�I d����s^�X��_З�ݢlӫ�J��+m6�tU�>B�p{y�4�MG{�+b髠���~M;��YiXմB�a�=h��f�P�"����Ǉ�o��)8�ڗ��y��	H�xy~�sO��/;�Hm���9*Z8]y��Ъ^�U�Lu����;���g�a+YM����4#y�w��|����l��D���0�ظ�/�dh�L;��1�Ջb�@�D�՗1���50��1��)�5��b�)��z�cZ�nA_�_@����GG�׻�x��+3�Kz���Lێŭ����K�ץ{8|����E��lp�ETvj���v��V��愼�L-�9���snF�a�k����i7&�������7�ڷ9�	�N��B�η�?\��=�&Ȫ����?b�e��ǆ��;Zg ����y��@��
h��|ļ	��o/ꪝ�'p��ΏX���D��R"��j�A��ō;��_���?��LRΔ��k�����N��V��P��1�Lۊ���ڐ��Εv��O�V��Nx�*3�)\��m��,=�1W���<�.b�J	�lP����(���4��k��dڴN����߶=�u�i[� o�0ܱ@�P�r>�;��TS-F6Ϫ��Q�[��
���rQ�����9o���Ha���A\B�-�/���S������(�� ��f.��hǕ��!�Ӎ�O�#��b$K1nնb�{1�y��xn��r3'�j8�Q�J�q��	�\<�o$����#��+cy�i��C^��W��預BA�fϷgŧ���1a9o7]e������	s����PK�Piʿ�>ˡl��<�r����cq�K_V87Sc�\��&��`�Wtվ����$���o�D�N���d�Qr��Y���)3"�ͽv3��1�* �
~@wG>�lQ��։ �	�FO��K��,�i󺬕h��(S��U<�K�!;�⻻��z�/.@ם��N>���m�ϱ�h���0~@{�V�.��)5�c�����VyT�u�K��e�����9�/��	q�����G�k,K�8�:�Ĵ��i�Kgͭ�<̯k�4;�(��aqw`É����a���n�b-W�3�4�-0�7#�Y��I���M+XX�?+�u��T�G[~	j��x�j��K��4���<�$�=�bܘ<���σ�y�T�̹��[Ea���9��=�3�0#���R�G���v-}x��݅𠦦�� ��o�l'�4���p���E\To�ƺ��Tm���(�S훿�2]�Rv��p��̞?�JWg��E����	Kxϗ��[����["\X(v�k�vc�@o����F�<�?G�+|���Z]
ad�a���:j�.��|\��O�[��0}�P�;i��0�v��H�A�Y�C�*L�*��&{NP��]���,Tj��8�Q�3П�x���?��ʠ}�ű�������Þ�!Jgh���{�ll�{{b�4k���u<ܔt�3��J�<=�.���F+w�+45m�!A�|tvv�#!�����P�dO���$Oj^�w���!���Z���o�qO��Y�"�ȏ�ZSۜ��t�n���Q�W�ڔ;x������z��;/8?�4��\:��[X��Ż�3�i�EA��n�:%���Ng��_	?1�۟\5�Hb=�	ir�Ι���p"W��̉��gHc8�����Op8���D��$��cH�(�CkXl�퇺~f��=�VsȐ�;-h�As� b�DZ����M�Ϭ���P�5y�H�#ӏ���8 �(��괘�teZ���^HO
}���.�Մ:��3c��K��G���{�6�8�ǻ�9!���ɥ�� �+����"��Ǚ �OO�V��=�G��Sl��"��oj��-�_�{c(���Q�U݈y�zu�	yf�SS��/ZHʧ;�8x�T�G-\��0H^S"�I�������eE�Md���٫�t��|�*5��.(䐪�I�vy�@ep�<�}�8��ʊ��U�[߉Tय़n�K�1<�[>�&����/�.�9��
�;��l��ݱ��k�;�
���*���>������J#EI&8bc��p!�Z���F�;r��g���on��Ŝ�X�2gw�]B��b�����M�M�2OE�Ս��g)�m��2��	+��@n�ȱZ�7���3�zC��b��d3i�O���f���b�NG�I`�w<̫���d��ښ�"T��������S�Ǯ,�N�VR�
��' �{)���/��6N���g����4L��и��)��c������~����y����t|EsZ��e�e��ؒ��>�1��1��3�#�'���߹�t��Kh��P�2��p@f'���i)Ἂ�b15��V��o�N��5T�y�1���U;�.�N�����ꕩ�O2K_��`�`2�3+�����RmG3 }����� Oh��" ���'�xJM�CY�<�V<��p��Ao��	� N��9_Ž�z�~��n�� �q����R��B݅�#���$�	nr�q��5���4Km�{Mb$�УSj|�㠭:��Ƥԗ�V����o�*�d�q[�N���S<x��b�ݪ}k`C��f]F��Rz�W�l���@ T7�$�����X1�U9���V���I��z�3:M���os�ͱ�}OZ?T�3ո~A�'ΰF����dc�}�j�S�V�HA��q�`��3D�a�f��cJ��F]з�`C�̚�p�`�9��fc56ûD����,~��8�zG�����������`1�We������8��յi��R��Xy�(��G���)^P8g�Hu��N`Hl����1n�BZ��W��r�q��O:�҃�\�dcײ���Z�*��1%/v11�C��w���L"m���H\[,-����s����mV���uX�EqnGy3�C��^��Uhoa�4���>q���a�ƋL�i��Jh��"�#[�^���h��U�X��k�;ͤp"�7|ĳV�W��c=g5�͞-P�e,��DKY�#o�u0��\�j0H�V$R�U�˥���F�q�b������Я@�++'F�j<Yz�&_����8q��H���tӸ�e g�~���
���m�4-p �DY�pIJH?�v-{��I��v�7p��:��ʀ3�.���㼥���i/.�vzK,���;9(	;�m� P�����p�\j�|p�"��,�&�y��+���y�j�ݶ��N6����	�}�WmC	�)� W:�>fF�8���f&�Nk�K�`M[�:�*��'U�<V{�����	T�Ĉ!ݚ���ӂG��5�L�lX�u�^��.����nD20�fy��}�j{��5C��![�K��ngӵB������]���]��K�����28�Npwgo��{�~v��j��vQ���=}��\�:�=��Ԯ��\��������spܖބ�����UDa�p�-�j3��Cq
�4tKq�|��q�b�h��s����H��e��Zs9�K^����5�)����]fu�{.�E��ڗ���b�ߓ�vS��	)�� .q�^m���l�����)��U�'h�0�zuF��X��+J[��}g����q�a^q9�4��;���n�f�YK����AS�fxU)��T�P�Ƒ[�b7a%�\O��Na���Guh�7���(���ڹԾ�E�v���Q���h����g5���|$��8��Q���e�fBV�\����D\��m<�X��sB��@�4��w�ҕ���J']Hd}� aܛ���~��m3�������ۉ	Q��293#[�5��F�5/�jI�M�PQ�,�.�U��rω��K�+_s�����ua�N�k;�q͵4�w]@�������6�.���T���UU�XMrY��3X��^�3���~��@��j7�o�~s�o�}��?:*wx՚#�(�~��78y7��AҬ@����r�K��uc�Z���p}r����_����&�=7�-Sa�H� ^�T�{9�J��}�*�*4,����"J��}���I#gۓθz2�g+�f�9��h��1k6�����'��,O�Mv�hX�?ǸL��=���#���P۫�V����5*��5G�_j��ۻ��E�������">i/������@�j6ԍۯ�����b�ԉ]Q�����Zi���Ra �kmm]��hSL���{#ܳ�H�O�dǕ��hq-�U���R.��r0��̝�y)����u>B��ȗ�e4=�L��ٝT>��!oN��Q�fE<�f��Ѯc�U�,��˜�Xh�{�G�-���}t)e��M���w\���-�>e�y�iwWj%�.p�%ٖ,�����li�=SyY�G�ML#�h0vv&D�N�էol�KN ��rX Dsw���2�I����կ��+�9߂P:gE��1���<���zm8�A?f�\��m��+R+��i��k?���A�3�Y�qF�ڶz�X磊M�C}��H
�3���%��ys2w�e�L�Z�5�*�z�)��������g�8�
 =\�'&̊�L/[��B���Z�R��i��3�_l`?�l8OWR����I���KĘd�=��N7�TE]qd�����iFU����K��iko��撤9����I�G��w��?�d�Yu���v�i��ģ�J����i������qƁ���Y^�~>0Y�gM�$3;��CKg���~�@�n}#�:n̺�ߺ�GN<���_/e|�L^$T�̠_�1'x���;g%-m{C�Mꯋ;E,]l���h��;�vԾ��r���Po�q�7���~�dd˚���� Sо��~{��]�\��2c;*S�\m�^;	�@q���9'�蓬�&M�5��yO��u���n�7A��� ���8�����J��K��-\�¸}�(|2J}��a���pI�vb###�̩�+1��=��F5�c��t%D���BL�d�U���U\hOF���x�_�ԘK����Ko�E:�����Kf}�}UɹWq1)ofJ̷�1���:����[߻�[>?|}���e�%G#�m���<�A*�K��� ۷�N&�7��+��j�򲓿�-3�v��k_H߶z��gdj5���LQvy��W����gA���oV�s6b�餇n��	�og
:U��-z���7?�� GYM��tKF���C��A��
⾥�y��f	�
D��t���\X�R�<�)��1����#"-ۅug�*�����8N�o��"��ˈ� qu	e��wԫ15��J������^�$娽ߦ�KV���Q�D��p)�!a4��e�R!��
i�0�����������UR�O^�߽(��)��M!��P��p���o�0��}��,r�>^���~6aEr��F�����$.��˩!�#"#���<{�#�V{5����O�e	��{�R���r�2�ҥO�x`�ҍ��G˶��1��^uB���A�n�"���U�5g���: H�b��/?����0X��u"���nO�+0g��9�;y�xQ�]��*�����F����z|��	��=�pѿ��
'�����_���AAÆ�/4�=TA��~'0$�I�ͳ`\��y� u���9[���~�(�1R�)<�@�1-�=�]���T�����G�J���֖a�O/0&����Z�/N�s�#��斟eZ��u��/�Y?�`�9�������}]���""��^����c��3�*�{.�#J/,h\�1O(}0���Ua�6�#f"��Їn���䨢�dd���'9� �8=� �|��I|纚����Ǝ������, 6L(��rP�M��M��}\����oA�#�sH��C��#_��9U�w���P̳kt�>PF��]�L�ݎ2n�23��"bO���ǃD@0��픗������4�F���'��2؛g�]'�����ۖ�/ߺ�q�ʂ*F���Ja[T3�9�"0�'0Mlw�TX���uY�	�OE�����>J{+ɽ
�z�\en�0ȟ}���{����H����f��]�0�u����7���Aۈ3���5�.C�E��/(�j7�F�i������;P]{��allP_��Z�O�+�l���_�ڲ�.���[�t�=6g69J�P�Ǣ�&�
�1�UV��(;�ڟ����w��S���Y��:?�w����5<�/���OJ1De��;�,�{L/�+���O�E�v�d��jGڱ�gF�û��HK��T޺�퉥�#�O�S�b����0�$�G��<B��u]D`�'�W��U����R���|_�B#�Y�)��c=����˦��fW*��
R��&���Ĵ
U���g��B� �����q��A���M�@HVk�����}
�-�l�˲�Hv9J��V{���$�;�B�~!XU�NUx�Y �y�U<%Tfdb��d����$c�6��)�:�����$�t������[D��mȯ������px.	��wD�\rc�a,t}�{ނ&м~�И��R�s`�rZ(�������6Ik�li��'@3(^�C���@kq�9�Z���`J�".�5�t���p�8�~W��pp��f�z.�%�_���ǚL�>G�?������Ӿ�1S�J�h2HP�I���\������Q�K�t��,*a\��4ϩ��6�6߼�;x�z���~���@��}�{�a=�Zm���:�t�Az���hh:�fk�K�x^_�崰 ������rmJ���&V��wYŘ�v?`3>��6ip�(���Y/k��C̻:���!~۟����֏�n�ĕ��&�ҟTqe�K:q�i}s���|	��������1Z.�\D;_��~����l��i9�^N�k�:3��)}L+J]i}y�?!K��1t�Xj���^�:	p��w,\��pF�X>[�s��*�������p�2ߝc�=�H^�z�x"��6�ou��׳`��[�%g1�
?@k��Z��{<,���?�����ު�K/R
���)i������_�D���7^�(�����x͋]Y�f|���?���=M%�
�Κߢ�|�$j��4�l���:�cFĸH>2쮋����CÌs���E[N��^�f #�����H�=�E��rk#�P��BWD���o&��	�=5��t�?�h<m�:�0򮇂O��rum6=8��H��6E:e���#,=C84�Z�N0�ʁ�J`�E_�H��HVL�I嶴�mg���n�2I�5��C�cq���T��u����^���GǤ�Q�r�����l��(���)�:�B�����wp_?rd��i�$��y�^I��������T��4�wk����su���d���$�|�߰�(��:n�>4����v���|i2��Y�E��\^��`~��H m=��<s�~,#.Y:r��������%���Z4�_��=��:��'�co��{����[���#Y�v'٬�9z��L(�W'6�DagW����!��Z�P����_�N£���.�`�tF�ԠJ;6�?�6T�2s��J��-<�2��pQ�<� �z����ٻz�ڻ���d�rF�⺓���(�U��gf�R5,ŕ���Y2xs?�_�H�^�Sr���`�AO>OB�(z{'�N�����A6.��w��K�.���������s�*q���O�5�$8���̿/@�s��~�}�5i�#�(nIH�U��;):8��m���Eba�t�i�G�l�����QGZ�lK�TI��Uoŷʯ�9
R#+56dYĳ�Re��7���x�3�wN���W;��<|�*��e��=vg��@Rjj䭇�y�;t˔e;�Rg�T�^E�֋C������z�%c$Me�D@��WU%\��Y>j5�	`q��33�B��s� M_�~<�\,�R�RZ���&ʴ��s��zV�ò�3ulL�F����]�%A��Z�UT�#)�-_�/ȵ([��S�p�ۿ):�Q�'���8Pd��lnΠ�b��:q�ϊ�+׷�Z�m�`��V \��y�8��v�x���f��U[�-?i5�|�Ǐ��+Ѻ��3��Jvk܇](w�F�j�*�m��u��qӴޤ�����kK̪��5�u`����Mͅ�gց�c�;�
ϱ9n���)�0��q���m�H3�z�
�,8�kipE��g�� ~ܛ5(O����`�m��Ȍ���Z^ ~�Ҋ�48��o��a4C|`mi3�q;	����zΰ�y���{�n��@M�Vi)�~�E0v����������H�Q5�N�_�� 4�N�M�e@0ߡ"��;�����>�<��P#6b3�cc� ��4�>�ޗnkh-5ȳ롇�%(�0������|;BY��g�S+p��llo̎�Tk#��;}6����s������\G4�x�,��1�_yҦS4+Pۘ��JgPr5�4ϛԞ��zxt���"��E��>��y�uDY<��:�����Y#N49!ķv�>
�&O��'fL��)��S |�[�V#z������uׅ�%n��|w	I,L�Ծb^��T�7`��h�N�1�a��[ �0�O���:J���o�t��Y�:������#��7֏ŭ�Vp(S �م �0�"��p�4H�DbKGu�:�l�%5OYW+�c>4y�3I��aC���f�ue���l�oGp�9�(��
��������S6��$!��Q�7������+�L�r׀����"^�E�2�گ��~����Y��fi5������ȶ���%�ft;RΥ�9x�wy��s���t����"�9F��6�z�@%����KӲ�C#���_�މ=�;�u��M���;LD��_/#�=I�����8�?�h�@6���~����{򈥵M?CM�����ǐ�6�-h��/Zx��xL�-��p��a���☃�B��� ��xd9�Y�x���E4o "��9H�'�K*mZ���*��o�ʱN^gi2ƌ��M3��.W��+-�$�lX�n3/	I��ʟ�T�����岹洠����Cu��j݅��d�p�Ǒ��2����d3�=��p3�j�^KsA�����RQ�k����;�=:���T������u�-7[�Pc5wm�z���&��>������?�9ŹPt�\���0#����I��Z���6�q�fh����׻��ȋ�k1�y,m"�K=�N᱃�͛<*JdS���s�� Vh�C�OQ�CP�l�c��xz�.R�kPQ�r1�)����jn=uD:W)\@��7ۼ$�̏?	�@Q��c������צ��?=�����nV���˨%bP�6@>�&�VN�5��6�{O�;$�����f�Dcv����L)���.*�LAdtν��8T;�D����V@�0o��P&�/q�b�#fT�tg��!��� ��6���]s�g[�3H�9�9�3B�K�����_@���m0��B4��v����w�o��p]<�9�MҌ�5Cz2Ӏ��`�ᒮ �b�j��]�|�B���i�x�a�v�Kq�d��rxg�Fn[S��Yd�I��Iz�����UN��C9����}?T�w�9��(O����D\��4�|?[�Fp�İ��9��P��G���b���urD���Sg*j͙\�1��*��\�#�0�#`�[��
�����'�7eK�f��:^��޴q�MuA�\4 Ml�i��Ϸ��b�#'�Ϛ���L����/�8� 2z��V�K0��Fr���j�u�&�w=���	�7��-����Q���mo��5|�u�M�\ϢX�c�O������p�D�0[ew�{y_"������yG��~�U��*�ˍI7<9�H���$��r�Z�#��!=L��S��h�}����~���z�����FAJ�:�?|P�>��ױg��5{�	�{�4��0�\7���ġZ���Ձ�c�V�N��;�;*�b6��c��
�~����;p8I�<�z�sǈ��֒�Y������P��`��ė��-�9���g�8St3��ٛ�����QfY��0�b=䧥�Rն&���[��};� ��|g�K?���4��)W�ɔQ_#�֌��bHr� �lf\�T�0a�[��T3��k-��[@m-��Pb�ȻC��_���*V)�!(	���໗������v�5����Ǜ��R���NWD	�}�8b�TS>�1 ��~���@�i쵀�1ICd�U��Z���,�Z�T્z����.T�n�Q�w1�1�6�l���>�A�M +��v�]*-:�����!��ૡ�[�cw��ϐa�e�c����n�'�<E�� ��h�����/�������'1��`L�Pl(�c��V�K+E������N�,��޺,➳�\J=Ag����ZW�[Qt����@mх���r� A�K�?P�,�ձ<��5�U�is��"�,1q��$n����{��D�o�e�V�� F�#/ӳq���.^:�(�Z�A�ξ����Z���9�J�쵦�;*A$����6�tJH6�O�l�lp�~j���;�?�7���UM���=�ܖ��Y*�>�3
���d}X�\�v����~�<p*_\̏ BvB��?	�;�w���J��l�*iS!�
��\'�OR`�����HXC�v�U�mk/ٵ���E$�Y&���^�=�h.>�P�,9�St�אcψ�)-oz]\#'�1I�WQy9��k���Tt�UXd����ZԪ"8�XZNN��{�M9i�.L�/�/핪gU��B�#���naR��|<�\� �@B�Aק�n��~�E�E9"�$Uw▸���ؘj��7U�L�6��T�Q�nV��*��1�,C�s�/G��1@�,M͘sn��Ei�q0@"��ә4�;S�X7��3�߯�坱p�Qg�3�. {�Vw��!z��A����Z���x�l�j����F�3���	I�=l�Ǟ0z3���#I;��r������[�U^|���7MY���I#i��ᚼ(f=n3�%�IN��L�5�>'���g���-+$ �y�,t� {dȢY�˫�z��VD� 7�U�Ln$&�t���ﾈR���K
�CA
�Y�qa�)E7J�&�L/�ً�q��gtd�A#�h|�\7<ᾣ��� �iƠ�����=n�����J]��9#�=<"��z�ٓ�ӛ}�5`�#eL6������%�Pm�J-��9� �H#�<�%�`��M1��Kb�|;뮐�T/b�?��&�A�,e�� �o!si�&�z�RΊ?U��4A�٥�*Y%�c��� ^e��]���N^��Ԡ7�wAh��I[�¢�6�'#������c <�����p�����\#�-�667Y�~���r�_�^~�4pϖm���rd�,,�y���$\�><p�4p�"d�[��r4�3j���Cn���旰�蕨���a�=ζzc>Z��i`�4������ݓ�P_��@kAj���d��gG�����geU��tf#��Mc��擳�;Z�Ǒی���/� �U��06))���38=�]��dl��vğ��%�'圡�\��b��-����Z-i�Z'L1R�{x����ߎ�f1[��~qk&9Z<wIj]OE �Bg�ڸ�;5��T�VT����8�������#�Udo��Ey%��������T�(
'�%�~��E��{�Aa�f�e��HLG�q�azG���6�y����X]~;�_�� �n�J�*
Sb��z�^>&'7��cߜPꓬ�b�@������e@L�6�'[�k�iVu]��䶔��Ff
	Y>N`w���47�[��!����<2�������otM���;>��������x���Y]�G�s��E�9�P6�(U�$@�A?�C�4��@�<���n򷯇�@جo������I�N�6�[|7����wD%x�#�ͯ���5��؜fl{�8Q��2��v���m��w@������(KJ��LS4�R`���xD�m�JK�Ap�̼�L��O*�)Ԉ�����B�4�����cC=-�N����/I�>��P�[V/�WHboƫ��ר�k��5��_�ȹJ��Qxá�82�PZ���૩u�� n󍰥5{�/k�D�Z}y/.�"�0�4#�!~��m+=�A���ՙ�*��4|o���pΩ&�D4p�(��K�`�C��̣~��u�Kc#��ha"�b�i��am��9�(�M��u�Jm��������^͉��A��P k��o��>�*�i��z��@m�%�5/n����>rP%`O��94~?�����0�Q��R5��w�Y4�:>o����\��?�'X3��2�y�Bz�m(*fD]!���;�("-����ڄ���r����ʕ���D��
Q�Q���Tu66!���n.t��kK�a��5�KdE�ڶ��E�<�����>  �tD�4NQ�����S�r�n;Ԕ~��(@(�0xjbp���w�qU��Zm��v���Y�������(��D�q2a��7dt��y�i��ᗧ�ӭ�>����̘}9͔�񀗗N��2;��f�<2�Qj����b燹��τP��"��f�n]��j�F������3��V�5�F�W<{�F\n!. `�wb=���ڊ7h�!Y�����cn����c������6���MA�ҮQW%.��[ wj�XP��7�w:��t%k�ߏo%����Q��D��B������3VAg��U�1�ڑƝz:����cT�W���3�=��/w�o�5���������óBW��"�Hd=O^�e����]Zcv]R���Ł6���MA���^g��5�(%���$��(D̲:��NM��#'I*P")���i)�/��tue���$������`��2�u�T�,^����
�U���(�ɱΨ�*��*a�j%P����F�T:ʬ6{�\Z� �b���@i� Z���CW��>����w�H�ʡ�8�m-\��l[P�fD?"�M����j�0^���FTX8`�� AɈG���t�RL)!�u4%��%z��� Rl�2=t��EEp����U�&�"5˕����?�w�G���.�>������C$+!QQLY_._jYPՂip��H��V�?�g7k4m���>���<Pʅ�¾��2W �p�Q�`�V>�R�\a�����f؆axZ�*��w����әt�\0Mh�hs�Ւ�.3�ռ������y�׿�+>11ﶕ*�%N�!���E0ҫ����]��e���3�ԡ��CB��X�e�Q?X��*Y*�ܼ<5�E���C���ש��E|���_�c��V������4��L
�ku���(��]Z�f�he�*HS��5G�x����$h��ٟ`�*�^Vh~�Y���v8�����Ln�:�O��s\�Jbi�=�s� o]����޷�2R��l�>�vw�r�����wyTT���V�¢�'���^'$�������)`��'�8����1��t�]v%���{/h���� ��w�%j**3�ZyKn� �_��q�:�z�� (����������+ݜ�nvX��VY���^��Nu/~��.�y����俍ZӁ��?$��V�G��>�E[�P�b��f�kg�{����1����FM6@�HV@LV@�����,�o-@jGPu�.�ѯG�b�|�|o�t�����Kk���:��r4��7�|B�:7ґ��� ��2����������G�db����f������x�q#[�*-��no�رqLQ�0毮��L%9�Ž�JE{A�|�x��yϛF�B���2"�g�u�>�%R�JT�-'揦��N8�)^��i���B�C�Ƽӷ�6UqopF�%}(G#e��6�G�7
�<�N��>M*<�g�����8k�>�{�[33���Y#�Ֆ�x:bHIUB�}��Y����̀��M�=]�x?����\�>c$b���H�_V0��ݎ��@)a*��kyF�Ӹ�M����7�� ��P����|z��\��lB�-�aG0kn�RPD�Z���.��6�ˣ�<a�W�5��JY�k��L��'K�$
Ncoq������KAN���&CO#�gy�����ˡmM�<�U�ڊ�x��'o3'[�	�lV�
����Lֿ�Ky��NS����q-�qx�P�ߨ��).[�-,������7Ij��BŢ�_+��M���ߩ�r:L,��eB��$'k������];�qp��@���N"� YS�|�\
|����GB��Ǹ����&�����-��`57�J�6���^��S91N>ߊ���N�Y4�L�����|z-C~΂IƲ�:	��V����٧v��p/VvH$)�<0 �`e��&���խE4�9�s�9Td�]2��W�>�R;�RZ_��^H��ʏ�є�����r�9�������[U��D�!��_�q��7Y\+"SM���r�<~O��|B[�F��wҾ�P��n0�ta�"[#��:�v��xa��ϣ���07��m�Z���	^�mv/6�\���D*�����p����w���T�3������qr�_��{��]�`��I���v�T#`n^rǡ��aq�_hTFY�k��R	̩E��	�H��3~�q/��U}ّ��y����/���l��#=o:����Gh�た�8P�U[�!p��B"b4����Vb���S��l��Fgv?������ֺ�(����W��=��P�x,��� {��Q��0���*�h���ܚ�$����'��*���J��j%Z�.�톎��ǭ��=zoA�a7v��B���\�@v<�l��q`$���_���i�}�o�.O������b��m`[R=���·�f�%fD�O��o��XS�<@a3� ~#V$��
/�LT7�'�������*ր��W��3��{����[D?�s�[�|���F����[��&R�_���x����X��9�rS�f|�7cX�[2Os|���+CX���utr�U�]������>�G�p'�_��>��}DΙ�ܡ�B�$W�����'Y�}z��{v!�!C1A�Pr�\ev�-��5\���Y!��m���Z�F�7 M���r̗55�>������Fi��%J.�>���P���}��k��%�L�L��#�[��\5X�:��첇��~�����X=\�<��ߓ��*��sO�Ʌ ���P���WsQ+�c��*;|s��j�dGq�c�ȖF��K-G*��(.��L3�.b��0�$`@�5�M����8�'Iֺ�	"y(w't%�h�>@%]V���c�R6�K�k���7X#�s;�2����7Z���=F7�U�u?���X>���7J��L��a�o�B��>��v��q�z�m�P���HKt�9w�I���nc�8bh���k�s�E7WT&��"����	�7��h!�Ϟ�Z絮�n\� G���	��:�02�i{]"Y,��8���%�5��;"�\d!��c'7"�� U@�����R}_ӎ��"G`�A����g��z�n���f���zKC��)�h��8�;!lI�?!b���b}f� ��3���X�jTS�<F�Qi"�b�N��GIU쥆T�J�6 u��`�s4;��t�ܪ}����C'b��������y�����h�A��Q�La-q�B��8��NGȇP̍0.	8A��j���혀.b�	�1')AX	�����s@1�ᭁ-0��f�쒅�s(K|6*S�����%T����s�ˏ� �8����'��-]��d���'w2ێ���س�'w��j;�շ����( �訉|�q�`�)̥�h;].6����'ܤ)�"��	�Vޏ[*�Z@��z n�2),Z��MN�4����p.�kV�0	�Tޅ��}�8��٪�����k|omv�lG+� L=�/�d�E�r��A�tݻ�
�-����kِ#k����Ϳr'�������n�xhvǔ6Fc�Y��=��kv9Am|� ��0*Ù;�Y+�AO�C���қ�:<=<)3����g���,fk�;| N���b���4�a.2"��@8��_e�hyv��o��+���ϳ\;��gԎ�f�^�r�<�2�p暼��K6W�\6����-��B�?��5���Vo��v�5���K\���]�m$2z���.P͋���\;�wc(qQzɆ.�FG��&Ǭ���H�6? sܺ��z2l SF�s4��~��1_�h<��|�����R|r6LN.wL%�=�H����l��]]���:�~�-���i�|��1)E���!�Elg"co���k�ƖH&��3��]D//0u����KWe���~���t(�4�zi��.�g}Տ�|�j*��Uu�n��}��nc�A�gE�l���E��Ye�sҖ���С�A�S;�Rw�88�P���oT�(VV �oaf���uw���yV����<ɗ4��e�#u��f�x\_p�j/�%ϥE�h_�(a����K����Y:�,,�������[���~'����8m;��~���ٖ�Nw�u��A�۫E�tr6 ���)�@u�.S(� W��,���
P(l�i��r��1�}#��W�>�eE:F����3|�Y��W緲2�R1�Hڝ�I����ϐ�em�.���507y~�V���?��l7G��-j��8����1�&o�V؞ )T��_�T��%��H���dUq��ז�d�utJ�����92�����t�
@���0Qu��0�5��I2��忾��ao��=(!�gE(�_a(8�Z��1L�J1� p�l�������e�&���?����~�]�x|�i�m#-�ȃ�.�����x�I���0��)�/�S���cn{�$w�OB8cL粧�#�a;1y�V�������7[c/-����W��G��#��w��_�)h�ݷ�෡���C�w��Ÿ�����q�a��{g���o�BO{>�`���w3�b�,\�|d�v�.~n�Y15��9�<x*H��6ཛྷ�Ms@�,�h*B>O��r�n⎹�#�;hy��J��ʕ�{�cj���?|��|�_�*��ٺ���Dv�RT_7�5�����[l�_���
�����L~��Ԡ����
�t?��,���ru�[Xc5 kB�W{����qR�<4�?+D�[��y�K0�>'��zZw׹�h��2)��2���UF��y-��A�r'(Ѣ�p�9�Ou���_�͞,1��V<����}t��ۊ���A�y	�Z�;2�=�(�-̌~?;��K�䛳��R�����_�*�Y����P��@��2��ox(��oA�\�$�Ǔ���קG�L����Z�+��Ü���y�Fkc�}�\g��_�P�˶Ȣt�����Y����v���-�9]���.�����G)�ס�5��0iTEJ\j���U���,<z�d��|���g�Y�:�D�k�p�0@�KY� ����}��[*C��t��J���d�k�@3{��$E�m���k�w�Su�%x�al���bd�/����>����.|�o~T�T�������� ��3�����=�d6	�?��N����?>�.]�����@������^]H�s���y�v�3͟ �m��ZБv���R��[7d�����'�����ES/��p��#Zjx���/��*
P�.�x�t��Hc8MsY�\k���t���K�._�u��M{{)�d��!C����Rִ8gn����tF�D���#��5IjM��ح�e�S���¾k��MQ7vʯE�P��T�{�	�F���$���c~3���)ha�Ȧ\�{�1�:z?�"���;��͊�$m��Ȇ`E1��*1�M�LgNV�%~LD�#��� -�QPEI�A���7T��S}[+��w��m��A+}e;Q�cTV��-�s���u@چ��g'��bB*��D��5��G���Lm~u�Gz��qjv�ש��#ѯ�������d#@2�@�����Y'�꽦�V�_�H'I�&_ҧ=ֈ!c]qWQ�%5A���+c��[�,l|e3F��X#��9׷����0d�1��B�ny�$Qq�ع!DLZ����a}��>�֊�Z���2≖*.{����Y�ȟy�Oz<����g�{�����N1E�ie����5�'e�&��y��Đ Y���q�
ѦT>��ǌA棩��Ѩ��L~;m��U��Һ��O��������&xL���Zu?(����>�/"R����h��OiՌ�B�]wq.�,�܏�^��SLYz��'���=Vس1�ST���}2ˊ��qq�)��V�����q�Q|q��$7���w�<҉�!?���ӽC���ڻ�����RIm`ߛ�U9�i���n7���	�lF�bb�dF7'�� {�	��V\s���[j��q66�k]j�H1�9�h�鞨�1e/�m��S���E]�,���� &��^�Ϯ���p�b*JQ�6���6�����%2�2?�����)�_qT_���9
L�{�tM�nG�a���E�d��Ռ�v}?���>"IY�^�8���D���(�?-������z��\d�[�d�ObJ����C<T|����z��}�ұp쳛|iߙN�g����I*IXL��W��e{�����4E\�У�,H?	�p3�,l���7>�׳�ӫo���rs��aQ$���r默����v��g׶����D��.O?�hƣo�ݕj�r���zmbsa'���~�D���s����oU�x���{j}C���>{M�-�h-���H�/y 5l�h1���D>Y^��m����ت���vNc�DS~�+��h��)_�d�i��W�B0? ��"��t8��5�*aw���X���?�������z���VE甄�,�VL�1�1K[���m�������Ҫ�W~'��v�3	��vm9�g!TA[x���ڸvKmb�;�\��9�#�<8��*����^�s'���ĔB�f�R¶QP�!��tcS������Eq�q������0X9��ĭ��2�t�:���.�x���Hӏw�2�M~���~s��۞{�i�e�n�Dɪ*�-��^?/����k���������'�ѓ�sЈzZ��0��<�Wޫ�\]]ֶfk�"��O���[�7[s@bR��td!�������>�#*7W~�^�RNh+����o�f~ y{��|m��S;EA��W��Ka�D�������N��t.��m�2(����B��@1Ը�V�~�D�^u�{ :<�
��=�M:�\~�u��\�di^/��\�%��H�8/U�*���iŹ� ;����ND�f�^Ju�� ���sb;�����F�]Z��Ƈi�'��j\��W�� ��'�>(�������o�on�$�ӭ�vbd$��kt�7�?Q�K;�h���}�}?N�6y�#�EQ6��	�����2)�t�&m�9��M�D��ylz?J�Fb%K�� p|{�y��<]��m}�HJ�ߢ(�;��TRa����`�0�����\QEfcH�M����[s_Q�Ҭ����k�
�\Vl9>J!������5QW��=s��1~�P}���?.�p��"����ٴ2Q�]�)C�*�֚�?�^�w���~"��:?�i���ݦ��@���N�"da���P������{$��~�w҇�R�Q]~,3Q8k�.0�������n��Nc/���<B"[�b�0Q	ן���5\0W�'�:``�K��t��l��.;ў�G�K�r@��SJ�K){��$�q�+�ޕ��z*��Ԓ�p7�Og�#j���u�Yp����S:�_�[�1|�(�"�Ct��h���s�`:^"�Ѵ�X�/t�Nz�É�r�~���1�!�Їt6�?[��TQ9fú�M��s<������ŕ�Q5���0f_Q\�D�4��)K[�U�M�cv���Q3�8��٩&������?�M�{�N�S0�xI�q(>�e�%g��c	��Ҝ~6o6臖c����84����Tϲ����죪4@v/?�v��8e�Uڥ_(y�� ʇ��:?�K��*P�S�|�q�����ƿ/�Chd�mT600R�)h����t��)�U�G
2FI���0<��\�y8
{76����w=��럩C�cQ��H��Ƹ�����,޷��>A�E�'��ǠL�(� v�O�rGv�My:�����/�쮠v�f���������}�&�鐎i���ΥQP:���ca��X�٥s�������?ߞ��p���޹g����g<��Y�u��攉�P0������.�5>:���1�����F�scd^�+�NXR��h\��]����[#x��K�McVZay/��E��W��:b�c���} �n�eh��>����i�K���qQ�'a��4�Pl㏒�w�z~|sm��r��`dK"W�I��eRS|3(�?e�����t���"��s���EU6-ǜj�+*�Q��_!�
�iM�F�CZН	�tA	p����<	���e����vV��d����S�L�-i�>�}��Z����������\�
^���]�[����R���b��&�R{�3�V"�L�V"m��L᫴��6���t�K�|�~x��X��y��%@O�[�C����;D:[�[��b�:wB9xBY?}�-<a-f���Cq�a���g����ԿىU)D�q���ʐ��p�q�-8*�fx��CN�1r`���g��Ņ�������k�joc�<���eP^�5�ض;2ԝ�)�Ur���?b����,�tt0��f,
;��J��Z���Q�t�%���ǡ���9�pWlgQ:�R�N^E�	~}I("a�u״b�ؐ�I����8f�&�ڰ @y��9��g-B��םЇ�V�������;�N]��jY�T��-2�ݲ�F5q�W H(��T��8c"9:ӊĘ]�V�6���)���_�=�2��m�z;����֣���bv����,�?��}���{���<|덵 �+��?��bS��81խ�e��q�� �����I���[qJ���W�!2�m���1�]��I(ܺ٢����؀���z{�)�`3�u�@h������C-�W>�m5ɡ��[rz��I�{� ��V�AA��<��r������\���ؓޢ��ȣ̋�	jN묡�mkiY�ը�V�\�H�;]����aX�P�iŴ�d��w�C�UPoZ��5���)EL5S��x]qeg�4*@�{��5i�5�����"��-�$�n��6�x���ϣ5�e9����A�������o��w�<��������F�;��Ũ��a�[�ArzU@ ��R��7��Y���\��c���(�~���.i��E��̽��^7w�m������S���M�Q�d�����1�(�6�Ӈ��SN�i7��<�8��y;l<�?zϖ}�p�����&��K���F���\W-�~�#��H�*��:��mo��`{o'����		��B_n���:��˸L?��￙�m(��%�0m2�,_S�����E��n}�v{��t�u������Ǖ�K�>{}����ѝ���)�C�~hh����a7�Uj�3�pfX9��Eu�+~�'����{8�a]հе�J��������7�t���ᖰ|E�a{�,��Y3�Q���in�qK��q���஧@�R5a=!�}*;�������|V����M�9�9���vΒ�u<����!J������ߤ+��B�e#g�����w����`����
��6X�����`K�[j[�%�����^'-T ����̈��0l���{��iio�Fp�H�wWը��$!�I9�/�q�n���u��w.b��6x��(����dur�o�@vc�Өr��Հ��r�L;���	�� �|ֵ�i�:��~�>�w�8]Z
3魣ɀ8�	0��������5!�]QQ�������fЮ��%����/�\ۧ6��w	���E��}�5\��`�n�^3��!�*I���:'�R��мaA�"�bln�aX�~�B�������eL�Ň��d���*ڗ�p�xV|c�Pc�%�,T����\��&�U�A������_s�"��7�&�{�#8k��k�r�W��:�ǒ�B7L��,���%酦y��[(�3��ϟW���{�D�5-=߽���ׯY��$��D�{��)h�����r��w�� >�Q�>���o��XE���%��SX�~�2G~{�1VN�!�}R�}�u��Wr��g�ظ���	wm�r�/��{�Ea������&�d��o��;��/�?S$�ɧڧ��=�v{j_�~>�6��yW��f�e�tg��f�j�#�3:�6�	���`2��0��p�جr Gǭ����@
c�עt�h�B-��NR%��4�u��x�M��B1zߵ\�­�9|���"�2�Y�\i��[ͩ�VYCj
B?�5Eq� �c���˯v�_"k�(]�l�(�D�L�|<8����H��i��t���
χV�X%�����?~C��e1�c<�,ܽ="���<s��d�^]��^�pm��%���>3\���6�p���)��˅���j���J�����^��eH�������=�$W�W���]|�f/�� ����0?K?���BL�.H���m[ �A:�݅�9�!��`ٲ��j���hY�J���p��4���:�F4R�ǜ�Q�>�5���s{ݾB>!�'{�9󓚪>1$(|��?{�P�����>n��J�w������omܽ�K(D����&����H�P�j;��?�lͩ&LA��Ɖ�||zoM툧������_�IV��x��'U����[�&T��w����oC̳�����I��`�\{��Y�+_ڣ ����+���}�������W��3��� �'�|F_rϩ�n�]ń$�>�� ��O3do�R�\S���l��t/2F��~Y��Ac���(�6�u�^/!�����i{�I�`،�X�����1��d0 �J@;|����P�c@0F������F` Feb!-9O�<�J :~�����z�̘�J��kH�j�)���O���`@�gǕ������/�
7W��Ύp������$�?���n��K�DL���Fq��74==�ޥf{�$���*1r�*�3��Ym���}�����b$V��5�V�u,��~+����x�RkRߥndK�k�F��g�yY�2�U�B���|pҳTC"���<9z�l͔�Z!�@���TWG+ �rVkH�`��E4��`'�f82�vb���\�%�_����,���JX�QƜ�
u��/���R:�U[�X]�K�K3D�(������e3z���T�]���wD��zJ�L<!3 �>P���:�F�*�4n����.*D�n�%�l�`~��bjo����� :�]�VO��Ȁkw�W�?=���=X�����������1�U�|U����rb��*6���҃Q;�'�T����\w~4N�_�]U�4#�4:��2_*K!wy�k
{���l>��<��7)&��3Ы}WR��(g�S�:R8܆K���_�}�}YԹ�C�,M�����R�@��S�
���v6`D�ѝ\�Pb��X'x5��4#l�}��M(G
ñ�3C|��X�ы� k�<}���2�Np\~LY���Np���{p}.���󚛬~Y���r��v�rHx��w�~���Oc�^���ARr�DcJQ��Ї� �o�-�Z>���m�;�Y;8,��;X1�����CEOG�.�6�?*����Q%*~��K3����e"�4W݆@���TD�XF��=�����T�Wn}�|�p�̈́M㠜�� ��#�I���%�ٷ(x���xFIh���F0��"�� ��}U��ى`޻�����z�����+��\DZ���D7�3Q��{�������-n$i�p�F���w��]M��9*�ՖR�g+�v���Zm^u��%nK�3���چ���yo&)�iC�G�}L�^���hd��������a
�a�j�$�>3�Q�*�ޙ��8��Ŋ�7��5�$�%���$�kף�%�aA�zAH�m����)�fj���� O�O�'�w�=N�E�i8Z��E����� �)&	��z+B+�;Kִx�Y��-J���h������|������4~h�Ȉ @����=k�ig��ҋ��ۋ��@Yns�[A9��~@W-���U� O�E#_r<-Ӎ��Ҭ%�,'I�i�<z(�i�ϸ�X�����5=1���z�L���@O �Yꐴ���SڶI���0� ��qm �}�Qv��$ZG>_���K��Tg�d;�À9ۺq�WL��[��]�N�]b(�2�7�]>�rS�}���<G�p��?s�Ňb�c!r���M�3=�mΥ	4�)�a(�ծ;��-'��/3]�{���/�2��ȋ}O@�����1�����A����fC�(¯Gw�*�����s1�p�'юQ�l�����?k���c�VVw��S�^q�D�3�(d�I��/��I��X�{J�\«�^Q��-FWS܏yO
��״Ph�X���������[��hQ$��Ef��}{���m�G�5QR?�>U���K'�a�y����������L���-�"�[3��/��v�/���ۦ*_�{�5��5A�ԯ������سn�3;Ho����OO1��R��GLk�� [��=�Kh2��c��;��v����eA��o-�����4����.a-��z�����J8/�E��g���0�%�-yY���]fj����~R�N_v"�^K������W���묅���>��L�B�{i���aK:T��'8�lˋcE{n�Re��L)������;�'o���I剏F{zt�3���Qv�l����;\i�-���M"�Z=��C�q�[Jz3_n5�4Y�����2u��}Î=�E�u��19���4�~��v98�&�{�@:A!�3/�'��ص�Ѷl���]����9ȳ�/��sV�۞w��~����+�Nŀ#�%Ґkg�p��_7��#�ჺ)��<��-D���	#m��G�;&��8c�H>�vV�/2������0?9��|�7Eڤ�E*���F�?��� �,���ж3`]YJ�v��J�e��7?gMm�ϔ��J��	)��yK��}��5K��*&���/�e�D�Y0g���Y����v�uF|t��L?���\���zJS}l�[����t��ʢ�<Z.�
*�d��`��6lpnC�.����N,�,��cϒ�&�
�\6�xԐ��\�z��0�o�����2�Vk��߱0��0����=�·���a����`+M�c����t�DCe􉭟ՄO�\�^~�;�w�ȣ�LA:�O�����Ydޚc?Ԙ��e�4O5��?����ig�`�s]:Qu���m��d粵#oQbV(+;,lqn�B���`K>҃��=��w%����&�6ΰ\����2��)����(�#V �=�c�W:�Ǫ��,�]ωo�~+����&����S4���+C�3��E)�Y���_�}�k8��+������}�lq�'܋<�P~��Խ3�7��!������Sfk���퀍���ʐ��F}�رUC7���0,��+Z%�"��F�C��������i���	�Ǭ�3��O{��'?��rq��բ�w{.�_{H��DS����k��� �f�{���NUQ���Q�#;;�z�\�������}�6�3D���Zb6f?L��'�Y�����pg�n��(�ޑl�?#��m8q+rژ5l���]�1LEi�B�ȑ_5�a6<� F��H��Ww��/
D�b�y�Z[�ai��دM�z9���fK��x~\m��b�7������q���]�R�.�v�3����Mn���u"�/6/� �?�r�%�,g����u�%��с噯����`�bd�,�}������VG��s�W��� Igw�mc���`ݙ	d/�o��N�<A�hH�>g�ĉa�8H�d����Y��"��\f���zJhe������.m�f$���L˳,��:*p�O.:˾J�f^)MK~�v�`1pIu����7�&݂R-9�&�n5W����m��ua�MC��AAl�4�����Ͽ��ɖ$�yi%P����I���������c_7��2�Mn�M��ͅ(2"��8��>�PM6�	E�?
x�X$�"�,�y�؎\���'����"�iZ��@��U^s���8Q�ŚE���w�M��o=�Gx�����������ě�����=�}{�vg-�������ʔ
Ᲊa*���'�Þ5bއ�.S�
�!l�|.��:+z��'�fU�� �E�v�`��{������y.	���c[�}�氍�Oo*�����)_e�E~���7�Tۨ���ѥ��R�����{Ӻ��	�#�����)ZS�)�/|`x�����8�n� N�'�Đ�cn�|��9���sP��C�V
o����i+�b]�?�{a�"L��aA�X3_�@\݆�]��6�ï��2���@	N*�f����O�6◾-�����V�G�>Id6���d�f��6E�rK�{d5�v�Wtpѽ/�ᛴĤ�l鍩�.���7��v���2�?k��qK���:co��_u �g�H�X�n����i�HB��)Y���C����|v+��Z&�+���V�aI�5���T��3�d�a.r�n�u�����λ�g[hj8	��BV�	[~$R�M��Ix�q��W��1Z�B	 �e�M@�����d?�3��U��w�w�`9W�[d.8�
���a:�ۼ��i�D�U�u�Gh{Nʿ�'��s��!sE#v)�GbǺ��f�D�C ��X@M�L��2Ƨ�B$�<[sr�e�׿qt�4��hv@�B�AN��7�Q�c�u��g�g?�� ��*l�W��#����谔�2:��l���-z��B�)���O�i�~��iZ�� �w��C�����.�V�hr����?��@���Z;m�{p�RtǛk>7ݳ^}#ῼO�<݇�$�l��ii��(�������ǇϊQ�4���(!I����M��G?���u�z�6I��Yh#�׆��y���v��݁���U���d�w��ͨ���G
�(���F�J�O�0/MU�6��$�N?��jg?����ֵ5io�~���,�e��Bt�]���<�D�Ah5\��-)�H��b}Qs/�:R"qK���I<��%�w��Ha����ف}�k���8��G%;θ���XM
sD��o7���>��.����~A��I2�P��%�@^M0`�G&��F�<�7��tr���^Aa4�-�)��i��j6�i�٧���0��U��E�U��E���(6��9�Y
4��=˙7l��A����$����m�ů㿋�0�E���єg��-P%�04��`W��ȝ�al�Ĳ�^�Բr��<�s$v):���}T@�R�^$�7�����V@����2%_�ܬ��u­���6.?������m�l�k=��<�*�����1�`�=���m���]R"ǁ�C��=�Caߒ�s	��3���/��(Qkd�3�t���?�E{/�"���+�[�Vܷ�?�ҾM�i\5���Q�rd������}z�B�̞����ȁw�RmR��t��zv����৩u~l<��s1�xt�K]��/Ϳ**X��;�"2��4�.��d:��$%\}+V��
!(̭|��Z���y�1+�䅎6JB�j��GԘ>�V���^��>)�m4�ֲ�I�1�>Qѷy��y���g|�4���쀡?�0;pmw�U�l�x/6H߉!.�9�������_ٻW�"Z��M[B�X[��A*/u�֦��]���Mf�0��?����H�E%p�X�-4�wk�(p++5R<�'A��V��q�H�p���>�~\9d0���J/���_>� V!���*I��Y{mY��8Г��H>KLb*�=Ɔ��EK5բ��A�K�^�	3���9\�r���E�׵��&�K�aF�N7wVmlہ��I#�.M�Ƽ���f��Ůb+�72P��P��`��.��kLKH�w��)�/"ղ��i���z��>�W�Z��pH��{�0�B��UV���[K�6�Ŗ���8�G����s#O��U^)��(&ؙ�=�k"�7_j$|%�uO������C�m>j�ˠ��7����ÿ��Β��h�WZ��i/g�s�J�;�'ؾ�%�
 ��C���ΡJ��Ѹ�&�s�{Fb$8E�D�����\`5�f2�?!I�=˅b&f��<]�=W�X�����F��ɖQ��!��iQf����VyF�8���ƹ�N�0�䳷����}���o�X�������X
J���0���?�fj�@Cz;FU���^��P0�C��}������`]��#�{�\(�+(�tv�Rt���#BA�}��TÇ��rQ�/�k�VZ��~ki[/g��Z���0�;���k`�ϻBשR�g��I^FkM�Y�[�CӾ��W�'x�PM�=`�����g��л�3y���Ы�7)�M�(ui:���c5�:�mwB<���
y�e&e�8���K����*����*]U+���������5��Y] �!ŷ�wW�i;������A)sͱ�ōi�h��
�kO�9|�H�#b'�BP��%�3.M��4��|*Ot��h�M�^�`��,ͽ��Lj9���M0R� 0�m_u�0C1Gq]🇩b���^�Uk6�Z��Ο�u٧h��=�@��4��+�`ْ�U�m��B*行"L��[kj����Z�o���8]��=z����F`��/`���2:F.�Sg"p�h�R�]���j����,z|$�FpJ������D��N�
�=풦�
엛��J����5����e�����ί�g�U�Q���M��yV�M��U1r����T����h0m�F�wW�'N�N}C���V*��\ ΐۍ��[u�.\�F�t�d*�IM�~�t �A�v���Z�����]��-�d�L�a�g�j�̞�
 o���I���ᴖ��3G'V��`�d
�B/͏�|�8> �.c��֚F�J�;%� fh@)�F�6Ȳ�u5�P�W��(V(��p�����[��'Y��hv�'������eż;�t	B��5}b��{�1�?�� ���'��\:A~�^��5CN�͎��\�1�Q@���'�5�.k3�OK�o�*���5_�k����h������:��_5%�!$G!�ǈ��#jVZ:���
���YM�_���6��訞9R��O4�7/���֜�<�Ǉ��R�Z`�{�h� a��Ҏm�M�}��x�]�������v}.H���c��o�̟�7x�K���Î��۫�T����>�EN�\����>I�T#�T����6FZ˚�T��Oe�Xm���N���}��?�H�i�ND�t�P$j˘�`Y����E�]��������c�J���NmK��zc���K��"�� \�|B�OO��ٙ�j*C'8�f�e0�|wU�#�E�ã?�9�Jr.ޞ����lݎb�f��O|�E
�I[�*
?���a�}W��Fj��q|���'����Oi�@U��QlN5���^�_����M�͉�q�sWtWGU!��{�sY�7Qï&�S�w��
���'K�g�G;�]�=k;N(ֹ{,�U/R'�p ݬ�geQ<X���r�U ��]�{m7�8����K�{w��8��o��.l< ��
���)�OJ�怯�F��]t��$в�Ρ�ױ=z��ex��o���Zɍd�9;����:?Cu��;V��?!3�Ie��$Z�\_�����Ӆ;C��ݍ9(Ҍ4�S��|�Ž�t�O�hL.�Oh�`�2&�w�n�h�XC!�'[m\���-.�����Z/��QA�6	�L��d]�W��m�u8��ZG;����F��3_��'#�5f��r_).~y��pr�ٲ#6�S���mFg��@�������U�k��`w<�����b��~M�B��m�	?��j�������$q�������Z�=[�sDE`-�s-`>K7�iˠ�po�"��ޡ�3~�[e]��*��'*��9����ũ��>�
��Dj��4מ�)5���Kc���N16j7�{,{O��.�'k'��q��O�l)ݭ�dJo����2%�-*�i���{t�j�4�A�r�v�U3>����Y%�x�oR�B��Ʉe���z���E�k��{�}�,#��������uҴ�Ĕ7u��W�[tѠU����=�h�z�#3Xܨ��-kZ�o�?���,v����v�����l�UÃ�]?�ϽA�A%jK�b��.:��N�4� ƣ����n�O��Q�u��vy{�u.�dQb�d&��>4�'d��j�t��Iy]~t��~� ����ɮ�X ,��[x�Xt���>Z��\I�~�&��ˉg8�	6�tӶ��[^Y���3�I��{)���Q��؟����5&	��۷!�Hr������h̖Zٺ--���#*/�U�J�wǜ� ���pו
dW��7�(F�%�)�}��d��h#y�M�s��7�e���S���&v����$��犏rF�^��5�Pav�f;�N=���(�I�_�O:�o�G�����Za�4�L*�hH Ӓr��JBg��b��/G[���֡:�v�76�k�;cA�y�%>���A�8��E�މ�~��][N��u�*�}�sm���DC=ghک�&�B@ �}�;[9� �+M��]�=�=�4͝'�����\67�E�������c����I�y��Z[�L`�@��X��SH�#�a��-^���=��"�Jp�^�\%FA�E$�Y\��/���O�l��ւ�^\�H����������+(�P�v���'z/ao���g�����qi�k0("x�GB�h�1������_;���;�'�����z�y*!��Tjg��hAz�V_v�p���L��n>4f��O)��մ�G��|�PrsJ5�1��p٧�ǖJVjatS�!����c��?�4�rb�݋�]ΰw�}ۍ�D�Y틨9I����r�$"�o�P�b,l��J[�A�!���'�i��Urg�٠����#����n\�\Xl��1�?g� =7��ׁ����ܬ��q.�_�nἧL��(���XJ9ӫ��y����x{K���ߵ} ��W/�Uc6G��E�~������e~��A۷��[g!��v�^�+@r"uH�`QgXPs5)�M�W�,��g� 0o�\G���aek����
���4{�H��}wkǇW,���x��7!^�#�B���p��v_��k��I/���ݜz`y7�4�����<�b���Ý[E�V�w(��&�.o�5�|8��>oOW�?��h��y4�E�[�i.B� ��[��
�A�e����#s�:�����5��(�j�|i������EaK���ȄT���_X��"~���\�(����{I���8��\����l����_>��9OQ&DzW]4\<ĵ��Ջ/H�(Z����>����lc8og�4]�W�� ^�jkTA��쪚����mz$X$�Xsݤ��.<�+;%�E&(���I_�! �s7|�α�4sW"tm��,�,q��|���<������A{6r��:$����˘so�j�l��=/��<$������G���}GLldV��K�*� ����	i��W�������sy����I�!�m��zܐ�a�p�u�O<r�IstGtwY�m۷gJ�%L'XG���n띭Vb��2�H�ق��*$��u��j"��\���9;<�.2~��Ν�{-z8j-�!��ޮ�ylP,Ao�$AaE�h���bU��K�o��/���0q���@��5�/S'�-XP�r:�EU�,��^����`���e?���@�v��<�d�є��Ә8����E��^�7�oM�a�0y�b<�F�Ma�i��=v)�x���v�,���P㊻LqcQ�F���0x��r�m}�WwOSI����𑼾2t�M��ts������+�ێ�R��.�>P���2�4�yr�-�j�M� M�X��i�圖W�!AQt��I��^�Ȅ��~�.��i=� ��-
ī������_�J��ז 0h�F���Z�<��-9>�B���bv���WB��~Ў366l�t��{�J腈v��j������v}�E'��֞�@.?aaaD�]Cў	d)�m���MY�87D;aväRi�*���J��:��wn��w�O�57�h$�&zt����� l�g&w���(]�5���Β���^�����oww�GXz<�%С���&KG{�{E�Y��i^ߕM]Û�\���vz�E�ibm����� z{Y�Jb�qly���0u�z�`1�=2���%�<<��<x52M{w��TI-��v�?���E���dc�}��U��N+��)�x=Z�F�
=���7�!f�[�'�v��*��[1@���d���3ߞ�K�ޟ�x%����䛻D�v�dF����`��4���8>g�i�������./��x�4�Pm�����y8�/"
�*e<��d��9x}��ͮHuʆoy�i;/����������}��)>�h�	o�]��� �������� �xp�jXl�!�f�>��t�8�Oa�3�-Z4��Y>��R^�J,q����OԿ'�/�cҲ6jR��`�s~�m1>
S*w��s��a���U�-s�����<"C�{�E�JUl���7.� ��L��L uAb�7A�KxL�5sW��'���q��B���׎��r�҄U3K�{�<yy���g/"ߎڥNL�&זM?X�-5O&��n�����|r�k|x �/��M�rҬ�������aA���x�J��P��2��&a!N��,x����M?O�D�^4��.��S�s>7M��6*tq%ʡw.Y��1�]����W��.
� kU���t�m ���tN�it�ܢe�*���]'���o�G��i���B4$�M�d5�wO+���\�~�r� �牺���0-��Wz�������i�û(�!��ߧ�1��`�wWk��ܞv�������g65��S��g�7�Sk�#tI���a�>;^$֯m�����|/>���Ý#<�
�I!<�O�r`��V0�)Y9vuQ�<Bw/^�����6�n��S���d;g�Py���.Ѝ��9��+y���I���+�:���h��ƛ�-.=�*�<���M��)����{��nZP�'l�HW�2�-�����Mz���N?fzRX�{QX��WY������_�#�G��y��nF� ���37A��xМ:��5��ݵ�)p��]�/&�=d�$�%�YS�%�jVnK�Ʒ�=�%h�C=[�i�߭�{c�"����|b�����:�2��jZ_ي�u�:G4�q*����⸽d^�oc�/HL�{�E�γ�J����BF�&{kf��0d*q�A��5�睙�g����h���bߑ���M�9���Z�|�r��5W/B M�^<70��~�
�W�;�2ف7�g�'�{_��o����g�EbF&R�of���?�}Q�����$ڃ�*w��J8��Α�z#Xp��z��i?���'�a?��c���qb���p���L�:����Q�a>h6V�ϐ�V8H�ٺ��v7i�ƴ8^�Oh�pa3-0�a�?��������1�K�zR�R\�2�q��x�%d)�aWf.G�w����
�=io�&��e�������C�R&����/tIp�O��ji{l9�	���x�8��7�Z���n�{�Udl�u��PY��Чd�)q����Q��.i.�������>�ϒ&�֘=�26�.vG8���OI��9iz��~�u~�L��?�u�/C���p�����>7��US�)��f���~�tX����.��~����BE��A��v�Ejc���^��Oӛz���f��y�A�����6N���N��7���lñ�	�e��*���y~�:��=b��!Sf�d�4���˦�������3�U((X�����$�F������*��<}gz�۾������G�w��.
QQW�̂'��P�%kT�q���&�ޫ��Y��Gz����?���_��T�?i����7�l�����{���D�G��٣f@�cB3��Ģ)~�O�����"�9*q�8���^�PΌ�'�]U�&���[��j��A��&�d����Em>thl/uU�5��~4��L�Gg���C��s�o�w6(`L�^wf
g5��
!u��UŁ��4��_~=�m-6h���9z�x�57W�3D�mv�)�C1q�q�`W�w;,g;k.��뇜�sv%g��3�(`��1¿`������B���q}�=��ӛ��~2�{��՚�<�|����9�l�t�\��w�Zq�Jb��cx�R�h�|k4�ۅ�����<�) ��*ʋ�W��%����kƮh'!lf�{
"y��y�ccq�N���v[۶R���=�h��]�^��8+(��`�SY��0�SA�(&7r����X�D8�����rA���e2�`)oP��� Ǽ�+$P�����x�8�{Uw#m�R~�-Ta]'��`P���1�dԧk�����8�<�2��8�l�;m'�=�ɞ!-��BX]�N)�DN$[ǎ�zMf�����ܒ�&� �������P��0?	�iX1FȠÛ����_1��-Rd��~���sW�N%:L�=�L7��+S��h�E��:�ziC4��� z�ZTbQm�����%
*��ro,i���sg���^/͗�^�/)/��ʗˇ�ZWiV��8���h�l""�ԟ�z�z,sɑ���*͕�̝ɀ0������<	ţ�_gNU~���u����)o~��ԍ��X��C�ʍ�o�i=��|���܄���vڄ��s۳X-Υ��������4H+�2ϳ��aFvIx�9s���W~%�rᅼ�9�Wbw7��M�M`��
��*������w���w��N���B�E�w)�DM勭�������H�C>Y�������J1zǮ��N|�&�O�PӀ�/���pgy�q�)u�e�kQH�{1y�j��6|p�'\��8��Zi���m-�Ϸ���}y��;������M��6�%���a��V(�1��9V��!3�FP�\�<�RN"H�.�����4M�Pj`0bUάL�벲/Ѯ��؅<�d�OX�����j��Ԟ�zv�,��}Y%Xx�ڨ���밿��|�-��:��Ta!s��_v`��4��h
�����b��)�w_D�=��:M�\��\�AP��F���1��q*?��C�'&33k���mu�I9���|��c����#�_^h��>�-�/U�V7y�ʀ�T>
f�+h����?Σ�r�{�����|�G�!~J�(�d�=��w�	��ha�Cj_11.{�����kN_����^pr8���˪�AM)�:�)�=	���F-���8~���m�r�[Q���I=����T�|tg9�"����j���}9��u��8)�O�8���wc2WHYS�:��ߪ!�Y��&�`�5���k����>������B(�����	+���y�V��m�VU��H6'��9�I��_��Ӽɼ|N�M�I	������d	�ʔ4R�e�p�؜U��h�!�/�n���SuX�2 ����F<���w�Qi�ၨ��L������ٕ6�@�b��$�@�m&��s�z\����L����{S2�����j_�/c�h?b���ܷ���"��,�a�;Π,0�c*�~��2wv&�RLkh���q�'��D'��w:���|�,���#3���ƀ����Vc����ҵe2�i��ں�|O�c�d�h{
n�X,����d��7q�S�i�b4/��nw턅��TJ����(9V��7���T�4����ӨMxoMؿ�����+��A6v_>0 U9Xy�c�4�������i��?�,l���Ǧ�߹�G�f�x�`\p�m�m��Y٠~��e���/��dL`�Ѽ@��>�3�ŷ�����~{�Y����R�dfssҠ�N�L��g�/ۏ��n�p@A�珳����7�ӂ]����ܳ��7���)���.=���� c*�bb6��W\l��ٴ2#/������'��b�e���e���J�7X1N�����MRDS���Mx�_�l	!ܨ�h���y���J�D��&�Z+w�QZCu�����=�`�|���}G��JA�I^z"�Vݠ�U�>iX(�O���{�^0�H�r�/?���^��(����c� {B��q�����Z2sm!-��ơE� �>�Fp�|I4�L�-��7��ѷ$_�`��S����~��|0e�}GK4�C�&����pU-��VS�:%����Q�����N��O��`�2��^�����`e�:�F��&V\��#$�$�ê���5�*��Kb�+�x�4y!8���{��֖�T@�?���b���908g�(�8����_1�N<�m4!
�U��S���>������Q�^�F=oF�X���TF��~R�uR#D@��έ��+l����߆c�Kl(��W�4��Tf��dkW��9F�U�vJSQ�5�EU23ߐ�9�>k	��4Gy��ß����J����_V鮍�Y��u�-�9*�9.>�I�!��g�S�j��dmt7�q��;���5����L�9�P��R�����b���B{m�ȶ�h���!/�5�����Z�b��(U�(
�Ҥ	�H�޻��B!V��T齗�	U��JB@@J��@��z�{�;����1����^s�5�|�g�"R �k��Y��k3�gI�^$�y�W_�?�$�>��{�;Zv�G����ɥ^阳�]
1�N�0z���G*���N�r�[Z���g�"L<Mh��/�r�D�ؠ7ҷ/Lp~�E�v�����=r���?'i�w�c� ��d1�5gv���
�۟�Ϋ��8-�ǆ	���yH��%uL���e�
���"�Ѩ؋���j�Q��oǴVj��x��#��/½Eϓ4ԋ(�/{B�F�'IJ�-�Ǉgj���� S1u���{��Q\���>�{�V��NAg��2`�S�M�_��A��z���4���3�]��*Ҙ�x���������O������s�\�Ƣ���.�]�7�N}8�V��O~���SO� ����.�_p��(�4Ч;�m�lD���d��G�s�O�9X_�����mL���<u�;��S�v��8iJd��nMҀ?xU�l���Գ���=�ۛ�sp�࿮T?�K�u���j���G*�@S/�~倽��G�O��é~TD-q�Nx�?/"�mW�_��ي#���>6��n�����r�� �^�?u����di�B��V#��P�/��a����#.��b���Y����[���>�?l��
�-���*��(bo����SW�rzj1h�;��Ɗo�\��	��M�(I�̯�?�������I���3;����]ɦ��PI�36D���6G�,`����U��u~�qs�qfYCu[.}�;�������W4��j�|PqsP/$)g榒���& +++~�HOh����3=�
�c�?���
���I�9��w����g�3�?��?R�����X����_kj�'��/yںt(T���OϏ��[���N=�'I?+�C�X�Wu� 9p����tO��
����װ���+M=�o�P�sﹲp@b��ݽ3^�Ά��'ٕS���a���&�2�@XZҒ������5j؁/�ߪ3 :��7OUsӯ˜;c[w���{z���u�5��WE���S�t3��/�صA�s�n��b��&��+^ZX7KS�<�Z�� Q�C�v������C���l|��ǂ?w��w���Ã��֐j#B���k@�����7�f�J]��*fv%�uI���;�	�Xch��;�.��p�Ź�F�e@�6� ��#0����[���}B� ��)1�Wb�RZ��4�U���&���!S�h!�?�P����I��|��ߠ޾+ڨH?h�?�Y��jg7�g��~S�#�yK���Z��D�� g4XUtWM���Oʼ��M�-)*��y��?�[$Qa�K9�`夈��QwD�RU%�����p��}�t��W�7��J���vy���	��<<�_�f�"����� �1��N���J�Yē���6ϵ��ꏋ|�9�?����1�{�e�]U(����k}��7��C�C��,l)fY��ī4crb�t�'2f~Ѧ�9D֟��v�Q{[#b��g��[4�����w���a nk.%+-�W��B�TF	��� %�fs|�M����\_�j�<�*7\A���&�78��B�JD8�T�c	3Wm�l�����8P����t��>`���|��!@V�h_;ؾϵ�b�ÈJV������LFa⪸��J�����q�H�k�1V����v]"��]�m���";^"�(��i�P��>�R��=���A絉I�鸴����V~`���Ұ�\b��GLx����y*aS�H����g2QB���?WrcOy��}��c��<�JX)1A;�Y���Q���ɭ�Y�3����VP�V��*"U�T�y�=E�J��h}s
 X@ ���6I�.l�d�Ra�����J����<��؉�0�;�������R�$dE]��d���Ѿ��W�
��J�P	C�?�j����������sk�M��ʒ9�s�Q�|%f5C]�g@٪�l%��o~!�r۳�G�$t�� �3d�q��t�q� �Ƀ��~M�OZ�;k2��݋��	&�G9'~p��촤ux������rN�lU&W�b��n�*&Z��懶�;_i���-'"�P8z��_��<�(Dн-��C�pҀ���H��Ae��간?�=��r/�_̑�d��$D�ٗ ={��J�/�� BWH��\��qY�E]Ku%�J��_�鄨���f�_�RQ�+�4�k��`��r�ʞ�2��:��(Y���J��q25jkun��Y�@d��f�!�t�|��\ ����Y�0�2
�g��7�fi0S8�K���yq���c�\0_6�{z
��j��[�JE���v��w߲i^/)�H!�@6/ʾ��t\��]�L(��̱6�o�A�B�q���j]�?�o�����p���˓閰{Gke�a�۱3᠎+�Y��� �Q��%-��Ei%0��%�'�=5y��/i)|��@y�59�u�SJ�,�έr3�.F�$}e��}]wqݞ�F��x���5s�?G[��}5p��>��k4�vbQ�6h�U ��8*���|"�����K�ma��e;��CT���i�G��A�Ǭ��OS��zYP*�U۾���m�1&f)l��I����b��C=0�!�z�÷�u�EM��!2�b�JB>P2
B�nq�N�8s��3�<��c`��e�z�_!��| �	���?&��d(���d��������w��uJ~�D�L�=J�f+ ���[� �ݷ-��}|�P���/�\��3�Ds�P=a��T�@�)�Ƨ����+�^�fz�fy�T������8|{z��|g)_Z��uڀ��+!���hN���nF�A
���]8�.�8u���Q��X��O�3�X�YÅ�8s}j�����Vd�d��u���E;���3��f|W:S�۽�z�	[Ās:�]�z�A��>$��uJ�m?��1�f��o>u�.�?�Yb+���2
��N�i9]0��d�U�J���Q@\��wMZIc����Ħ��k����� %:I��}.i�����l��w����Ԟ=���c�)��K;�����'/�*w8��y�p[�c[�?�
����~U������Ө��?:��tS)�:��n@۴KY�f���QF�l��߶����5
Yt%�<qyW���(w���U�w'�Dk��j��U&�}���Q��4'����>7n@u*�o��屶�� ��n��^z-��̈́W�N�?Y����Cہ�3�������_,6�z�(n�4�l~��?�Bs�V��Ů��	�pu{Qdx+Å��`J�����藺7�}�:�y�]��E�����7C�w��+���>C�"�=Y�]֖���	���G�o��V��>��0^R�tatY��3��*k�8@%H�|u�
�o�?l{��R�*ڙ��v�Ig����a=ζ'��7s�`�K���+L[�t���Է ��K�Y�)�]������kL��^6X��a��9��
)�s-U��~B{�^��ʹJ]S�G_\��[-��f� V8���}�U}�<���� �k%"8�/�2����7"��fsK9M�k;Ks�I�X=�GZ���{UYwMXY-a���Uf/D���c��(��W���Z���4��o����꠽��+S{���zҤ�ҘH�JC����y͵�1��0K��^5ل,��,��pt=)֨hV�3^�߾-�r��{<�mo��{�5~��G@���7쎒���Qq�O���h�&͘�T������'�+y�&�z;�u�z��>�E\�(2VF��8Y12�$I2��O���nj�4t��-m6u�E�'5����{T'�Y��QJR��e�_��}��/N=q���^G�#v��`��?�kڱ'��B�|t�crGi
�5 ��FlbI��ɶN:��`�Z�7�h�җH[&|�E0��`q�P텋2��)1�2<�5M�`�LW�2�4L�+!WpzxJʻ�R����2�/]��+ȫQC�����ė���j��s�V��U7�@ۡ����b���^m��Z+���F�T��W"�I���i�s�(�oզ( �^l�#RK�ta�H�RcR�mj�F�����F�f�B�򲿓��ʫ��^t��z�?�AM�l�rў v`֠�,ђ�zQb^�,��@qo��,p1�z=@�.$%�L��u���@�	.c�p�=> ��b�M��CD�B�@������>(*�{4;��T�-���w����G�Gw��.��Z��J00���U<G%֩2=�d�r�N�KK�������<���r)l6+�:������g�p@�bo1�W�F���m�8�δ�C��1�
�0��C�}{Oy��ۥ,��;��O�
O�^
&$�غշKy?:�ijb��D�̽5�P���X���{ v�1Es��H��߾��;.諤��=>f���5���0����҈���/^��V|_�:/6�]�z�����jQ�_k���!C�.'V�#�P�O�>��Jl�3���`n+��j 3
��c
4k����/�PZ.��b����35���R�p�f�xڢ�ӺJ��o���ލ��`|v2_��a���Y�! �X��W:�#����F������������ɠOڵժ�q�;�:W�	�}��ȈR��?�����k���	YuV�?,�����"��ι>0���{���	j�D��5(P<�ǆ�:_� �B�� �uR���>�,�F�zPGW:L:"��075�֚�>Y8ah���&좘Lu����qs��L���2����-k�a������pXס5����f��mVHt������Q�leZw�;��Gj��oB-o%�wt7�Vhѽ���_'�"i�ʫ_13�
->_����=ǻ�G3�e�3����hԈ�]DD\�j��UԤ5������==E�(���H_���?��c9"/�#�vaĥ$���1��4���9���L���ǒ5����t%݅�9�#�Ɓ�\=v�1��Dw#�����.i�37{>�$����(Cm�B��*2��z�ڡI-����wpQf�/����x��d�ʢC�o��^��݁��/|3Q�I��^U�:,���:?��~I~b<�e��@�kG>4��ܴ�;�222�/�����U��?Uq5�| ��v����hnR��媒
#�z����P��j�P����=�ۮ}H��1�(���hM�L�1X�2~ixO�����ѽ-3�&��Y����]$�z�=����Y�ǂ��4��@CJ\�N��S�2��GaN�t�Z�j-G����P����r�ȉ�<���L��~VZŅ��0�=�M����u�67�Ǌ�L�6ݬZ��a���:^�3m�E)��M��+9:������Q�o+?8Xn[�!p���S��%��zVן���l=%�x�\q@�(ØqZ���Dw�x(G���v��i��tOgQ�F�q���2WN+E��\�?Ej��je��0�à�V�{��̸�fr�lG47��F��..�(2X��k�s4�j�hf��´/�%n�0�a�U�u�"|�OG����ò���>4!G#+���Z�=��+JbE�MB�vv�MM&�s�R���P����gh�U֩�K��U	/��>�ޥJ_ch�]fօik���n~n\qt�Z��E<O��*\���|=R�K~����6��޷#��{Q���?�'I�k,�N�Z�l�%*ٗ!������N3d���6�J�frN�/�Bt9��#
ա�%RE&相߷ZG),H�:��ȍP����Su�OH�G�(�����60��i��_���96Æ,��.����{K�h�Yu~���7�Z��l�a�ѐ��p~��r7I,�'�O�𜽩�����f������[�*F���ho�����c4(m��=�եB����:Q�/��6ם+�^�5�բ�x��;�J~ĭ,Ϟ�����В	�����u�=\V�2��j��:Μz3�}��Ј٠.�X|]o��yx����r)��6��A��R	�dNg�>e�r0�s4�#O�q񙚖���T���^tcHy(�2���'l�pO���W�-W���zthx)lE�&���5���J�e
�;�E�I��\G�)�"J�9��&�OGȸx����@�&w�Z���F���-�!�#��*O�q%2j�NÉ�����V���׌��I��#oA�RUB%�������D��P�����{��f��tI��v8E��2u���YT�Lf�]�x��MC�>C�[ŮXl=���яO����v�_g�&I�O�85b�M�ZY�w��V�S�;TUGc�"FF#���OƖ�!~�z��a��b$<~�N�T���xG��hg���!^�=�fLP}��,εW����D\���<#d��>����>��tKT�y���n,ڒ~k�8$� `;�����ItP����-X���lW�m�P�1Ři}�[�{p����+�$��M�r1�}|Td0�o�u�cLG�Ӌ8���*B���A��&)�o�K�����'	����j���ڱ4a���^��G]V�;��x��;9��ъ�\�����M��6ty��8�?J`C�S��^�9^ȂɺΓ�
��J���4Yk��<�R3�����a�־	-qP��C����V�&�ߓ��C�kQ�衒�d������w�8c�A����D̗NÝf7�������@���!lP��MϠ�޴��j���Q�������F��b�^�""�8݅-�qmw�R,�<\-�2'N��0�������d��)�a�U����N:��Y�ٗ���Y��9hf���v�`J4Q�C�_��\��y��6�E���ib��|�3��^�opn9�\�:����H�
es�7(5�CY��]]]��n��]���%��"彉O��7��`Z�{��ߑ/��۟qN	���Ū�qɣ�j���kY���y��r���8�f%Ƨ�u�tu�����p!��ަ]����e���jcQ���)oN3_92I��Lt�1�K���MF�~�hX�f����s�2�錺���]�(S��d@����2�4��l����`Kv��w����{���4�
�>��yN��Cn�����dd�#��ǀ�z�FK�	�Y( ;_��-�5H�·m_}�:�z��<V@��ʱj%�jsӬt8D��a"}���h�˧
db�a��G��GJv�j�����Ven����@��T�ZT;� &}ܙ�#���yV���i�d�4�~f��)��ϬKJ��h��kg�P�z���P�!3�&�� ����e���ݱ"U�Hu���)�\���Z�$���k�U�sC��@��^���b��l���¡m�Y�)3txW���+��Ɇ^�]���d�7�J������X��pT�\kN(�|�k�af�n��w����.Q���8c�M�k�r�+�O�EM~��
J
W���i;��x$��w�����ζ�]�^"��6r{0ˏP3.�Fsr|��л����e��T)z�k�/� �J5,-�ui�Y�h���Mr���Cr#�4����%�Ұ!�D�͇���\�(ʌ��Ȋj�D��?^�U�К�u�/tdN���#�z�Z =�Ή�1��ڢv�(^�̔}��k�K�h8<��|M�H�V�8��vSP�o����k���ӽ��ow���P�(Q��.wpQ������6?S�|�`�ٻ̞����Wd8D�*M2�&ŉ�� �X�$���_w�俗��*"�7�ܹq���������I	%�#]����G?���dA_yB%Ȯ��r�> �&��&%g�x;264��ө����à!C��A7�tv��D��-�
�=7�2�<u��Y��ְ禟3�(r	�%@6��Fc���ad�ݼ�����FA��ɀ��&�:`�(2c�i	%i�1��1�؟���& S��88��n��.�=_������6?�c�U=�`7�o�t����
<����N#!���)�� �4��d?z��qy����.:R�N�b��}�1{}���wѷ�W'�h
b��`�^S
��~�ꥄ��AUkߕ5��v1ʠ�`�V4g�<g��C�g���FIeU�fGs������H"4��0܉K��,�L��h�,����V�Z�,ʣ��2��?��FM�$&��N�L��_���F� *q�+�����S�qF��'����%����PZ!g鵣0��Y/�]B�DV����W�,= "n�f�vV����{�è�'�E⫯�)�7�U�D�7T6{�Ͻ�6�`�Vv�N���6�Q�N���2�J+��k�:�#H�2�y�y�ic��z0G%%��;:�//��1i�Es�gi�h���4x������@�G��yF�؟'����m�-���\��e�P�����
P�a݌G�����E�Y�ć���F�W�p�O`$��l$w��k4���?'���P�Z؆���yrW��������eSM>P�_����-�k~��=mr�����݋Qn����̶Nv�����}�u�Z�P�]Yj�x�w��0��"��-�b�o��O�r	
K*{9�7��K�ɡ�=wc�u�ރ��W�$����0*"mKO�n=���p�;rꚓ�2���ñXi6��/���ь;\��U�;�÷������x]�!z���6)B��,t�E{ý��(�'��kg�I7��<�����Ҏs[ԫ�䳫>^A�P���Ql�R��-��v���O�X14�S0_Ʊĵ����8��r�������tW����?�	P�q��N됕��{���|,�RF���q;֑����'�~U�ļ]Y�q��<@��#{aLC35.a`5��ͻ�|�fҼy��2c�d����>�Ү[����C@oy�ß����������'2�Ϯ�WS���B����$r��V��r��˔0>�+���-+��Gռ����A�р:e��/&��T���2��YN%;�h��=�b��C/"�]l�������'֒n��/�Rd��$e��O�/"6~Xl�WX���w�S���o�,E|����j� b�E�����V��o|xx�!tg�#��4�X��ɼ기�g���^���趴<���N���d�;$��D�E3�د�$�m���6E�=xi��}�qA�{���リ s)�>COp�*>��kҨy�f��$2�&o�������ѷ��Mgv�ō�owX<Z�/O�����u���R ����DH�I=�^��"��[Z��1�s�m��x�V�O�#,G���GmS�	�쑜ʪ�@U�g��9���q䆥IW!=Z�2]c�7�?�੨�"Zz�7gN���{	�GZ�1��ua���<����h�$���"����⎚��V�7x��zU�����b��K�2���P��x�YL��n��?��[��c�%x."Ծ��������a��nh��>��ȥ���<_d�����[c�#���/�E��Q����$��:� ��&4G�%�o����{1I
Š�⼩�ōD ��j�Œ��ɭ�~f�^�hgm_(���uykB�}������E��T|�gѳ�@6Y\�]dEC�Էq��MW2�^�m���e$�i�ɇt�s�,���o�S��UM��G�\��7IJf�|����Q�pحs�'-n�ey�Iz*���\�7�"��D����E��6�8�����H���^8�G�#��}���6iV�
��/wʁ�Y�'Hg ��z����5��<�,0���鸴q��j�^��q)�2 ���[L�<2�)�I���/W��A���Z�)�W�_ί�Ã�����r�QO�6F�U
H�d^��^�C^Eݦ�9
��i0��@%%6��a0)��/�r�6���m�]���Z��vc��+�$Հ��X�5Ϫ� ���r�����+�y�C�CT�{�H%I���s��{4�n����6�l��i;n����q�q�vje���;v����rO�FG��n�~9L�(?|nu�������O�l���u5�,��o~]�99=y� �T��-��%����C�u#B*�߫e��?��}�G����F����٥�|��*:wn(���C���Oh�B��n%���Lқ�'��y@i����M*�� ն=^e
��b}5� �,�c t2�6�ݍS�([B~�����)�J������<rUɡ�})� ��)��"1sA��vk"ì�~��K�����<��D��l��w��A�\�i��@i"�<I���$U< g�!g�L	��
?��Qu�8�I�9�&b��_X�ZyD"�j5�	ο�����4��̮�-[�,o��5��#Jd����Q"�e��yl�+�*|9Z�of���"D���!,xH���[��'��/6]�*W���C��D����֪�j)r�h�nw�g�4�I���"@��<��B��W^u�g�y~K��B���+�B�,~��y�� 	��Xi�D���nm'� �г��ib�X�� �Lؕ���<G)3��*V��z�r�a�z_u��vR����+�Qb�\��O�C�Ki>i���Q��l�\\*��/e�vy��0b'F8�G���N^��`��	P�U�pa}�0a��A"�M.���2��d�����lO���E+uD��).�1��� G�́��Zl�,�.���Ez��Q-o�T����X��.r��+^��=,��Z�~0��u]��N_aÃ���Aֶz��Svw��;hB�#I㔢a����?��1K+���G��v�|K���L!�G��jY�P#�&��c'�f̮��5:��+/������ߏ4��[߭���*f̆����s�J��]���h��	|-�K��4�z�	��Hro�x�*gy㽕�F�ށ=��{�����.|��]�ȼ�1�ٵ�#j���_��N�_~�v��i�ze����4�¤�2K��e#�;F/�j7-�TD	�b�\=���D�TQtſ{NX�i����%M�w6L4t���L��<�G�6�l�|!��*e���u�J��K��ՓL/V�ԋ�����q����-�{l�;���V/�r��X�Ԏ��k���P���10/mc�e�Z�nT�����=��F�rV��ML��D��h#\d��u�'G�Z����}U�d=ќM�y��Y�K�"��b�� �4���/�c���Y/)�Oc�״$�Zv~a���1ȣ`�1���� �b>A�;�l[���l�Z)r޵T�B�I>�9�(h����kG5;xǘ� B�7t/9xx�n�����=9(Ѥ_�C-�7��WÃ5�]����Q	�H3a<�5�a���_G|�����W_�V�ս}_�3/��侑_h����� �=�yc�ۺ��\=�ɘ�Z���,��RT����̳Ýzҋ���L��c�"��r��,m�̀�珮a�.�r<�W���{=����,��~�|T��R�ZBR����/�sz%���0��{�ȸ��.��v��5�\)G��|���-�v�{��'���%��UK�h�y�����4��^��P�-���j�u���C��>�?Oq��~q͝�}�n�[����J��/�sԱ��{ڄ���jTJc�^�,oU���O&�_q�?�'iN�-<���������;��j�:��h��f%�t��n�f�*����`	�-zG�3M֬��)]� �#>���?��^���PZsv�O܀��?�����l�2v���F�z/
f�����#�fE�.�q�+�%5���a�7�Iu'o<�����N�F�9�<�,�����FrZQ�C���kC�s�LM���4j�˵:8�n]�/p���(��t\��\;�\����Z4Ł�=0�1�l7�ȉ��7�j�J54��I���R�}`oy1�� rb��^cn��=�䢐�`��{?7t@�Q'����I���蒄����V�7�;�U��cr��B��t���	�O1%+�V/e�t��s�?���D*��\��]E�<
&Q����;f�c��7��(��YK�����^�ch�`jY2�S�R1���ƆJ�����g�����ށ_5/kjӱ�b�y���O��K�3�tj%���B��sg(q��o��7�n���O>X�d��LJ��)�ْȉ�)�T��x�"e6b�g�(��A:~?+��5�~�J6�}�3��f�Yb-B���\�����)��J�D���L�����#�B)=5���˲���8
׿}��{J%��E�&}愚\��eXW��R�c9�|�U��}��vݺ�p�����	�'����Jc��V��g[d�f��l���h�L�h��k���� ��eWٰ��z�(�a_�«���c_�Ce�Y��7�JK[P2���^+[z`vu�*<�0kv�3~����Ҭ�����j���� �&a% R�?.WG��C]����B}�s�~~3h]5�Q�A�EVYr��C��標������S��Al^_����@�����n�c9_EM�f�4�\�$�D�.��I\�m���4H��U��N-_e�:i4�`�b�h��E� >��^�:S��|���4v��_&QF�����!��S�j�9�V3�)CL�&������~.�G��5^���\��US�l���*���U	��J|?��0]�0]Bz�O�*{��;���P.T\��_R��Z�����#���T���7c�5�i.�4L��Ƌ<�4�"+)�S�TUm�Οb���i6���7;�i�6[���UD�z�sL��h��:B�;^�ׅ轀Cu��d
���K*aFܹ9���-�Nۑ�d�=vi�p��}���س�u10�Y��y�ud��׹���������4F�S]�[Ɏ�D[��࠹�\e���Rq�(Z!���\8�GS����X<ۨ�|0��3�q~��χ9��]��~H�:�N?O}�����%���5i@![�<��S)���:�����uV{p���^Q[���O~m>"��l�Mx�S~����g��`�U����&� �
r�g�W.�z;�_�z\��`��k������HF
��U�ؘMf�,��`��3>�5Br��e��3����,Np[�ѫj�k�̈��A���0+�F�-#4�57�$a�2�Wf{PD�v�mH�]Y��EAp98I�	}L�2����|����Mb� �'�q�և�Kᦈ��#����g��S�yz?����i�2����0�`]5�� JQ:�- �߃�ud��VF���?��G���`O��y�b|~ga�/e{V>���wl$Ug�M��z�W��5�.HCܰ�*���fޫYq�؄.q���o4�w�}�B���9�~�#3�[w�a�z�z�[���'ԝ;	W��I�R��:�
9�1J�9��p���S��1n���������fn�m�2�;+˾@���!��AP�~ޞV=��^/�/�~�=a�e����ݩ���9.K�9��f�/3��� g=Ϧ��s�ӛl��ce�Z��p�ڏ����/z�*��k�M����c��&��cS��T�n�7�L+�V^z�.x<t�|���I�n�<�Uia֛�>��ME�}�����E�q��TRW�w��Nt�ҽ_FRV�^X�5�rH���(E^hU���L�zt%B�t7�t�{07� ��Q��N5�tJbw��,�H��-
�k`�@Qަ�]�L8zwg#���K��P�����gr�65�\�Jyk0�$ڑ�I��#�=�fؘ��%^��9k��Cq��Oߡ`�H��wZ�Ay+��0]���_��xu׿��2�NQD��}|+�xrx��-NW�h�/�$�g~���)���5��̴�jz_6��dm�r��)�ձ�$��ҭ�R:dKBݨi�*�L2+�?j�����m����ݛ
�H�R�����HE�ۜ�ШI�K	��>��cڢ��G����aܺ��Fy[��m�Ҕv��e�ۯ�{f��3��h�q¡���~Ս�Y���Y3b�Oa��wH˻�LN�I���s�|��&R�"�d��Rx36(����n�30�X]Pؚ�SY>�l\�x��C�A]+�bF�>��٣�+^y�G3q7�a37��2Wܰ�<���=l�A��X箵j��H�gd�z�#i$���Z[y4s�|��t�T�l�k�~�����.V�Aٛ�V�w�D������U�&`��:[��^RTr�Y�It����T	�o ���������6��\8��B��ZQ��]3J���7�_���mW,�8\�ΊO�b8W�o~�E���
�돹"1N��T7e�͙+ϫ��q�V�����z��H.�{�[��E뛷&O���ŏY�`�ʀ�g#�8o���י��J��-@6`S)fS⤈��lE����A7Ua��U�mx/v��wIn�q'����Q���߁�-����M_�΀��[W�H*�j�76�)0'���lR��mk�nJ`O$��E�]�����յ�$'�^�;+�޷�:v��u��E����4Nj^�+I->���l��\�򾐡q>-�㕓��b6��}-��~P��Ƒ��dCn�\�\`T٫�j��;bo��M�ypW�r�/V*P�z�]b��4�?��?�%%V�J�[~Ww؊�I-#Q�~ӓ���3J���s"��1�	�M&�i����}�1�r�bG����VMF�ԇ<�i/a/���`�e�h�v��f�V��?�j���.�6q�O0�N�L�yxM�瀝.���gh8�p���he<(��|>��c2	�v~�=!�H���M�\��M��UE���L��=R=���������}��\ƢԿ&�Ɏ�Usj&ō���_s��9�F���'V�1`Ɗs��_�-�U��K�l��;̊[����Bm���<o�1�|bj''S���x��R,�]:��6���ߟuh�w�^�����C�b�$nc�aqP����\~����9��aԫE���_���@ƛ�zuW�C��T��*仂�{����Vep�a��!I�q���>��N��9�a=�+�@{cYw�T\���{3�>���2�A������A^Oֶ�h���̺�s�]B��]n^���wh�D�	EJ�v����.��]��
Z�X ���Ͷ6�+�����PW��;ty�w�C�:�5���x��dW�024�M_9�c��:�OO�����
�CA����`�2ńR�sN�'at"M�1�ٚ\�EV�^�B���@��)�rѪ�bS���'GQ^�9\-;\Ѩ^��z�<�N4�����sd����> ( �o�I�a���
-Jm�Sl��ՕV嘙��L8ӏɓ�읛���=i>|DmÏD��3Z�BW*���77 �˦���Mq���]�<�R��A�cbYe��������Ý5��,?�M���/#��FvM���$y_�2���x�L�|] �Ph������-w������n�o���enySX����g����W�.7HZfJ��_���I#_MN���9��ȶf�".U<6��P���XA�lp���ϗ{(ص�������=��sjƜ�Ѭ����l%b�x� ��� &��N�W����f���B�5᚜U�:�j�H 9����#����f�����gi�6�z{{./�Uy��5���/�λ@F��t[����qƹ�Y4���+V�Eݙ���{�gXf����e��~sFX��Fa{�A�̒%3�E�u��ͬ�{,�%Uv�3>?Y/�O��R�-���� r]X����Go5��^>4X��(�-I��� yp慯5m�x˥	!~���؃B��m���"y��_�kħ��R¾�d AX
����H�j�3ˌ���Gw!t[��/-nM=�����r���mPè�kKIێ�هo�:_(]�uujUO�Y������N�V�x~T��,�@ݠ��'�g�V(Y��=[�O��Y�# ��*5�]����ۜ4��^�P�Y������*{�Z���0�孠�>P߮w
���Y�4����uὸ&��̈�σZ~�� ����J"�5���7�سh'��ܤ{�wz�ջ@����+ɗ/������$�or/�z��s\��z�*a�����)?��[����2��s�β�^~J@'��\�E=��ګ���\�<S�&�2��nd���[:	/��_z����I*!7��Alޟ�q�W�ǔ��ĶW��y�?s�+ߙ��C����`�sCF���X��M��e���9�A�x���R⫸R�)`�6X	1���(�Ad@��yI3�}��)*9$]ت\
�mB��l�]jA� �_��=���QD�}���#.~i#���F�����C�M��˂]@�ڝ��o���+��59��F�Q����%�z��7�'��SL�.����@�q��,7�'�1�Yy�Њj�v��S#�E,��LBsL����?������P��셉,M��M�ks��c�4_`S�#Hi�s���ڙ�4��pdp��;�D�$OO�q�lsN��V1S���õ��3��r� %�Ɉ����w�j�?v�՗~&�G�a
�$a0z�P�EoБV:��mD@ �t�4�GM��<��#|���U��R��y��jl-2G	��"������ɴ�]|7m4�YJs��eER^��C]��F��-��"����.�?G�LT`{[j�?W��:1z�����w�(koT�s�e@�P����8��C >Cor�RG�O��ug�ݥ�R�F�-J�#4�.!��N5����fRp4�Z3I 	Dv���')Ƶ�PN��Eq�h��v�h~ɑ���l(Y��Qz���,������!�d����}Zh��ڈ����/��**�n�m"A"@����w��!�qiBp��֍[#	��Kph ��m���ݧ;�?�6�j՚5k�޽���^x�Aq��V7�H�����0����ҫ���↕�������hj��)���q�o�%qL�����NkU����o�CX�)��Z"$�j����V?�k�-z��33��w���?25S41;�^`����M=�ar�i ���|�i��W�J�r�/8���H��*x�^��/�+�U���lk�)�0�۬�}�ǣ;U�<+��O�Jt�0 ��r��Z�+���V�h�<~�K������
m:j.e���iJOw��1�� '�^M��Fh4ԋp�U�ׇ���t��)ד�&�BRN1<,{ej�g�)�{���I��@��k�V��.J�;'��i,	I鑫,%H�c��ybV��a��%qYs1{2{N^g�g7���������?�f��cY�������n�)��;�XM�k��L�y�Q�A�'����\_��:z�N~/��H��!j/��-gf�#��/��`A��⡘؏RO��i�%���F� O�ٻ̶C��y%��x�[A�´%{*;x�������x �t�Q*�8q���O��${��^�=�Hau�$"|gj��\�2�jP_@$k�ph�dD6	� ��{�[�	���x�Y=������+e\���{H���ԉH�l�h��R:yE�m�K��M�fEI�����I�G_�BD{e���֌�˧j����ƭl{�h���R����[F��
���2rO�N�Y�L��IS�^���m��
��IW��1�yw�Y��H�n�$�E4�~2G6]��P���){�� ��-�'}�n�%�?�ek���>2���t� ������6����蘃��2y��663yT�W`V`q7��"�ڮ+�P"Uŋ��V���U���tk�h$)0Ӎo_�V��ca�)�ᨥ��'�0��Nӊ T�z�^�� ��1�.�YG�?���.���>�lt=�P�k�<������w�6�6U�6ӭħ�6z��i���T���tL�W�F��Z��b?۩�2�3�^�9�r�P���щ���~/?�fV�d��� z#;��b�������T��םc%a�ؠ�aͺt���iM��6�E��!{['Dƀ}�������7%��H�t��b�{�~�k��K��X$t�^h:��n%]9�e�f�b�7ظ~["eUw3�T���+O*w��߰�E
�^��dP�c<m�r�����E�v9!��������P�L�G
<o�O��SY(�����G�gM]�j�̤�4�W~��$���$�ؙG��-�5��Ʋ ����aG� 蚥��x�@ma:~�`�m��9F����iEg���$k��a�Dcx%�^�:~�J�#�ʯ�y��R���Dq9�ok_�H��Qo����2�9��յvc�BA����uq���jpt���a�9D�N҉'�XCk���ߺ
�AX���&a_q44G�
	��[X$��{�ᄳ@��)]��ݹ��=k�'������Ց:0�w�����5ABq]�F��s� ��-�����H"ЈN�����?|L�����#�5��������L|.���6^��X�WP2��s��Ja�s=X�~�k����h5�YM)g����=�?�S�*���;@�4�^ؒx�E�(/�ov��W)Ĥ�/}�8�l�f�k��O�g�-4k��u����گ�px=�ȩ\_t��]�<���5 &񆯍�VD���)h�jl2���=��qU�AZ)5���o�'���n�&��aT9N�����d5��e�5�׆�;�U�Zy�D�Ap����b2��=��_Y�Z ��i��t�I��h
)� �[�L�v���(��p��GS��Fz��c���0pb4+���~�#���rP�ґI��5bDC���H�����ϯ�YG�
w �uj��zd�Ӽ��t����3N�.��_d"n��]	]�lq{�67��4aR��#{���^�;Y�T��	��U)�;�v+�d�aE0ĨV�eV�Q�l'�0}e��8OK�`��f5�j��ā���Z�)k
��eqz�
":2�����g�#�1���~�	�A�@ƞ��T�F����,����Y�KeсZ�|!��U��@�ɕ�m�ϑ������B����� A҈��pU������	˵"��M���s�����\Ue׊�^(�I\zQ�1�&RC^�P���o��ne��o%��J�9nG�ˎ8�1��,���J?m��u6��>��}��>��SW��,Re������PdpY
���JqA�ϤV�_� ,Q�N��맩|v2�m�~�u9���٥�.�̉gv���t�;�=y:��w�ٌ1�$�˰��T�Kw(+*B���4�q
rI�$�Z&��Ƴ!7Sڡ�Ɩ؃��~��'�L_^M��6Xŭ�
������-ر��]����k����>(l��e�jؑn��_I6��������q�Qb�Zk^�/XXN
�$�).XUn}3���4jYC->dd5_�d���Ԙ�NY�\8������U��L`l-\����2�*6wg��t2I�fy^�fk�ֲh�3CS�u��+�C���Ga�Y!�zi���� ���ZlU�	�s�8�o���n��7��OZ�`X�]�J"6��g�ٔ]N
��E�s�1���W�q���%#ӓ �##v-�6�f���7A3��7G7շ1�:4��O�w�Ɠ�G䱴x���mF��CB�o_r��F�<���U��u:Q���}EM�@�V�ȃ�@��#���<] e����N;Y�7Q�pDlc�o#��P[!�|��E���i�V��]��ө8i�p�{����-�N����\-N�E�M)�$���#����+��g
�tٹ�m��i�?�������+�1�\��a�1�|y+�o�V'�,����$ھ�\L'~Ak,Cd'YEa>�a"ufb�DO�n��$� �M�f��Ԣ3�{vP��Y��Ed$j��UsU��W�*�6{����r�\��Wq×��S�R��:����Kx����q�:�n�BG3?�(LR�zQ�A�h`�����T;]h��It.�볖
��3ͧ\Q�ⱵMW6Rj� ��02�����A׀�
��/acFX�R�`��ǅ��ACxo����8\(��2�q�U�ջzh�O��E��Q�Z,C7�4҈+���uM��e��	� �a�ĤYQ�-�Q�nsy6�Ȯ�b��$������l�}�9{2��\�C�i!��O�u<rI�걡��tC�}��,!UyC�rܲ7���~{󶱶��,&"�K���<�>�M��&��U�Oe�?)�,�
���+�?�@��T椔�|�IQ)9�+s=�����GbdJQ/���]��V�fv�e�O�ٖ��
�r�w�/�?�>����CVh����!&W�J�ce����N�,&7Y��������d�$V�ѳ��^��J�*������ ��;�j���_�7�G�<�ڙ�/�'�Jy���c�RÅ�?o��M��ޑ���A��Yо�u�Z��m6��BS�F.��&���>�����'l�m����l�z��^�K�U����a��h��V88]�q(�)jɹ��G	�9e�E� )m6N������pLv�5���ncv@{u����k�A���D�T�ں��?"1�L��xFR�5c����t��ϱ9�X���v�7Qz����yZh�5B#p�[6/�������rw��>�]�IӅ`~e���^��v����E��O�E�Hw���*M�?����'?��T����������?���L?=����5� w��$��Z0콴����&���hx��^�ȎA\��vq_�w��Y,�\<��p��/��6�6�9a#&Տ����7(����L�9$jv!�/I3��g+�xǕ&���w v'�OJ�]l��^4H6O��v�k�F�t+sv�#���}�����v��L�d�P���0r��e������X�9l�S��jdy�V�P�bL�t�aWJ	��m??��?0�aD5\"F��jB�����|�����]M�ѕr�l�o��Lʊ�j\ܟ�*���
C��z�+ѵ�úezҫF4��H�s;uj<OiV�����8F
���T��/f/��f ��̝}����G�+-��C�	���������f���N��u���|�G�8��C��cP5�	Y+��S�wZ�*l���R
����@>�*���(d��j�V���ѭ��v[�{������7��<���IL�q�;�U\5u]%�&�m�c��N��|�W]�������r�x�m����z�d��/��|?�xY\ٚ�x��~�[jq���2��g���`�������ķ��$�s�L2?Q��*SO+��C㷞n�U�� !&�:������t� ӹ�Q��M�f靃`�O�Ċ��E-h�4��X%+�A��ZHkl�|��^�:�`�%�t�����
,"�?*������]���'���2��g�����D�>]F �$���n��%�af8Ǐ���FŧF��D�	���2���O��34W�4Oz�L���H��I�����^׉Z���l�d��L�&b���l�Iv|e������Z�����i�+÷&��L��VD��#��Q���N;)kX�`)��8]��>n))K|�p�y>CRj{�ؐ��Z�vN�N���Jx�I������*��=i�g�&��t51�R�d�Ƈ<0�-:d���;�v�^�q�ז�.���i޼�5��tZY�MdB~��mBW%c�r\;^;�/yoV63	���"5=a�~�$q����-)�/s[l�SP�U�?4Լ �C��
 ŋ9�>���Im-�b���$��/��rZ#O^�0t��ڊ�W��7���ӛ���X�|g��X���`�`:��K�✢/f���J*����;� �蚔M���O-���'f_6���g�*��N����{M�����2愵���C�3cy$b����1�Z�p�e�W���G<�L0���Y���k��?9Sn��T�%,m�����|���k)�!�[F�:���*í�h5��Y#0�C��a)����A��ϳ �k-���.U��^�k�z"�>��N�2_�kEM�q�N���Ѓ���Tnc�����I���y�\����쿫!&����"��F�j���}3��4]O��b� \q�����6_�qԷH��N�t������5���a�̘�,��	���%��o�X/�&�n��;���e�Lt!���W�O���k�q��S��R����j!wl���@)|�R!1��4Eli���J���D��&Np��1lf�5������q��+[���ޤ�����c���M�R9PpU�^~���Ӷ�>+���8��־���򠾏�skq�r�j3�rU�խ�Z�e�����o�*�M9�N3��%������;��ϹT���/��Un~;0)�	��捘c� ���̝e�l��t�I�D��
���>��#��������>�gUt��-�EqqWUI��e<�l����$�4ע#�q�g:f����Z	�й�����_��Ұ����I�ci_�t0	�m���d�`����IB|��)�߲��a)M�*����F��F��ӻ�ʾ@-�8�$�s���T!��s��f��di�K��,���gv��JPk��	�z�ay�V����v�Yi�5����c]+��?8/,(�K␛����b~=Av_�o�jEv��Z�����N	C| �Z$^Μ0F�Tr�t����j���f`�ӞQ�پ�"�!�b�3o7d�Q�ťF԰f3��2)�I@�0��#���L&�v����Q�М$�V�>�-���ȵ��x����o��5���<u?�y63|+����:V�M���,k
�|�� �56��I����d��I���GQu�o���M RU׌r�����G��հ����A��z�O��G�2ۇ�C���q���Σl�s��A`���{q�`�z�(�W��C�W��� ����4H����h�a����~�'{U����CQ'�^ &-d�,vy�	V�Pq����2w�`�f��R���������,O��nj��9O]�db�j��[���}8��N	���gbS��W̦��ӊnAq�Y���!�lM�i�f�3ȥL��.s�yfF�&?Hm�2��*�kCǻKT��F�R(ú-bǈ�`����c{����& d����%/ �1��3h�n�˽�Ku�6�i���j�c�ȌB�{����x^��i���$�����g�/�f�깤��+��J�V��-/~p��]��Q��͕tԊ��<�ˬ-�~Xv����y���\��[u��x��<JX��dB�hX����y����~ -�(R�j$WT�Rh���^�������p/��(�䜹q �+���Q��l��^�3wO#���NQ����N��g�9OSщ���Ņ@����L�a�U#i�i�n�G��;j�Уŋ��p�t��#1
�����}����$��;A(>L�(����7�iVR�N�!����d�t�V5q]���<�JD���z!�y��� ߥ�k�Q��n����I�EME,��{�v�DVK��I����rZ����Sd�u�Ӊ�I�.�*��M�B(�������,�d�oV����Q�OL�2�|VէØ܉#�G��D��Fr��;+\���W�3��������4��蚭����V\���u���K���+]|m�P� �Bw��H9�\s������wl�l�z���� ���8��x@�w�����`��𕼼(#���o��	��L�=�7SM�'�;�'�e4��CJ�&E4�}�g_dOB��~Q�5ʖ�Rl���bSy�61c5��a$wIkԎ��]��h@_zK���:��l��G��_s�+�-*�3�x��,'iemH��	#VH��Ɠ���]f!���� <l��I�;^��BQ�G�^񕃳�E�T�p8|v�����Ԇ����S��#(����G�t]:
���3�~ d?����D�Q�g"�@2}�Q"n7�Re^�$f���*�HZ:��*N2�c�6�چ�-�)�&�������{$�I%|Ɉ�!Z�i�є_셜b�)��^cy2��V022ʛ�M�@xV�H##��Uf.��'���\9�g�ȟ|�?=��K�q�/��v�҅����L�-�+�����g�NHQ�������4�`tި����Q��%��3�مH:���B�YyҷH=����q��/��S�U������v�$�5c�3��H��z����|�� ������)������AX��C��t�=��be^���YO��#)h�F���DL�XL�JL<jǮ��B����+�dٷ�G����q\��k���ʔ�ي�:_���K{|�����_�W��?A��7 �`�d��t�}��7T-4Ҭ��$4a�yTb&@�d�X3w�S���<�5�ٱ�z.->}1!���ugd�|Y��a�V#uʰA3��hSk�"�t'�=p��j���{����y�U�l�����2	'4VJ�FvEs�H�(�!�cna�!%�ٖ;d	7rK��X7��M���0S��ST�<�"lI���/K�f��`���$��d���P��)�>:6s,/�����(��!h=��*H���ōQS��<�7�AJ �?��=����X)E(�d���S!��u����o���r�d��wf��Q�����1���˺�]9d&'7>�E[
��P\��M��ˣ����d���ܗV�z��4��'���m���� mɄ`�~l,!K�vxY�:+�B�r=l� LfZS['kh������i��&���,���f��o&{w�%��
������#=��T����xW����\\\��(����U0Ր��x�G�=JZ��k
6�㪙)Ze�z��^��2��L������vQ�<sgm%Ʃ���J��@�e�ӂ�u8�ܳ	�J�m6>4��B��&F7�tS�r,�=#�l��~G�U�(�Y�,"�0�Q9q1��ux2w���*Z�D!3R�ٸ6�`
]���ZH�.�BS�>�3d�9�����2\iV�}L�%�aI5׋?����E�|_�yp��O]2F�����4�P���-u1���Y�=Y�w5�˃Py����� 6e@�⊊�U;&���u��DZ5�]��N?��*�ő8�Zm�p��J�
�g��9��[6&�O�"���������_u�à��[K x1��ln^�K� ��c�r1 �I\]]Ǉ�IӇ�����c�3 �LO1�e��k?��.�!
kf��eg7�I�XQ�=Kԉ2bbud�>��_̋���؄}�ߡ&�*jE�7s�E�����HN� �����K��h��y��P �.'�#Z��εH[��_��`��H�?!�&���qy[�:ou4�S��@,QwQ"�n�@*�Į�H�N�:��#5���A6>��	&@�y�b��w�E߻�E�P�~*��X=�r�c�>̠:�gѝ�������e�,�w���uD���_��q'�FT�U&"���VN�DEe��+O�j@�z�tv�vv�в�Q�v�q���㣔�xת�4�
 �R�Jr.��������L��)L#!U���D���ie³�,@4d�H���(F�赪�ccS��ó��#�~z���ѱ��^#55�bv7�	�i�~|���� �᮫�\LlP�t"%��k�9 ,����F����-�#4$k�n����e��x�q�&q��{�5O�N^o.?���e��`��伨x�U"kd�ũ	�426���
�� �r8����]�EL��w�R�͢�l'� j|��E��R������ʲI�"j�O0��7[�E�O$vw�^��m��0���:1<���)� ������ˎ�n��8�<@��Ȕ�����O�ɟ����^��s7���Ij֮G���k��pJ���2�G��Cwݼ�K�.W��a6&�<̔���\][۷�������@������9ܞ;�1��^�}��9>�*:�j~��	ps1N�$և6K��Le#��q
�P�q����G'6���μ��ݟ���3m8�[�H�;:9�-ې_cR��=���/K�n��BT��Y몉���De�����{�?�[�OvX;6:�6�g6�������,�Ʋ:_q� N��`��c�ϧ���� �~�H�19�Z]]M�ֻr@�z���&�T�C��PS�.�׽h����/����\�x��Ws��u�]b���s�%�-{evG�.�E\��G<Q�0�u�j[[[H0�?��B=[x:���w�l�8J���\��Ռ!O�"��HC��|K���M�`l��	���3^�d!��f���,�&e}�� |�Yq��MJ���2 � �Q
w36��� ���.OcT�����4>I�+���"#���}T�m��lƯ�a"�P���Z��" #B���+2�	�Q'}!���JKK[�/n<+� Կ#W��V{]��;�;�a��UWAd?����+�]D*��(���_��oH��KBB��������Xo�_c5_��_�~er��]V�f���ӹKR�����A�l=�����5֭� ����}�Sq�lv<�h��3��oiw]bF^���1�+c 3@v�[Ɠg��Ts�!�ܴ#ط�/?��G.�Q{��^�x��0�'8Zp��8�BT&'�����o��R���Lxg��2��^�ɻ���]jFF��go�P?�~��Wb��zB�Q����Q�F�%a��=�q��h%&�PE+C	&�#�/5Gr� ��Z�!ݓw�ײ� ��'�eC�����]�B�u��w����G(����kȨ���mE�a�xl����m�+����L��D���xGX��[lh�gס�a��W�����E"~�>ܑG�*�z����C�&[�,�b��SCL��;�nmL�~���"�Ra?ŧ��p�0K��|_�"�
ʭ+n��?:�ffl�]��B�,;6��+�+ZC|��5����O|*m�_�k�w���Z����AC�!��>1QD�Zu��Q$iL�t�;@�i��jH]�""O�N�u�ߦn�D� ��d���&�@@�m����p�)�w<�_��~���ˣ��{��=�HM􉞙��v�8ߙ�M��tr\Q�(W�oEf�̴��M�݊�Z��Q�0C�
m���m�)9K;�9���Z�x����>u:q�*������b��R{vΜ�d���j5i�鰙�sv�B�I^�_ʪ�|�x�#����^�+Kg��O�Pc���^���~�R����m�ju�!���6������r���Q6[\xj�B���?���ݥ��q�~I��/�s�Hͯ��%m����
>�ͣy<ƶ��)�D�P���#H�aQ!˩J������O����QquQ{���ަ��v���d%�Z�c)�ع0.����D���sny�EW#�.�n.γ�[�^�_�D�nl���{i.6�*h�j謯��mH�_?��i�G�-`��pc�,�ć_p�x�\�*�.��^_�s�h���͑䖇w��Ȫ�}��UhBaD�z���=���"ڕ[
0���Й+�JS�\K����S���� ���+|�}ԖYm�_�^�e?{�s-ֽ��_����P]Yb�2��替�[�fN_ub翽
�:�5���+|$�V��y9�y3��]?�t���x���{f��	�e�	eU�R
�Χ��*B��_3vv9����a����-:c���8�ոO�V���aڒ8Ƿ����R�~�� R��fr������!��#�7Q��D������	�{�ё�{��k�Zy�;��g�TN{=�RKr��@�1)y�9��H�P��2����X8�����B�C�p���R� �N9m#k+������?�z�^�O ~�)[�3y�(G����O��)�%(��!�FU�H'�Ae>�5���a���g=$����ѣ��;��Y�<�f�P� >��V�x�+7����{�r�琞n"�l�]ڳ���j��<w��.ێ3`)Ĩ���&�z�H��{��Cp�&���m��Un�&;��Ȳ�&8F(�o�s%jp�O%�$�y�h��ŀ�/���(���l`�������3�vHL������(C�տ�}xge��<Wڵ�Km@�Ho�O�S2x3g��#o|�^l�`�v,�HxVT�k���2�Q�+��n� �ߔvB+w���^_��^o&K瀓`H'Ď�>D�t��>�2\$?P��:�Hg�L�7ѫN2ȝ'���,��t��H�/,?=h舓�蘽�������z�^�H/T��oO���Ǥ��J�g�lnV�ޜ9@���Q����|�	�0Yʷ)�\�J)
���&g�S����q�>f�:��G�2����76�?-�f:��o�>EG���l�!Q��og.Mȕc�}ϩ��MO���T6�]1�s��C�����%����|��wT�1�o����J9/@|�=���8G�#�D^k������BG�jC�M:�<\$j�M�`M�,6�I�k�R���	��rF���n/Q��_\���5��hŏ�5�G�VHb��x��{��k�j�caIޅ�M����H#e��kXv�򘑽��̾����~���UGQ�>���=3fkT�~o[�C}�:��H@���E��!�>����K����l.�+[��Pd	6�Ȑ�����U�F|��ٽ,��_��Z/�B��ьy�����Y�z�mĴ �ȫ�7�5�5á�!�����B�H��M_z����7Xj͆(BK��RJP��䊏r�afK|�]�=�ϱ)̜+�ܧ��;�C:���M'����X&*�M�Z����d����D�����{�%��Һ2�Xt����^�p�s��\7�)֑��k�X�A�Z�W{��t�����k^A*�ӡ	����5��v�z��ԍ�i&�?�#6�����_��+P$:�g5��c�ߓ�iV~A=��Q�fv�ɷ�r�M	���yJ��vS�)b֧g/�\�3Al ��sn�9��_tm»-Q�{Vi�z�7TŘ��ݜ]�&���:]l/�&���-?M��E�'�P�7����	�-�>=��MG���~�J�k�����8�����಺/�3��� i�.<;,cP��9\��1߯�E;���kO�����Xb%�!�/SL9����#�qh������:���P�����Hk��63xQ)"�m0*G��r�PI�����x�Y�}�<��fr�����'�1d6�̂3B�{X_��밃n+���d���e���e��U�V��E̟�Th�%��C�����XoQj�7gdGb�D���Qi����<Yf��nJ-�|�Cj�C�u�LW�^E�'K�[�W�N�����}j�+}f��{��Tz��F�p�N�=���6���!y�>D�o��'�2}�x[��=*�'[�2Q���o�&�~5��6�n�%Wwf4�ߎsÊ��0`~,�C�Z�_��M�����ǝ�$r�O��ި�f�Ìq�>�dNԦ*�����3�'����QG[z����fF��w���4F�������
�p�K_/BU;]�	䕭_xX��F�Mӫy��an���GD�+� ���Lq~;7�M��6|vr����-|l"5�����]�w"��BP1��kY�g��l��{l��F�����z��^�s͈duW���+�إ�1��$Ts�bj�$�ϭm}F3��H_�N�uݬl�̯ ��˽d��&'Mʧ4�=*����:���t��w� �<o���M���빏$��Ԯ{�K�K�E;Q}�]
�V�����q��rk@�蛖���g��?*vsi��a������S;H`�hO^O��Ĳ[pi1����+�(�;m�����P��g}P�	0��p�:��B�1��|P��M�W�ʲ�:1����8��tJ#-����b�R:�Owt�G��u� ݔ+�J 9���VX��-h=���;�_R`�R���I�j�O���P�v�� 6I�*Sj�N}��S��+&�+?/�1���l��)LiECo�;�{�l����Pt����I��U����� Eo����͇��F������Op���"J���]$�������f��a�M}�BX�#��y�+�ܴC��#��$j��^Nݩ�>.�Sv9�v��2�d�\�0�"�~��[Vc:�4��Wn�=�l��+w��iv�W;j��H��5������Ox%['��ve��w.��lp8�A^�~W��G�2�c�)���q0��v��ߎ����tff>���~L����|$����7��Q̢��MM�鼍������٠\�_Ax~����O����e�u��]}hr���PbΛui�ԧ���I�y1��*��lΆ�LհK���qT���p7~.\s�2���U|�YC&ؕw3R^� ��P���$��u��N*����O��tXX�F��ҥ���oI�L�S�e�&��R��p���<��f���.�3��#�-E	��!�>X���}�r�l%Z��%�*��j>?����?6����y�$�F�߹������t)i�-O#*�����$���-d��qo�������7��E,'�Gq���4��ﴻ�BW��W�\�iϗ��*\^�c$w}YT6�C��b���hm�P��t;� �]�Q�}5���0�M�q��8i%Va�r�G�W�� ����iK�k�U�r����woTcn��B:�c�m���
�dS�o�R��i�#�0�7|#�j
�%W&�)3��9</�Rd�VA�6�N��jJ(q�$&
t��q=tQ2ti�u��}��g�g(���ص����j�h(�}��K0L��a*��W#�I��D|뷁�h�W����sB���M�0/��ߟ!�Ba���㝔9��>ؗ���߷`�n��أ�jᝌCgbɟ�v�o��Ԫ[;ߠ���M�::���b>0���.ޞ�E�3k���ky��S�`�R`}m�y�&Z}cC7��@���|��3�h����ޫ&����:>ϋM�qR�6#KV�jy-F��[S��Dr�֯��ވ0�6�6>�ʻ��E.���5�(���_��op������6S�:3%
�y�F�&�Ǎ-�9��ۇ���N��Yɮ���IF�9C�d�@ݩ��j��it��ϒ�Ϻ�+�!VI���Q�Xj<	�HH,����ɲ&| 90��ӵDQ~6\�	�^/��V�WE�NZ7h�c"����PK\��j@�n)�"S�%�:bٕ'x�?;�,P"��;�$�7�b��ZHI��h�_�K3���O�|�e���
3������M�aZq������j\3�3�F�i���w�R�����0�9�����^�;���!iJф٪��n��o�7�B��O�גB{���|+g/꥟QK� \eO������`b�zLg2�/��2_�����u�H(�~� �k������~q���je���q��/�,�%��|���P8q)��)�(��r&���]����刐1��ܷ�q�kq�s��)#��\�rXn�r��M�T{�W�<���2�˿�P�7M���A�%;����U���Ւ^ ���'�Ǯ�����&]T*��_LX�)�B��;bp��b�S����aVm�I�Z7W#O6ϸ$���"c��F*}S�������� 5}*Q�WH�m`AYa:���7��7���*"A���Q�u];P+F���t���M��'H��dr&*�h��Ѕ���Q�ϭ9��P�=زm�K�%�.)/WT<>�o�u�n�v�ة�)��ԕ�0�&��5$��ۓj�����m�w{g7Mg�~��޿J���w5���аfmW���`�h��w��ƳVo��mۖd{�|4�U�3�9I�F�إ���= 2���S�^Ǔ)�b���H�`�:�����!Gu�&�Pչ�7G>XD���.��V�m�r���~⨔����s���'�|P�3�d ��.(�~��<j�7cx
Tj\}�J�N�"��Q��h-
u^a���|��e�'�D�4�Ì�$�MR�=7e_��guv#v]#(�J}C�����<�f�v���6U���I~�CyN��,��ϕ}B��6�Z>� ?����f��J����UT�3:H#Z��\q����$�����Ӕ̓؈u��57;�q8�T*1��z9]-�������p��F�@ؑ�������+�𶢭���@��蕊a���pe���'g�@"���1�],�Y.��R6P���c/��bs$��8vx^Y*۔蠵#����6u��vbAC]#E�	�%.>j7M4�R���t~Pz~ҽ�%v��M�[Y�c>�p�F�Jv����7�F�	҂~�&��o��k()ړ�����4�*Q�zh��F�����'�޳���T��ۂ�I��8���w���`�[�a��0�>�PJ�O�����nyM�f�qa�ja2׍���$���2^�����/ŵPl���1��&8v��G��8���:��K��o�tP!,!a\�l�����~=>H�"/tu�p���>���յ�p^�:R?��YpD{�8�Y�O���yw���!z{�nͩF|n5�����q����Y���}>�cwӚ?��L�]NO>ʼ�SZjJ�#�?�U5�}][VQ�S�r+����.��� �O��kA�A⥐�S�ع0�:*#ܦ�d�v�n+�Eٗ���=�=5p��t<��Z��ީsyx>�6��!�ߪ�O&�z�poyK ����9���w�,!t��{d��ek���i��;�|����ml�l��TP`�":�4�{��S���+���֫۫!b��p��e��"3ݤ��x����Y�ҹ*y7K�kG�{���dW�R����}�R&�-�[�E֢k���5����]��rk#��H�=��UQ��̀5H���}6�w��`�Zes`����ƮA���G�H�8��UE�'��3HB'�Ѥb�+�X��~��Nҩ�K�����dX������3"T���; ������{D0m��e0'*��llq��Zi7�*����8p�V�i��g!/�e޻�e��nrٽN!84!�Զ���A�%_�O�E��mP�ؚ���O�����8k3I���Z�u��Ē"��)�n8��̈@\���|__�ā��}��(��~�"�K�����*~��!��eԴ�s�8�ҟ ,#�K�x����O2�j����U#��6���+�R�N���o���Dk��081�K���ǈ�݊ �0��Bo���4�	,�^�ͮ���h�!��a���h
��jM�a��ظ~��u:�-ي"������q���-x�!�U��gR���>��-��Z:u�-~d�<T��p(ǭ|u�s�Q��L���=�̘��g܌�|��)�j̐�|�wM�������q������@�X�|�L�Q��#U��A�1O�8�{�u�v��B)S�L-釮��~Vd_�4u��x�q�5�+�}\��o"���z']ա2�?���_7w-Lwe(�"�����kN�zW
�|����K�@˙�I��� �v��z�T���lu*�e��xY�;���X
ZS�E�y�����Aq��m#��=��3��9]�NSs�s^�1��m/�p�s޼�����ԁg��Q:.���Z̹XE{[�Ƥ�~�ߺⷃ�-8�vN1�/�� 3����Ί@iR��K�����[p��,m�,�w� ��=����kp�w�������n��Ν��?�o}k%!lf�U�U�Uݻ�;䯙O[�-�R����D��ͽ��w��Β��vr"�pZ�T^BY2�� ���,̴-��QɬN!�]���GJ�^��Fd�* �_8�$���/��i>zJ�z���DJOIB�hd�V�[~nU��4�w��tg���&��"�8<���hO��p1�?Y����ݪ�d����}��$s%*��V{�y�φm�P?��<�@�4x���A����� R��fy��Tu�fcɺ	�����۰�#���2򡏽��i+���Ų<�Yy^LZ�~�]n[�Ȝ8�L/��|�v�Q�
k�4f֣r�L�����| �H ��}Q�Y���,��1�-�w��]˹��q�mw�`����-��#D��2j}IatzY��,���OR��;��'*��(HY��Q�@�i�v�P��d��K@3֙�9Պ�AF�����c��Yڿg�0U9��w}Z�2�Զ"�cP�	�H��z�`�$���F��΢p���{�bF2HJ�����Ns(|R'8��.��e����;����ル��*}�9��n�\e��D�Y�U�}_�h}A ^���ӭ�@C�`�ǵ���l$���q�o%z�yvE������e��L@u��ёJ}��$0I� �f0��vM���b�Tѫ�9���Ϳ�ܻ�gU���᧱�?�5=��4e�7O<�� �9Fl���R�5��w�����)ߘ~��ㆉ�U�k6u�('װ�I�MW0�6)�,�k��u�"��F?�6$s�2>�ɶ�%��j/``S��{y�g:�u����i��醞W��WG��o��DW���6�]�G(ZH�s����C��6�����8�#k��c��7�^�d#?-�`�|�5z��/�����#<n8{u�2�B'���E�iP ���y�ӆ�y���J��z�>``��h&�	��'<��8j�SZ3����U�5�Zn�@pd	�9	nk.�I��:WYS>cvK�]�S0�ճ���|	�/DDf>�-�l���>�|��0��l��]��3��|�BݢbLzZe~��%(�f��(��#�1�������NT����L+@iYD�@7��Z�o yp�N���+������^����x�b�'���-n����S��g�;��[�$��O��I
6~#�A!��Ø�Xd�_�1�����bΡ��v�G��3,U�]��`5ܙs�կ�4G�w����5���F,�){�H��٬��ܳ���� %����;8۝�S@�n�ۂ���gKRs1����.�S����k�������M��m�y�Nj�scX� �o�&�U�NJ�����I s�!�vΥ�������ދ8�z49,��[�7���M���qя�v�z���b�������=���jE��R������@����W����<�*��<��G�����;�V�m節����ӫΥ�m+�����/�����A�v���`6k����W�k4���*1LyUO��M�H��w�|d�`����>8+���rE���_L}�C�1`�j�Zc2�]]�f��D����H��%�����"�^EU�Ȍ@�������ʯ�k��瞜/���6��P�`�F�~'@jŸ��;T�r�L��$R�l?3�z�N/��b�"����*q����ݠ��U"U��ǔu9ڰS���3�a�T��e�)�7P\�b��PY�Ua8�9��g���vV:0W`�Գ��R���dGH9 �X�v;��2���z�y�|A�����ELb���tJP�w�7�QME�����O��=o�ݞ�x�,�iv����6�ԕ���h��tn#���C��ͽq���S����FVD������^1����¼���ŵ�I�7ƅ�d~�ΑzIDeH_q����k���~����Z���)�l��"�!l!��	��(O-�&9��!aq�I��PJG�<}�E�����0pn��5��R��P��o0��T3"�����M=O�S�q�<-םO;?+^�C?ջ�� h�	H#CLm=%�kx�ӘP�?߁�+����wm����g�	Ӑ2�JF��gb<��D����������Fz	�'��0�����l(4{��0��}��;ߘf[3��#g_�c G���+��Np̤=�ZQTX�U���_����5�ӌ������f習~��pW�uA��z��s�e!��%(����@7_ F��A#��s1�߷#���":-���zV[Ĩμ0�}!ǱC$�"�D����ȹe��N�p������K��O�>���pY�yC#I?;I�[����f���4U��V�xZ�-��a-��a}������{r���{�]6�y��0��/���A�3����B��K�_���ϫ��nz�!�T9ZO����n�MD����D۽���6�S�K���H�X����a���OEx�[-�G*,�w�[���I�������QZ�Cw��F�9gۃ��A�E�Z��E�0_���
	d��ѫ�[�V '���/΋��3�jQկ�8`@U\{K3��>ȫ����!�4C��N�7�a�i,��+���8Wȑ��H/��.I8��mp���c����Z��Sj�v���{ij��0�
3���/��Ѕ�bN�_Q�!r�*�N�(CE k��Kr%�.�_H@Nd������#����d��;�
Lc�c2���!�i�:%c<���Br �U��#��CY��>�w���c�L�(��~��|�a��y 'dF~?��-���1̙�=���y�`�q���,t��,~�J}�`̸A��F�Y�{Z&���%�9�OXxY��;(��R!Z�4��f�-�r��~(b��ݛ55(t�%^����2>�W���M�|�<�l�UԱs�˘2͉���[�����?W,jE�q5@QL�[��BB��iJEs[��#��Zsd�C#�$=�����G�:��j�ь����$���y=\)Jo�ޢ�6���fF�tJ�ׇF mj`{.����;#���?<�*@.t�"�8+"������.��� [ڀe�{Ҏ���~�� �zc&ol0��L�Ȣ=�~����w{Q��/���c]F�b�&�t���1�[d�H����7d�x�w��r����T���r��z�Q��U�ӥt
�0D����(�O]N�k+��Zr����5Y�-J�am�2\�x\����ܾ�˱3Ō�a�?iA��7�vwB����j����y��b��gg(o�Wo��Un	0�Y�B��8V� ����������^2M�a����
�i�;�N	�$�9YD�E����<��R�t\��9����l.�c65���?�pmd�HI�IKg6�K`��ݏ�[�o�ӧp�w�򵔢e��B�.�X7�����>�O�K���c�'�-
 ���r{ܔE.�~ ��c�	�-į�Q���"�;NTu<�Bj4@{4���q`���'5�b���aC+��O4rɠ���N�0�z@��N�'pY��j�ڻ{ϡ��B �7/?y��,^�yó�-TD��X��Dc�ˑ/=�n,�%8��Z��t�	y���[�y�*��(bȰ� ,���v��g#^Gf���Ҥ��ORj1�v9ko�<>�̉Fv�&�&�N:?FXe�^���:�b�����=d��G'�W�V#�!�5�Q��Pb�K�m�����f��.-[��Oc��FB��7������Ăw1'-�cJ����:���-kє���dHxsiF��̇����6��f�_���
����D�6vɚ�ܷ+e��+�j|;���y.�]�)q|..��d�TMl�g6j制ƃ!���9��I�~'�y�)���XLO���u�ݤ�BNE,��X�l�gw����*_�����%��[���-��]gB�o�t����_���7�ʧ�:�I]�،.�YdP��M�'�6o���pl� ��q}
]��TG�-�z��������j�G!���E��¯Q�nϚaBL�h�Q�.<�ɺ���b�j��Q7��g �����1m�n(����T�q��c?�?ի�J����[F���9�{�@f�2��c5N��.TI�!"�Y�;��-w���˥���Ms�e��*M��
���@;�a1�ۮ��� M�U���\{<�F@��_v ���#8����y�f��q~�L�z^l2bn8# " �4<^�?�kc#c��t�d���r׾^���'F�mpu�X\h��	8���8����-�*�f�?
Բ�Uʋ�/ZD�����{�aP�f�?�^ZVx�/�����6���6���)I�>�p���%DqR-fP��=�6�}�N����|�g߲1��F���5l�Gy|���M�9g��Ua�Ķa��e���w��c����Y�\�M��M�*&h&u0��=������I��|����S�Rגf ~�4�[�ĮbQm���J����׍t�C�#��	uol�,�Kܺ���k5�N^��������b]e�^�s���-��K���2�\�RJ8`q{������p��g���q���u�FSێp�@�a����-�nP�6+������KE�T�y��J��c�� �YKtY
���[���~�Bu���/��X=���md�mS4lzV7��0f0��Q'H���Iqh��'F�7��n:h���:t`p������A,=�����4���
�w�LL�1��-DQü���Լ��� ��E�tF�0�]i����u�wӳ�
�rݎ"@�yu��(�:�
x� ��is*����n�k��u����^Q���ͫ�d�b�����l ��p�*~�,X��Xm�j����O��ҁ���@��i'K�E��n��R\K���&�i&���u�2�ܙH�!?�귇�hM�Ԣ:��+Vu�.x�ֿ������a:4Nw��C��)�MXn�7���e�����		�<��~s���VG��k&�'8��"%z0�bj�>��~J�[�xې�C\��b��B�X�_���S�����_�"A�\�G�C�^rA1����,�va��I��sE�%�7�	�q��=$u�8�S�d���cC���%B��^�'{_�������B뽃9�YQ�-[��5j[0��qBGϵ��g����i�p~�6sj@.TrO�Ym(r��vAs�S	e�ú6v�r�e��{%Ļ���cskz��������p^+�M� bŹ���A�]���c��(�^� &n#����:X����7u���<��`h�	H��L�]����6���B�뢺Bɞ�p�>�48�}��1�1�'��ʓ"r��ܘ�q�n�|���P�ԺD}h���h�'�|+鄳��}u�-���ji�`��7��F�2넪6[O��'dtUA��kES��*�Ұ�#��%�������7+��>���+�ݗ��V��bϿ�wk���?n9�{l�>�Z	��O�&r�H@ɽxv�N����%���_��������0}�8�)�i��uR���E<�F]=����{/��;o0B���P��Gx��4�*�D�0��\�tb�jC�ڀ���(GQ��I�)�]�P����>X�a� ��؜)k�#D������'�a�~t2Ց�`�Q6�\�0��0��>��?	;����r�}'�������`���c��
z�!���t��"~_��Dė����U�ދQ�S�*ϧ,cn͙ɂ;a�ݘH�a&�j�mvL���5�E`*/~�}�^�3�b4����X�ԡ~�ʎ��sꪨǱ2�T΃#U�����OP��E��jxW�ɺ�A��;�jj��VUy��ʁ��1SsOg�^�-��[iBB�/�c�ʃ�f=�uS�������^-2�@��෌��`�6��5��"�����_�A��]��T����f�5�����m9Q!�"n3Է,��\]���[�����Ջ/�h>II��^s?��j4��=�	o�z��fyU���b�j�dn�w��]���d"�J�o+��/`ʗ%ps��9S��1K�S3���W���X[M#o�#����P�W����UYҲ܋L;R��-
f
�Z�N�y��2��X�i�[����O�Z��8�mC�yX���!��������'�ܕ��mg����zc2�����Y���j:��Z�\f�F�*bNs��8l��<c�ֲ�АT�e�<xr!��%5t�����u�ܫ��j?/hcÅi��B�P�����p	g�c�|�p��[���%~6��i����(K�1���z�J[;�wn�6�$/��$:P�)�@���'}����V0W� ��%�D�լ.���#���s��݅A�X}P��}V˝[����w��*[��?���?r�b��1)N�]�=���}T�9�i�պ?����I�e9R9�$�� K�ŒFq��,�M�`!h�}ƺ�**�5�_|ӡ��b��ngqۿ��Q��.��H�3���|��3��.B�*�����6T���!�n���#���b\\�LE3D�@�|��
��h��j}�Ce�ޓ4?��>������R�4����a�9� R�TcA�N�ƃph�]�_G�|������ oMS��_�������hҩw�Ϋ�
o*�䎚Ė�,��O:w��n����Kx�!�œ庴z�v�Z?U�o�d��z�$R�"�ϣ
�=����x9
��b�#��݂��_�3��̗E�E���\�?tY*Dbư��2Ud�چ�J�8�Rc[����5���*�}�QW�B���>ݲ���r9^e?iV�S���#���w���8�Ą���,f��r3?�`���嵥�����1�$�6p�[���Z>/"͑�Gn��#���L�:"�gR�ՠ�"8�W�Z-=nA���c��;�3���x|����+�����8=CE�E��%�"�I�wIM�m9 �;=y���e����J�>�Ԇ0��-�I���uj�]��#dC�N�.ԅ <X�;��L�J����FSz�6�j���Es�	~���g�vg6tS#ɥ:�����bX�X����
-�cVq��)�s��V&66��5�>D/_j�I��AA,��r���nR������MG_�l�@��dέ�'?�-
T� _s+ǲ��G�`^-���FÊ^����IޗW���fL���-��+c��D]�={?֜M��7Qt�yR~�B&��!�g����Ġ���d�)4q�*S"D����@�0:t����(//�ߔTA��y��+�XYW�ͨj<��&��y��e�]�A1'(4�z����:�Hi�f����4;P�e�,���P|5b��R���/ �2�S�9f�Q+�U^x�M������|6�W&���U��"��Y�/P�rTM�T�7�:�Q�t!qt��)ie���i�E�����2�	
2�&��Ϩ!��e�D��=.�D�~m_�G¨�AO�
�"z��/皌�=�2��!/8`ur\�YE�8g�Q���^�e~�j���[?�s�g��]A��p���^��yԼA]y͂��i
��~��3S�Z��`u��{\�n�,r5^�PW��jGz���� �ߦ��쫐��~>�&��*�㵛���}�c�ؾ�I�dp����dnM�,zv�@Pn����=��!�%=��C^�c�!��o��D�e<u;'�P��iΡ�2)�'�n��c�I������ν
�X�����ʍ�_n���ؼ�������̂Pg0Mu0�O�>�X�}���i3	ʽ���7�Q�UP�g-��7�����'����oճ�p�y��i��rV�k��K�}쟢V�3�1[�z (�;�k=��+�|P���!����@^��Q+��x8~�p�Ǳ��QBX��.�!�2��a����fEcs�ÄŦ��jI����~�9<��	�0��3�941���Y,�EO}��OS[�R��b8ߤ����BZj�QF{�x���(�~H�+�1�����w1�}m4��c.C��R��O��V�'am� ��;�_�[��{ZJXی�����W�+�	9ޗ{�ey�4d^�B$��Y���ٕ��~�Xx��.v���K��g�L_���'4Ή�ٝ��=ҭWF�P�bˇƐ��d�ѱ�o�5v��.��������b��V6�����ϥ����2���F�tԣ��כ���ӽ�����L�a�r�y��
}#!}a�!��ɾ`��ܟM�Y&��W=�"����`�ݶ8���z1䥿�N���bn��*#y<�"���ݭ��|��u�qs��.d;��$��i��k��f(BՑ�k���f����xt=�/�O��{� ��!Lv��3&Yo��i���N�M�e��.�\�G���~8��P{�v�E����֋��a��m�g*�9�]�Â���Y���a5^��:��slXL(CIK����ލ5֌J4�ao53n2[��bv�����aƪ)��
�B����iߙ�6_lR��Nd���s�;��Z��Fu�	d��Z�<ɑ�/��:�Ob
3j��p�RD�0"�Iyw؈�_�Y�"ॳU����/��2ԋ}���S5\8yo���\� ��+|>va�d���,�����+n���g��D����&�_���z�x���DJ�EoMf��\�� w���ݜM3l3Ax|s�����6����N�q��ܘ����c�18k�sw۫K�a2�t����JX��%���m/�k�T۞=`ڙE�:�h��ߒ�hw��Κ+g�6^�1M�1r��y���Sj5͞�;D�*�>�~�$o�Ȍh��
��Wy���n�R�.���ݱǋM�P.��m%�sB��6��(2裬hU�GRA��y���2d�p�l�W����y��w��8"��C��S�lu��ۨM�wˊ��l�1�Т�+ޅ���@_�x��ם�o��>��г�r��>�"�?�p�#���(Mn3e����?�s�36�f���=�#Y�PUg8�4ͲJV��ܭx��'�[o%Nd���XB�T�0�.4Ճ>[���R�c�������-zчl�G+s���ɱ��_{�Ʋv�2��}<��[��Z3��%��G����!���&�i�*D(�wI&"�[n�emF���O��)�r��L�LᏂ���Y����H���X#K��!���n��ϒG]���RE�.����/;��CP\��?;wMB����z�u�vZ
R�4�UZ%f�_��!�
6.ɳVxX�.��OQ|�
~y*/7���i���(^l����E�_��?��ѫ�����3nns�шe��	�|�����C@vj�pH�AV���pL�Ѽ�"hd�S��!�$9�-��tx�A��N��j�$�w8��Ȗ�0R� �u�������9t��r����1o?}Š��k�b?���>���s)RI!gZ�{�{0Q���@W���@i໨���=@W�����:�P��*2�u��;}�lZ*ZV8�|�?N):�$V�c����(u����r�:�|�v�W���z6�"9�D+���jx}���0M�o��G�����+��=�A`�$���ibqn�hpȪ��_�*aY^i��[�� ��j�E���G���
�ю<	}��Ռ�=b�=�(�u����k�Oy�Bb��2��Q��S2Z)_6��H��F�VWk����=���nΓ��{7���.�m�q�m�c��	��/8�ډHHNs�(':��6��n�B}�k}��;S����C�lY����Nx���H^��գl����A�	,��x�Y1V��6M��[X~�j)s�e�\?U�a�F�g�i�S�r�șQe����Y���d����/�Χ�OX��!|�����:�HV`����/OXʅ��B�bOt��^�A �CXc������!�MVi�K}�A6�x��7E<�g��bF�P�!�ړWa���L�rr��.��8�$b��rQ�#t5_�j��t�I*�G�a�y%S�9�:��(���̥�/k�Q~�ϓ�0`<�o>dB��w���HƷ;�ad_�������-�5�ʕ��E����f ��u|D,ਯ,�ět7�)u�5��$���������g����	�yn�]d�]�rm��{J'%��Q�y�DtR}E?q-�t+OI�pplY��vcQx
y%�k�YKt*���,�>�wQU���>�Ԡ�2�,b��Rڨ���6aGx�r<���i�0�M
/�q�tQ{����ڛ���]���֏k��iU��4�O�+�1�=fqo@���fEǥ2��&I��*@Ä� ^{�a(N�G�.`�䊥��t�|l�/[��}�ݏ������q|����3�������CQ�P�1	�,�Ì�]�W��`���ZQ`حz��X���xWG�O�S�'�\NWvD�����  Pm��Bw�L�s5}�I4��G��!��b~�?�0(�	�Y79�����ݳѦ*^R5L��!ƶv�v�46��5�z�;ݞ��}���O��t`]#�1�@���A�KR�q~�=[RY���Q��E���}��I�շ�^"�!|G#'sk�����w���cj�'8����W��^b��0*ߕ�/���J<�O˳2㚅�U:��2f'��nƩ�w�n��:�K�AC�C��F��=@�2��$�l�غ��5(T�3&_:��Yﯧh'��⥚�~��4�T��6;����.��<��t�d��kX
q.�&C[]�1BD�˕�%0W�Yz�7�z�u�� �j ������+�7xЖY���Aa�W=�0̃�c<|�W!b0~|���~p�t$��r��"�x;JC��	�5�ͫ�v�I�����N�F����&3�O�]N�^M���#��D��@(�V���t���<l�w@��2�6kHz�a�8����ia�r�o�.������! H�{L���Mf)?�����plU6�!��_���*��V��㻼���\e�h����K��o�&��^�%�G��>�ʭ4Y�R-SUt��?�8��\b�Ts"��O�x��K�y!�W�ڽry��z��D#��C�&<��1iKtJ0�<'A�F_�ް���F�d�q˺���< ���P�>/�Bwy4i�`���G�5┯؊������	������������ß�wn�x��bȰ+�D(�LW�`0��Kz��!\/��n�¡��j��)���\ܣ�p�
�ؚ\3l�2py(��v�����Ǐk/Dy�|��N�C���W��fSF���n�s�|�6���Y���Z���q@b�cI�B�U4.��<���H�o��{v���P��ll�׾d"��70�EX�����g��Ǯj�R��<��R�kv��ܡ�_ܻC^��6�c����Hn�b#���֊ÁN�{���e���!G����W�UY|�y2�`=x<	�_���iT�6�L�*3"�z�a�i���P�$����)�@(W�.%��ϛ�N��>~�}b6�E9�����$΍zh43m��UWǫ[�l"���%��s$㪝��+���JVg��9�^�����u[�<�$���@��(dv,����5LC9�p�����<Eo}�L��b~	N�C�&�
4�@�`�Ҟ�?`��mn\�Q��ӓSk
{���;��{nlZ�r��������,t�2�W¸[��m�·?�)��kE��PZ7n���/5��/������a����W�����zeo���b�������td�%I!;K�+��b�m��\��y������Tߔ���y��������&��6�ƶ}om8񱱐g�w�O���O�#�I����`H.�[�W}f���7%��(O���l��h.��V�>�`#�_��g���	T��md�הA���;��3����p�z���u��.5A�kU{���N~,��9�^�"k��B�z�FW�9:,��c+cJ���yX�kt�T�=��?�p(-�.l/�L��KA�v+^>u�xg��E����VLp�u��͏)�����^��K-�fj�1΄ ����[�d*ҝ+��f.��%���C7�Ʀ2m��֘�w}�7jû����\#Fľ�[B ^1�;��#�o���N�3SNGɪ��;N�D�3�����:���t�oٍ�zS����+��ܳ��M��b��%8%��2�|�C�v��V��w�6#\<���V����^���T��e�:9��,�)3�4tIL�W�q?�G�e����
,{����ߦ��||�Kr\��xDT���LS`��ͳ=�9D��5T��p�����pp��f�?��0`_B���~��Y�tC^�����q��U
r�.^!��xQi��i����Q�"�j���Kf�ƅ���R��3��������ռl}C>��~N�,��I�������9�i��fJr�t�J���������)۩S���Í��n�Zk�6m��ǘ�-$ ���]P*!Ha&��w� �����3�����i��ل�0*���%�.��#���^ "hd���uzX̫�JG(��2�/G�.��{~B�+���}X{�gI�u���Q�Xv���?�5�{L��tlRD����w���oy��kvM_�d��TX���c�6��kpM�;��`�\(��_��l�.��^�L�y���Ly�U�S���Q�Ec�#����{z6�j�Smr"�Q4��n�g��麖^&�*����x���m�|vs�;hݕv����n�F�Z?�t4�u�N�ȩʗ�����a4���+!�N��)�m�/~QzUx�)e�#��+b��O�	z�ڥI��<�yj�*'�ec�.E���mm&�/U��iF�:����
�vR�W"^�jl,��/_Av]b�ٔ�]���"_Z̕��c��y~S��؊��|����_@BR�QW9e�V.�cb�62�ѵ}i��[��)�S��Q��S;��0���$��31���������r��#ו���:��X,�� ��t髞3G+���*�E&�A��]��:���*�v�G�k5���\��u���[E~b��ZC�GF/[�µ2���vF:�ɕ@l���r��̟��u�2���ͱ ���_.>j9��R�)觊IO]5u�@G��]Z���S���DX7r)�������lس�������6ѵk���9

e==c��ےm^G�|��a~�u�ޱ�!�Y*,��vⓅKٽ�[�4�/t�R�+&�	3�Şb��?�^��9�)q�K;�u�y�k�y�$�9_��8<`����8D+��);����*;��$Ѝ?tx?c���[J�W��Ugn����ފ_6}�s�&+�jre���Q��b�dW\�iQ	e���]~Tec{�[1e��oWv�:���3y�(pɐخ�f'+���������·�B�־��i�Zۼ���tH�-�$o���[�^��Фt����E��u�q?,]����Ӆ�/�8[AB	<�DVg�˷q#�f��G�xGn������o?LsZ��ġ��7��A�tS��p鶫�y�)���>��S4�_�;5��TL*z�Dz�ą��u~d,;Wsu�y����!�vkN��Rm+gϐp��7��v�V$�Re��ب>�'��	ce�`U��'��11.�!�I^��ߕ����"	xmR���9s�7;D�E���l�t��.�ћ��[�;����W^�cNg���Ặ$��a��a�k��|�Y:�'��'�z�_ �:8�Ibf��t�T�1 �8�ې5�N�\��D nF�ly�-����{�OĞB@DA/�q�$�Q|����l�v��������./�^U���Ooo�4�a��C=�`�;Կ��_3}h��u�G����h����\��ߞ��0�mzO�������ш��h(�T�̠��_��	L�udC���LW�4 :Zh6}vJz��R�f�ą��!��� .�����<��Y���C��0;:�����2��Q��*�i��_,��W�
V]/����eU�n(�p�q�@��H2f
1^����mf­ۙiut	�v��H�	��#�@�.�E�e�t��l�~���1�b�eK6؞��zjf
�U�""�������,{$���<v0��9�Ew^K�_5����X�P-a������;�K%Vs���9�$��A�>�<|�ɫ�߸ޠJr�eh��Q�k�8-Ma,���e�򄇀��%����5���%��u���I��XW+�8��O|�!����!��ߞ	K>���g��� ��ϯۯ�KW˶�[�����R|�vј-&6�0����-��"�5Xe��k� �'C
bD7ͅ�M���1ne���>��J�}�r��vp��f?	��H�D�`r@����b��;��O�5�9��f�U��4�tv�OI1y��i���ׂ_@@|�X�g�'�����y��-q��AjY�CL,����9�x�.2ӛT����!#��F{sō 5�	+ϻПe���.�:G�8X>H�\5�oQ�]��dPv ��>ة)���1[{����_�������_Gk��.n�k.��7����~ms�ǀ���x��k�:�@��u?�XtT_o�,I�U�KO{��%:��U��R
c2�>ltѷG� �%��� ~b����el�&޼��bCXN��;&^d�'� ߎԺ	$�bq�G�f0�	h$o�2 ��Ǧ�wU|P��O�F #&]�;�兏 7fE�j|ύ�ܫ�	���q���s�Z� i�%h1����ف��~݉����?ԳMȸD[j�'S{Cl�i��s���l�+���/�k�#� �[���Fe:�����#<��qA,}}$.�B8!d���P����c��@��j�� t̮�;��n�76QB�ѿSG�Ҕ��o��J�a#�y+����������#E�C�j4$R��(-���-���Xԥ9@>^X����u���LV ����߃��mB�N��VjBڿ�W:1��Y���,_�\M��44�5���F��/� CK��%��8�y��碥���̈t[�*�_�Y�Y�v�|y�i�9���&m�������Y��G�+��~�)+ܗB7�����.}�^���ޙ~�۹�܁ט5��O�F�j��^T�|#��/9`Yd��-F�e�h[�i�8W��,Ǭ�w+�	�$�;�{9�պ��}�vm9�"�T%�`}�)��b<nx]��C���������s��R�(V�s������Êءl1�LĐ}�\[�н�}V(�2I�KJd�3�S�J⑒�W��i��*�����Ѻ����RY׎4|�@;E��:�(�umdm��[�� �jӿ�sM��?����n�>ڃ%����'s6a�8O'�� јq��.VFn��&�2f�3�aӻ����H��>��������UW��i�B$T�[�1�u��c6s3�(1#g�Z�|i��ĵ��
Pڽ;sKhk�0������7Rp�p0V�=�� B%��n�D]�`��l ���M�;V��?�uaid������RH1;�<��#�o���򦇾<euj�g�o��pi9����_�0L���RX)�����c��	U���9]:�9��R8	���4��\x�8�N�A�0K8�_Β�~k��5y5?���UŔ����v��cK˭V˔L��Yi�qv)Y����s%�����R�#��M"� t$?�N8ٹP՚���q�SM�t�!H�{��(A��5Gx��'�<�*�u&����9�,F�~ѓ� ����kA�5?�_���n�Z��2BV]�e+��Ǧpѱ>=.m�Xh����,9ut���2�@�[2I����ielU�j���Kf	��ZJ~n������B^ZP��/�.)��=����F�L����J����?�O�g�wjƖ��'�y� anYL���k9�5;�>��o�%JM�<��[O?4����S��������N�ջ
;"�*���eӯ��?�#R�,/4E~+,�Þ"N�m<m3I@?��n��p�n]\��i2Bc�@0���`x�(�:����C4#g@u�ә��Eu�W���j�����H���
�%>�΀�Ǩ����ӥ�E��Ӧ.��l�]�	�.G���mC�	% ����l�<uyj4�%?z��x�tjӠx,}�q�7m��&$#�}|n������[Zec�l�6�d��^�쪮@��B�2fq��M��lm1������ƥI��0��jز�KA�p�3��8m&J������}�WO!jP�$G%��hG���'�c��ѥˍ�3�8�����t���E�Y5\";�������C�ƚ��Z�!�Ú?<�㧓�f�U\���.	^��Y�B�������a����v��E�W��
&J�xv3� ���Jk�� #oh����a1W���_�A�˩3�	����n8��R�����e�x�69���B�J�l��n�^3��i���3'��� �ߜ���/�ڨh.�LOPYHQD�n��=xJ<[�)n*��(A3��h�}���͑��~p��ߢ@��y�x@/��Y\B�+8o����4��墴|��AE��U��Cs�9%��o��]LI�fo��$�4W��:M�G�~b���a��GQ����
�ʥ��}~�$�ڔ��.��V���/�v��)��j��ڴ�֭�$zI��21�ޥ��)�:�[�g�Z��՗��?m��ITZJS�$�՘��:BKL��J�x�i��of�Fժ$[>��O^Ĝ�*����P�O�.@q�`���lt�.UD�->R��2�3�����K����L��Zr�`	�C�3R��׻�`��+�ҽ�n��y�--�]��o��ڒb����ԣK��u]��D��\�B�Ȉ�?�?����]�F~��鄦k^~�/����G�F�5Ɍ��	�Y� Q]���r�~����i������j���(
*%"-�R��*RR�#��{���! -���1B@�;FlFo��������sv�n{���y>���Jj�q�MF7�@#��~��ssߪiQ-M:1�},w���t�J�r�.I���{������4����6�Z\���P:�a`�L�X�2?D|�C��z��l�;Ș[N��\��{kj���L��h��^��lZ�:�%�<�d�Y��i�A��L��d�������b���:sO.����D|���3����tba��8�����27�e�P	��M�oٔ����u)���D^��8s����r����ӳYL�ڙT\[Xe��[W�����X�F���.'��2�R;=�f�3TĐ>�o'Z9�6����ly��\\�̀�W~���:>���"� @ד�	'���N��V'���u>��@�BCpm���Wǌ¦Ûu��~g_3���K*�oKe�:@�ӄx��p�v?f.A��j�������w,����Y><�t��K���ɛ)�3 ���"K����<m�N72Lm�dP��}T�oy;hq�`ݘ����ٯ���YE��j����D?��xHU�0�����qi�7�۞�� �`�;`j�Xc��vc��fsur�'�D I \g5۲T ��MBt�7ǩW-3a��5��P��Ʒ�W�/�IG���*X�uo��O��=��X����n�D��M����������ҩmq<tX��V��)�\�U�%�K\�ϕo�eZz��e����F��zt�j�v�u^a�Z�mU@�`�g����.��W���.YY[��bӁ�@�ٓ��]SAD'�v�)$ѱ����󂳘�de����t��\��#�����Y-�mTʳ�'q#�}¬�g��w^r�	Рuvq.�]�"ꪎ�P�OI��'S�e��!NA�2a�B�AzGΌ������O#�K
k;a��r[k��?!"��A:
�r�ǯ���O�s-���O�M'5����Mk�����
�D�?U��V���6�i�M�ysmZ�w�0i�D����~��
.!��p�Ni�m�f��PP�Y\�����X_𕏞׻	��0J���!�"�`m2k亖Z�e=��?�l̖?�2�kh�����ag7��S:VD����s�ֽ��S�qF�~��Z���f���w�4���Z���觛��\UU�\�`!:����OK���U��ǃg�bW�����/��DO��,��Q�����.ʅ2��g1�R})ǫ�|�m1&V�񾱫�ŀ�K��E����'e;W����8h@}���d"��	��݂�����I����V������C��*�E:I�YS��q�� ��H�.-�NI#��n�OC�PV[}㮀��C���^�`mTL�k條�}z��x��q�k�Unz�<�<?��*T�;���/1:�h����@mLĶ9���`ۄ�|����� 	�	u�Ӥjn.1��j�p���L3q\@F;�����yu%x�}S#��V6��RC	�>|=\췇N�[���Ӆ����V6��b�@K�L��z
�i?��o>Wk&�Dǒ{-g�,�:$��Yz>��C0L%{��AgUv)n^9tNT�[{�0`�������V��R��EZ�2h�2�0lq&�i�hrQ5n �7l5�T�8_� -m��:n���X
�-��u`�>؋�G>��e��"Wɥ�N�<s�Э�������vH�s뮩u%�1�������xue�.�f>'"��n�"�S���D��4V����E1pE�����/Kʌ��(�u(.�𖛞{j�3�a+�q��3<zc��Kt��#I
���_ A�%s���6$�.�A;�`���qX&�el:�<^q`hͩ���ƴTQ� {$�A���(EWV�͈���#���W��������Ҽ���T�~�9�ڸ�R�tc��@�O��"g3f�\&��_�ذ��E{����"�����7�c�$F�p����0z	��tf{;*3�������ߦc���� ߾d�:��2�p�,B?��GZ�����._�?e��1�L��Pgj��Z�8z��"P��ݠ��m@̈���%Ԡ��ĻX����Q!���"U~�2h䦠�E$��'�T8b�ۅ+`4נ���c�0���Q4M�USV�����ݢ���Fx�
R�]RR%�>�M���lZ(ZT(�K�)�`������NI��ivyǶ<���&j��]�cg+kj��7ފ-Cu����Az�>�p1	�7�d-u^�\�{ƛ��:���(�\Vi�;?�x5̖TN���>����T1���w�����@�/=��J٫b��8h������>��a�u��G �@k�L�I�,�^Ɩ[���pXm����C��V.M�]��+e�a��g6��g����5�&�&��s�&�o��7�7@�=,$����W��������󪽌Om˺%2�:�[o=T9�T�	����07n) V�������_c5ȩ+J-�\Uu�u�O;�|�H��n���e�}P���v��/s\�Egd�gRV��{PX�#���Uv�e굢��6� l�g�u��'ZG���H0�� b5��1}8�j�5�:Rw��o�:{AϤ�Y����{�4j�ˠ���s6M�a=s�O����P�g�2B��2�/�����d�'��V
ěj��hN��1`���Aodb���X�/��=~�Z�gr�l<?J����e��;C�`���`5���2j�>
(l_�-������`����ݻ���$P�;�C����	Cj���\&S�Lr-�rF�!-"G��M�1����+�62C���T�QHE���S�;��v����-� 雎�ѽ��̨0	+Km'��6R�80(���Fl�F��/��H-1�2��C�Z����.�Wi�.g��΃��=
�)ʵ~8��.�w_ӵ��K�+shq�y����Jx��йղ/�3�Ü��A����ef��:M(ۦ�.u���8��xz�OâDi�~�A�{J��9?���%��^��6f/��U �����e�����3����/}�1mk�U�� ��+[;�/<�TQ�)��o���-�(�Ύ=%���7��d��(�zeēw%?���a�	���r�6O�I.�=t[����y�3+X뿟���Ns����Z-�2]o��64I���w�A�QL��"�3���$'�xo7���0$���q�����%o�rc.�7n�~g�wj������|�\���]Hӛ��L���5%�:��~�Ġ���cߧ�ﱯ��2G\��#�UC�q��Q̈�'{(l��rج�z�ꅴ�qA�d�xw�W�T��/���:	:��>�GC�ܼ����`���a�m���e��f��\�]f"�^���pVU�cs�Pb�����!M2�(��h�J'pU��m5/��]H#pY��Ɩ��R8�wq��⛍H�B\�v��l����(�)�Um�B��0��ٽ_D	��fPף��5Ou("3K^(�4L<F��&Lm�� )q+�}�#v��S��5^�+�c?s2@�C��)4\R&�!8Y6��K��-�&$M�%.L�����O�kG<w��7��ݽ�����D��p�h�)eY���T��J����<��犦�pt3v��B?ϝ�^�/���ֶ1��-)wDҬ�Յ���;�t�Z�}T$���T}2��Vyő��	x�EW�O�wŁ1�������f�}g�X���;�uf����
�?�o�ڮ���G�!;p� ӽ�Bha�I�8酁cm���'��sI���j�T��Xo�"a}~�^�=pz��z��_�5QoQ�C����7��tiQmQ�X�A���deq"�G��9����:�J�K����c�/ ��7����]h�U�2�/&Z߬�Y�_��Z�Sk������D[­��:�h%��X�r�.����x3�G�[]�	
�-&��!;�3�tu��z�c��Q�@������~� [��<�d_%�t�,
q󨃪��������
�.��֣W^>(�$Z�}��x[�VWS�[�[���6�Bn]��?�Fa�@�������1�V��]�z�(�+F���P/��������t���
cy%r��3ӈ�i�ġ�>!%�4��H���w��ѻ!%�X�ZƠR��˛�g.[�(GEz��7/&���wb.uHS�����Q��}���T�7-�2�C|�|1' ~.W��3�A�b�rVF~�y�A�o��T:��@6(��׈�M��f��}`���x��S��j�kz�fGb��Pڒ��~�EE�M�.��Z��I�[�[#�8B\m6�bh��͸�����j���;~{�j� �Y�m�u���H:~ ����|���%�I�u�aU�L��^�Ke�_�5zTy;%Bl����b�{�t�mC�2�5c���g4g�C���tS��U����Q��s~��g�}��b
��LG��_"�oP6�S�`��v&&no�$�XS�F�:^�@��Ic|1�9��֫NIۂL�d��Ok3	�[��3Д��� c��@7�����dT�{m�������i��~�H�,��e���� ��3 ��Q9�2*}6�!vD�Sf�F��yP���3}dՙ��d*z}Ն�Y���bEk_�o^*DLR��v�K�9��-�;���L�䠂�Z�z�9�+��ɮ�J�'��k�W�]��B}(�`Ɨ���b5�s�$)(�r�Y��$a!�Ҭ=��� �˞O8�dH��
�%%���DL����{�=ZOe��������,��`+D[�n�o�@�*�^G�ϗ��1A�3M?�n4��x��,I�DO�.GAx�ܻ�����#���(��Q�hj^�����sKw	�]�>�v1=�b1 T�0�i��n�25H�5�i�v�?j��|�cI�Z�#JZOk1��=��9����߽!�1!#�2��q��
HY�5���2+���>͓����-��G�b����^y#e�=��)�e�ހ�;�SL�u�B>!���Ċ��W��&�k�"�0��Y��AM��^_��,�#b�'�=�~���,f���T���TՉz�q���js��[b��~�Y����A���0�/��+�i�q����BT���a�����ֱ�c�L�
��_lᬨU��W�Oe*�M�`h�5��Y�^���4� ϸ�n�Z�>kKf{r�ʉ�$�>*�+a�K@8��ƫ8rАPˢ}��������7����"
��QÐ�+Kڅ6�^����tm�ǔ���`)�q�������"���O�ю��9��H��i�pu�kЂ*��}�M����BJy�Z����c*�%�YYa���n��_kl�1E�W�@�Y�6�#I:_c���KQ[�����/@�r�������9L��|�Y�Do�٪�I~�
O������w���y���؟�14��b�d4���bī��T�&]Z9��ٛ��[,ϑYe������� �Eۿ�y�i����1�M�mUJ|ح�V/c8�2��;g�!���fq�"���Ba>�1����N�{�o?|C+�c��M��/��:����#�>7����awP���x(�rҺ�.fy�~b�J:���q��ߢX�₃��(���7�/� 7z�9G�Ǘ펋��QN���Ym�:L��͂|�'+�6����S��tA�4U]#?�q��l�K v] +,Њ��~2�s[�ޅ3�T��R��-���b�|�Q���I���ӳ/�y�II���%�J��R�=�Y����L�ɏ(1�ɓ�#=XI�Kp��K�~��3��v!��85��H�g��7��v��"p:�1ʓ�T̰W���1�y�<���(�
[�=v� ���i��`4}�&�'+I'"cm�/hÒ9�e�F��~����͔o�wB|��mם�X�N��nN��.��t�^��K���ŉ���i��b���
˝88q�+��&Zwd�<�ǧ��/�/&t7m
lG�T���B��q�v_�4η��b�g�s43�ˇpO[�@ַO��;�Z��׈�l���.���3-k�nJ)D����^X`Vn
@���qS�b��evc:�)� ��c���++S�N��N%���+�+���4Aa��d*Ձ�b��suԳIw�A������(+Wa���
�Ig�����>�7��7��%рs�ӕR�E��R����ڎ�&���qH��x#�l6ݝ�7�Յ,�����_��c����g��>�`Y�i �b��O��ޞ�E��`�a����t�g*�j#�8�k�p0}1�w#z;ϰK���Ƹf�&�=���MB�S@=�&�{����
>�ᬷu�U��ֆ�P�n��A&�d�9�](8k�q�6*�GJ���Ci���yx�	�i|[zG�kV���nο*�`ꡙ4@���V<9F�	+�P��h��A��^/X�h�%b3�����9D�B��T(@�V�_�H.P'��ck ��ó�8���J��@k��V�@���e���T_��: ��vn�`��G�`�7F�_�k�O��~��n�0�n�h5Kʺ�v{�����p�����^$xج��������5�f/]+��D�.�{�h:�GS��͠��?�G�K���f�N�#�[>W�� s�FJ!�e�}�6bbF@C����WE�O��d:����J�����z�hF(��J��ǀ7�q�,�&���Xޱ�t/�FI���sFb�u��s቙Թ@cb���~���۩�����LO�5�]����\��16f��~uc�{ϫ��/�r����as�6��JQ�m���3�i0e�N�׳Q�������h��4�FW8��2n�ɍ=�;X���� ����+�/��+��	֢���\���L}�bח���/2��6]Z��=�c,�k�f(&���Y��b����Ї�ǡ�ym����e�M�"=�x;�:G4=r�T
 ��]������ܮ�n�`��F-�#�`�j@o��؟���Ͷ��B������(�tX��CZ�k�FaFR�頾'Zj`��U:��������n۳u�L�B?;$�`���I�#b�v�t�
��/���8��I�
:��7kտo~f��gp���5����g��U*��t�cta�W�"dΓ�:��qC���L����7'n�����f��3��G3��+|�6qo�"M�N�Q.�KxmBa�h�<�xqsZ�ow��e��:��/&~�q�GѴ�Y��dtje&>�g{�A���M_m/�_�{��B$1mkL3vӱ���6�g�b6-Y������:�6�!ţ}c,G[5V�/!-��`�7�}<«�G�g�^o��'?Q8<ݬO%K���l�%�����a:�u����<�ClB�p�Z�+�K�O��Z�1w4K���PCӃ�.a��j�×���ǭa�k�V�q[�o��8i﷔9����8�jU�����,�^#�CL��:�Y�f����:�4T���������!�Bw���[�l��.���M�_eZmm�,Y}p��,�1e��xv�V����YgT�".f���+kGK��+�8�S�X~zf06��w�2��B��j����^l\�Q.���)(X$)���}�֡��B���K�c
Q��|��~��}5�d���Z����Z�-Fk?�<[y+��<1����a~��Ǹ�lTZƓ\'!�w[g��>�*a�`L�����=h����?��R
/§�v
��SՐ YKh�A�0�U���ß�m�b�2�����;�S�����g<�7�[�eE�
��g���D1~H�e���� ��ၫ��xӹ�~�.眝cB�N�(��_����E��P$[ |��:�b��N�r9C�Wp�	�����/�����fq�ɬ�tä�_(�bά߼�+ƯI��}wm1��l�9�J%M������{Z7��8>��9*g$�sz:}��A֔W�8�Տ3؍^Y.�z���$�׍b\	Q�����d�!(�NmGUq�����������e���bW�9�2u���P��[�K�|��6X�>E_6�-�uA[S�|�-P.kP#ζv/ҏ8�?z�d\��+]%Ex�%����~���M)�O�x.��Q���XS�;8��ټ�$�.$��0U�]i���m�C,Хe���~��G�괈�WKD�6P�O����F�G�ˑ�Ķ�둁<\������EBm����+ўeTޡ���w�^�����n��G�=�!ۆ�@��Zo�O�x��, /�<R zW��}A�QkN_���.I�ͻ��"I��=y�AR��}��}�R�C���>���z�����g�� ���l?ę%x����
��z9�_�uWW^;-M�@��Ŋ	�>�6�� �T��Q-�@[t+�b����zEy��۞��%˾h#�@��$,-,��2�|Ii� <Y��Ks�����5�	�kx��V<��_աL��_��SyrW�ͼb�"����i|_�]8Y��Qh�L��?5�2/jȚ���M������:�0
s�sh�e�Bݠx:DQs���'s@B��HV
 ��M&�a�24��a�ˏ �$� �d��ԍA��2�̆��B��9�>6�랶��r�ܪcS)����-G.��}4=� �u��l���$a����X9T�?�8���Ѕ��w�.E|���z�<Mbb=��M��P�x�S?m�������'���;��"���5h���	y�_Of�
�L��\�>�����*�?"~�zbc9�d�5��,��r�Nb�hJ�]�&����S����8?g�9�ð��ْ��PT���N ��64��7�,�Hra�<Xg�թ5�`$�nq	�ø�u��X {���h����71�L���l�vm�r�#!���7��P�!���I�E��5q_FƂ��O���ޫ�n:L�꫎'��2�I�5�3�����׫V�Y�hN�ˢq���5�F�(���|�7k��+ R^��:�X���&ېkw<t���9i�浛��RB<:��}�/Z뷾����r��ё������o���5=1PL�7�^�s �k��W�Xd]�t���B�f�Թa�2Ш&3Eً��gX�\aX�z�9�fqS���hN��Aol��ɉA���n(�w� C]o[o��P���:w�?���G��:
������
L-0`6�1�)lo8g�M�z���3��D`���~��I��n��cR#W��m`��qUp�x�H0�B9��qӷ��x{�f�T�n�� Ǎ,�={�oR��P�-�u��г9�=gQ��B�EΞYy���V[R(Zj��:iK��7z�ij�a ���>�'`��G���sN���mĨ2$��en�ڴ^��w*�M�K���>B�{Q3	�O�+���#�ۢ���m1U�'
99W��8��ڇ�}�A�h�9n���$�)4�+���c����|��65����kRuj7�f�w�-@��B�Zy� b1� ��]�tN��Q0�-�_X�ȶ�r�󿘘�������U)�\��>��*�3�L�]�y޷���f�\��UiW2?壋_�sOg���T.u(�k�Z�u���S?��ь���Y��Z�,+	�g�0�Y6��=Mg�M,\zx��cn����6���¼�x��I�f���eK���zb��k[�ˬ3는�,l��c����5|b�)�S%Br�}�.E��� ��'����'����H�;'~y�Ӵ% ��Y�܏ѭXL��wjB�2g��6������1��^�9 c����p9�E���H��e��K�q��
��[�k� m�.o�_%.��$���w���j�G]�/�'*�vS]ޘ����z����d��r�6��:^���B[զI�vuebo��a����2B��`@][C��Kw�z��w��G�M�1����������g�K�_������ik�go!�j���-��d7�{�m8�40�=�%mӛS��"�8���9��/b��*��Rtї��p�7������M6�7�q�Z'�=p��Ďv��p��L
n�7�Pߌ�I=61}E�@�mU��v8�u�S�BA��.�	d~��\���rrA]��I�sq���[J���[&�@�;���9���
"JZ�->�4��x�S���A,R���y�<Z!�x�Z���')���(7��0��K�*�)G�4�O
~,����aA�����&h쌽����;���]��s�K>"-];2O�
-KY����h/�%�Ԭ����a�t��J,������ ���3��C��lթ;���w�p��wҤ$t?�^"Ď3��r:�i�6̩�\���d�G�Ǔ��R��+9\��=��^�$���Gp����y�V�uZ���-Q������ra�IQe&I_hwZ��SЧ@�=b�mQ��� q���oO{����N/w�^��6��,+k;�����.t6]��G-T��1_���?�.���m������]���U�Ұ��s��?���<��&�e�S��N\j�akm�f���%�����X�}�˻�������:saO�@����*]��T����g����]���#�\A��˽-�������٩/9���Y9��[}T��j���jĉu>�=}6������~�Z|y�m�7���YM��E��t�{�l������ZS��;*��}Ó�w�Y�͘�z��}-�p6�bK�%���%�;<[{����q��S����\q���x)C2�̺��
��;Y��vk/�ͯl~��~Ͳ�#,
ĥDMZIF ���R�������Nk��ݝM�z��*o��wH������>��I|�H'U�[�e���������m㨱�g���9�TKZ��z�c���g������#��Z�캢��5d�i^���/�\f���
���Dv�(ڬ���ie/�<�u�f�!� j.sƐ���ȣ��w�%�<�����*�x>C[��q,�F��c��K(�Y�a��xk�І5���{�']�w��u;I�Yb��J������2�P��L�N��dщ�|G�ЎD���.�f {��v�y #� ��R�vc>^��l��Y����Z~f�PCLsR���~E�}	�5��~�4�]��EE�hN��y���	��_��j�nq��{en�k����y:ſ�k�]����9�f����d��B�5�Ǒ���`�d�a# X�֧q�lv��Ϝ�������uFs��%�T=͡In����?({j-��>(m�؆	����a� �VnS�B�%�d�d��bڹUb��e�CxْSl���>�!d'E�c2�.d� 難�I�7�;0{�]�C/��p�\;uc���g���boz��lbJ�9g^b4�dHd��\�>{���
�
	�c�L�����CVNV�3�O�b��"��!����A
#�S��1���P"$�/u�}�������B3�G�ˬ�?�{!��	�%R.�*V	�)�H��~��^���+�Y�.�A#��3tt�u�[�m�3�Y�_[Ȑ��w�,5����}�$�/��k+ ���Uh���5s����ͤx�6����UQ�s;k�Bd*#C!���3�R|{���I��42o�F.񟫿�����$U�G��헴�����Rj���G��w���H:JkȤ���/ϻ��y��r'j� 7���sׅV�9�s��ΰ/Yə�y�ѽ��!ד��5��a���]�-^���6���OW��q�u�/;ՄՇ���Myi!]����j����n���w<�K�|x8�5<�=a7�jB��ִ����/`���jXݒG�x�h��#�iT�ݦ3�y��<;�U��̦�C��m�������T�7�Ɓ��݇h�x��#���"��G�eAx��G�|��ܱ�9��;.��O�5�
ߨ�<^d�,Mv{͹�v} +�����Z?�l�����W�а��T���ݖz}�@����^|�,֙� ���zE����=&�DI�}����"�\ٟ��>m5��)d蟦O�|`�Z�u~��O���� %y$�>��{&V��`�ֶ�����I���R��������4�B��l6k�*���������זu¦ ���E�"Xg�@g�+��ϞQ7����vX��=��F��;�kH$�e�N2+��Ej���ul�I>�(t��O=�T���s9�w�W��g=�d�F�_|�6W��1����WK�_�^�ڿG�ZO��W4��]��oR�D���TB�Џ�w`j`�[�F�1�(I���_�d���.�P��5NL�\#���ƕV^��q� ��NUH�e�aj�`;$e��*�T4g�U@T�w�(�8��ĝ��HM�8��h/>_�y����3�o,��vͳYaJ���#&�!T7&;D�'�TJ�|%�N]=�7��>LX���)�5��־zͯY����ɰM�]��z�W3�����:�yD���}~(�ܻ	Qwy��1�7��6[�{�aǒV�Ts��K�����&��}e�;&��@e�hMY��-��`��������I�ힻ�X1��%g�)�cXPv�,wh��%���H��,t*	�R����s�7WZ/BԢ;�Z�,8��=R�����)'NK6g�|~ڰ��b��/������q�Kv9�gE)�}���N�X�rY�kU�H�EE��e���X�ɓ��N�P��d���n��	�LA���t5eGSp<w����u&�5S�U[>O7�$߇�|=l�����a�Mgd�G�4�ޛ8��}�����
��SW�ŘBc���r��}m>�-�3��]>��g�4����5��}}Y`�jY��[Ol-\�r*�5�#e_����\��6��:m�v$?f��X�7o���Ձc��`����茒|���������2��lU����	�҂W~����a�:�!Pr$���oL#��җ���G��뼴���R1�!zFI�y����{�����^\�
�]t,W_��w�wS(��ɡo�+����^�λ���DP��h��*R����O��X�9a;�>2}�6�ޣ�n��.s��'�Z��$����'��ƣv}��.�>�r;%ڊk���A!�6z~w�>�/���+(��Q��@B��wwo�\c�w�_IS(Op8���=�S�R��0�2wû���S��B��Q��v�O�a%���l3[��==I==GΚ�w����8�Aя�Q�}�=�	��ɴc6�ປzg(�gt"3GSi'�kϒ�m��;��m|�H|�ta^	X"��z
�Q?�G����]�z+=_  &��\��+{�F�|���֣������"�Ѯ�?9h�e��R���Z�l�����b�/����$2����� u��U�O������zk��╷��X��p8��[�'��I�.�U�
)__i�a$�Cdz]�E%+����U����Z���Q��/����7����&b����4!ډS?�>Z2�1�j��%����-����ua��8Z��Q;�Q%�S1��B
�7p��S��>�k�����2B�5Ӽ%=^����mֻ�ڠ���m?��k�Fϩ�ϗR�.N�+  Y��4�o/-(�n����,ʀ���f߿I2!M_U[S
EW���|���4.���b�&k�yd��x�
<���(3����o3B/89����F¯*)�U��O�x�4��{�<Y��$sQhm@H����aa���]��ꊦyFߴ��SM7��`_�r� y��y�����ͮ�J�LV`��r�+L�q�`�#��y��V�Q�F����X�j�s���#�M�g�^B�jJS=7��� 4�ߑ�fu~��	��}2Z+�>�KV^];d��F	��~�Q,f$��"�����p�{��,�Y����,嗙�b��!��y;g�a���)qf]a�>hs;����k�y��1����r�]��OR�+�M�*����*�MLgc����2׆��Yƨ��~�>�����X|<)����^�6�d�6_WM	e�b��b�PK���{V*Y)~�*��Ӹ�h���&�h.��J�A�U���ӢR��f�f��Xo���1��l퍘v��%l=uݺ��M��{�Κ���/�����ˤF��fVɼ-�("�*�Z��Y1��+��-���s��v.V5�08���TF���V�o#U�Ph)�K?���D��"9�I[����aסf��s����~��F_H���B�"F�r�QSi*�J �T�m��:�4X�}-ͼ�����i3�p�����%��dJc���Ij��r5�G����rC�*z����r�s7�Ɓ)����|}�ʏ�.���*K\�݀���`7� tǧ�#�\*��x��R���n3��7�E<"��\Y�-�J�2�O�hq�Tto�c=ȿ�nzƺ�TM��%�m�+�H������)�d��K2���)7W�'1���h�X�FDP������:���Z�p H����r�R�w:��.r��X?H��Cb��D6w�[��wv�i�Jɧ��3�%�5Y�L�u�3T���Ju?���wE@��md
��n�5)�d�n��b���f�D�_�k7�ޙl�;=P�q�oC��}��Hq��K�DC�Y�����'�qD66w.[�O��8�
�F�8FQq��9T�� ~�������[�b�R�G.�@V$/om���4�2#�E3�.~~H��b�T<^�u.��~��`��Ꞅ/�VP=O���x/�ߛ��'��U�`�'#A�B�i/��*�o��`�I���t�5	���*(���[�����B.�i�%�(�eͪ���5]�,��1�R�����ު��w0|\�ȳ���`���[�Rs۪���ϓ�� ����Z��Q����9+6�{�v��t�������B�uJ���0"���m������/��Ala�\&�Ƒ͈|��r���3�o��d�s�|�e�K����e�vC7"Z������n�߾j�}�����N8j�`q��a�5�yq���c�|B��@�Q�]�]��<I�e"P�XS� ���l��ӫ@��9��h��\���M9^.��s���o�X刺�}d?��pD�����	UU��a��w�4�%� ���o>�`;568�w���&]m���|VAq~=<�I�هk}�_BEܵ�q�|y�xHݭ9�;ʶfq	ǽ��(hxѳN�v����SC�%���\Þz3�;UtnǴ�z�/�:4D1��r�>,�N'>S%�4�Ы�����^t�_G�'��'���e�"x�苦t�)��o��P���Q��~��y�w1�N���u@=zuHpn�[;7�'BZiZj��>��%�諧�����ԨJ5_���q{��ʃ�$0������Y�֜U�	�o�s��76�
"����rp)��{���f�i�g�<ͨ����Es�wJҚ_��G?�5(3^�K�1*�	w�.dr6dx�~ٿ_���M�rt	��n-�S��/�v]��϶nOH�ڮAks��ho�z�R�]��ه,��{��*����n���B8��|�!��/ђ���#︤ο�����D�5�ҝ��%���䶣hc���D�]�z#^��_n,��A,��(k�wM@2���BZ�<,�8�6�w4�9g�������y3��j�W����T'�۳���᎕w�UR��,6��PuN�[I������x�}�G�eϨW�C���U��f��ֹ�,}4�m.�e��O�jh����v�^	!�H|��{%}D[��"���U���2]&����h�\
�gt|�J�jJ�u�u(���X�a�x��c�j`�OYQc�ֿ�A��/��9����8I����Xejn��T.���օ*[g]�lч0Qu0X�20){��m���[E�����X��ۯ�\*�ո ���p|�Q_n���������et���lNXh �XÃMR75�'"�1[�VbH=�G�����De��[<�-�J��̠Otӽ
����p+5�R�����*F��1;v��iy�kVY���jv����N|%n��U���ܱ�v�^�T߄�Z����<t����v�y��|�֡䒃�?.\c.8N:߾;��ثh���Ǥ��Y_r���|��.�'4ur�m��W�rP��T��!d��J��S���89$v�hr菆��w@C����FM$�D�v��̈����BJt����	�S��Dt���D5�|)��(g��cOԺ�:(����z`�輋��,�w� ���^m�F}/SQ��׺�g���nO�E@n.�V�:��<�#nX�5���v?yZdG�,'�ⱹՙ�;��,;/�ђ�ۜ�먳;>���!����&���߯0�o��EL ��B(Lhk �k����c��΢��ǒ,⯲2?�r�����m�#�as��Tt���-a���*�����"Z�Vk㓄 �y��i�҆�/��gr-Wb��0�0���{K�>��7���{j�?��x��A��ozzzv�!�>&�:�B���'���oZ)~h�<5�b�����������*;E��s[r�D«�U����!�gI����_��[h+�a`�M��Ьރٰ8a{��$���C��d�<���݁/�>Qf����4^+��zk�Ǿ_0�-m�0�ww��k�������,����{pׁ���L�9���zvQST�={�����Փ6z�CnX<���T�obgg�����fd�%�d�BQF�,�Ջ����WU�d�0�04@��#����i�\#�X�$� b�KH�ֆ⚃�JG��k�_T& U+��Ss'�m���܌�%L��8w(���ݵ<kkX��m1�����f�>Ƈ��3,+Q�G�ü|%�\���l����@���7~�ΚRd�.۟;/9��L�T�t�+ (O��/6�c�o�I4%�~��2��1�n� �=�$��A$�ǉ6�U�gF�iyѕ��:$�]�>fx��)�`ѷ�jC���6��X�����>��30�[qO|ơ��N����,V^w���#*��/2��[V���[�Ɠ�Te�o�W��{Qi�bرW//t�į�pl�L��F�Elu����`8�H�n�l�~�� 2D���|��W����g[�U�����X'��*�7��B��ֳL�W�˗h5ѝ$�1D���@4�" m**1�:�6���.�.��vM�l��r~2��C3�#��%��M�>���"�\M����x�n��dg�B�ƿ[��`���GеWn�GZ��s���壒�vl��te?P$I��+�Q�c�ػv��tO�q�]Q�H�JG]Tf���?$sl�QUH#]uM�@�k�{�m~�?ْ����o��n�xd/�q��&���Q����qP���۸\���FI�w�M���������*��M���- tZs�drUE1��:�>���k�H7{2�8)�O͂&�y��C�I�bG�Rh��i��9��[���A��M���Q�[ �@��q#
E�c�!}��0ac����ޟ��~|�j�H]�k(s-�ul���{!������������߬�r�������m�<�b<�F�{G� XX�g�hF?{3�*z+��K��$�p���7�.5@S�jJ�!��~s%\$��M��L���)�<:��7h]�iEGH��L�&Ҭ\>c�G"A���;�B&�B�*6lL<��y}�yzr��<��:�����B�z�Eid�~�p~����k�/E)�����Y�`��a����fU�G�{~���e،Z$y�k��R�v�&(=�f���ҏ�-$�rϬ `�?����P���7s}X��aJ��Y�39E��5�[#2FgU��˳�yy	�����X��'
�<� ��OU�?�<�Y��흉1a9`|C6 ,�5�++k��U�E�Hg���E�Z���;mD�k�Z�	d{x
y��X)�Q�����ѵ��}v㪱�"F�S��({���k���,�$/ǟ7^�eY,p��Ws5j"}+���j.�P��Jj��r�#>��L��jJc��ޛ�j�5��2]@f�V���܄�Y���4^�+��s�!B��z8�7<?�� ���Yv�T1��N;��BHܙ�x����7��hZ.)�;K �*���w�Y�>�%p��Nb�a�>��}������"�^����zF�|�}�x

����e�����P��uQ����S�^)���A�^:7��ȋ��u��ݜD+�y7�����&0>Bdk�Ν��{2�Ί��� Ye�=�֙�v��iw�{���������F�RT�9㞚V�0�!8���ǈ*�Z�=u�I2���y��D���E��%9a��!xp�Q���Qr��'���SX�p�=�N�]����J��
4ڲv8��S;p*m��L5���n�y[����2\"9)>|���~��ު�l��'�+d�b�����@7�ӻ{	lH�>*_��)�Z��'����ɲ�n��ZM�h�
�0�p��Ѯ�#?�p�r��cj)�8e~�΢�`�+�g��w�6k贍�7[�~� (�Y"߫�u�K^��]m�ӞE�<�����F��7�����6��Į^�]\0G�4%'��g�������|�p+/@;w��K�9�jw͌�jܤ���Tv^o�^c3#�\<5�{��9Xw�G���kX=.Z�#!o��0���c�r�P�J�+�cZPt��`�<�o3�_[�i Y:���]����:�<�.ss��+���Ȅ�c�g�F*I^��w���w/�5������!�IL��@Y�����qY��Rӂ��3�a�7�@y�G#��=K�G���1�8�ʏ�N}��ڢ�jE�ۿ|�s��t�r�7[zy��`��:��IM�
���&���ޕ(�1�v�!dp�B]�㼊<����γ��)�
�;W��'�`����3�����&H��"1":sGH��7��5�}􋕼#%,���+��W�]}�(���tx�[�5\.��[6��y�mv?|u+�dq,�=�����@���(%ލC���#Qv�'�?���l��9	�����'fΆ-
f��T�<���T�8�2��꣝q��v��	��;��b%�-`��V��4�摆r\q*Si͟ƀ���f",���1f'Mf�~%>BG��P_*_F�[�V�0		ڃ��C_�(�$c@Oѻ���u��1���J��)�\d�VعM������a��lн�c��n��~��������z3�<ͷ>l���ul�Oc�1����%�9z]}���h��1x�9��i�ڴ�CY��Y�'����h�
S�t;X��`@� Py�Ŗ-=��2M�'<�ˎ|Yj?�{V�t��wyx]��U����Μ+2چ#���O8�<�-�C� �ގg�A��^X����N�I�iq%o��X��9�K�a��lXD��n*��t�Y'��LJޢ��Cж�Q+�ewp�E`��$����7!g��|�\;�T��Im*�0(��JE����|�Lh�}o�[ >g�jx1}����7F�v��:��@�\���2��ѝۢ�s]�8Mi�+L�'��P������p��2�)tL�-�X�C��U.�^.lך;cR�5��^�TO� ����̰4��d]�h��'� $��Q���FRS�"���(ā�}$N9��n?�C|�o��+��ܪs�G�gz�����ܣIP��,248 ��3���:�w�Q��X�Ǝ�m(��i+��y�M2E;}���@��)�����j]g1�U�J��!I��OK��� �����[������_�(�!���}��U��<�b�3�����N��J��J���֝_���@E<7)�V�$t��ԶzV~}��it���p��r���l�^�3YD�����>M�����1ce=�iTy�|�%/C��pOofS��k�O�kQP�'��L�$�A9G��c�Q�xp�����	I�bk�;��q�z�D�q��d �P�ԉ��� �Yo|V�������!՝W������-=�[Ѡ��~5�xm�rA���T��1��7���|�yCg��L۬�7^; <mA��"�]�vsL�����^/���P���d���|_m���^6g}��P�)I)yۗS��,���;s�q�V��k0roy.z	U�y{,�6����[ᴢ�:H�MD�w�
?�x l�C9��R�����Z67��;��Q�	��](;�����4�'g��=�8*hW[�X^h���g�M1�
�,�W��$^����m�;��y������V�b��i����g�!-�g3�<k�V ��T�6���JT��t�ם ����W1�d¾Y�Sc�Pb����XU�58k�Đ&���V~φ��&N%	�n�3�
?v��Lެ�/C4��{��(d�V�y_�/Hk��
!����Qzl�zsDO~�D9�	"Ĵ5b�C�%>oFͧFf��oknC�;Q����]_��]���?�~�l�r���&��&*n2�Q��ܴ��/���N�l�N�;�7�;QQ��ʧ�¢��ًE�x�,�E�?z�s�z�&+�O��W��T���H2�X_ip@�yLoq�7����a�����ud��}Io�ފ��3QH"�
��䓙k0Brf�l��+����J�ڡ�U�t(ڣ x��r���<Ty�>4ke7O�*9�|�m�������Ks���AM�<]n ��G?GǤK����
�iV���4w��Bd�m$�%�·c�#V??�A�06@�D�W�<��z�8�;�l�^��c���xwIVL?8RUh�\�F���C�	�i�̻H +v�EPo��C{V9�!�hϒ���3�5O��Ms{h�ܷ*%rʅ�r
��q}�p<HE�G st�#�%M%��9AsH-� �P�����u�u6��q�&�zck7�3��kp��:��N>~���e]��ae�����?SbzBg��l�aՉ����9a<��,��`(�! �Xǐ`�aCg@^�R�꺊�o�h��Piu�7T���R��Ʀ �֜��f]�`p�sŒ{w8V��c��K���h��g��;�.Ӣ�x���������duQ¹�b����.�9���K�����nN�w�\1���^��p��$et���Ol��iJ���:w�z�D�퍫#S�ʩrɋ��OY$�E���3���֏�������2�)�l!C�D�E��e�~N��#�XDR�&��0��lsg`(�0Y��v������y2�a����n�����cY�߬��)B�Q�:�1H�L���V܁��h%�zbƑ�C/f%�Q�]_�N�)]���ߤ�D���X\���&��ap�e��qZR�+�َ|�c��IS+Wט��w	T�I�o��c[��n\�ܿ7�P��\����)7=s�i�$��ņ����:R�#�z}���cU��Y���3e�`�j�%b��ٍE��œ�%�Ph=~�	�ٚq%2�x�����������q�]�T2F�=B���F�in�Bw���/��E&���C�������FD.��ʂ���yW'Q�7��T����Qd�T��}?�Ɏ�TV����̝���]��Mfw�*��7zl4N���^r��}�_�_RY�Zn���ʽF�#��Z��	��:{�����T�m���W3�>llz \�ËyB�PM��q���[���j��|HxUS���(�^�bq]�f#a��ฦ�]�փJ��p���[��ꞓ��obI�t}�[�qƱ��:]���y��N�T��M��ȇT5s�8�W�f0D��TG"^��܂]�v÷��Vb�#cɆ�B�X�!�v��M������>�n��.b��..����۾<�P}\��A>�o��.PX!z��u8�^�����pA�-3�_��ޓ�{%b����h�X]�HZ�W�uuс\X(�D�&.8��&6K��}&�?<��Q�;�FA��5Z���=E���[����x#�|�E�����(M���_0N��$Ge55�,�cp7��^��N���^@u��N�����ң
�����+��:<@����O��6I�O?�PN aUɨo�z�����1�̠Y���jv��/��w����L������Hf�D������_��7��J��C�ߒ� �$��Ez�ݰ��ml
`�*'d���ͰY�b�p0��'�a6�4bڴ�#�n{J���(��҈\o��۟��F�ʴ5�|���"f�>]���x_���,G}�'�w�"LʝAġ���45ɑ�K ����[ӝ�v���z|���(�?��  u�3 pN�͞�ҽ�D%�f����S��v��h0�,��g4��br��O�ˉv)�7V�2�Go��gh+T��,e�,�>%a��(���� I�`��r�:94��l>aֈ���*�s�Q�_����e��?�S��Q��ce!&Q�bd�AW��K�'�@������Ҧ,�q�=�g�;�-I�Cz�n�npNQm4�ѱ�be����h����K�2�ew��L�UI]��@Y�`W�X���� ܴ��3��;�#G��I�*q|�~6zZT
g��.Zp����J^!sX2�� �����EIH�ƛ�qB���$: �S
#�����K@]�o�\����G/��3TƜC��`Z�R�,��6�c#���DCp�5¶����b	 �wj�2t�mm�1BZ_�1�Q�� U�;_l� g��� M�͔�s!�Fp��3,�U���4��+vOs��xI�f}r����!�m�\��//��=K��d]����u*ȳ����۔`S�-:<6b�7�b�Ѓ��h=�����	j��O	^�lDU#84��O�ht�7`?7��;���/d_7����f��Y�G����S�	�*
�K+������ٷ97�� �<�k��-^zX&�+��edU2�)�y���ۃ��n�Mn�XP@�Iձ�ZQڝ�����#
z6 �(��|�����,64f�tƵx���P�m"�+� D��Wg�oN�ܫ1�X�Q��S�I���2\͒�&Z
ɀ8f���h~�\U����ɸL��{�D��:�O�!�V�r����4t33N�������E�d��7��q����N�1cMNV��gtΊ��;�Ȋck�����X<�ɨp�u�9j�|�|3��
(�#&������\Z�&���*z�{W�	h
SR5� �37�z=�C��߈�Ŀ�BPA��r�-[��g�W}� R�	��K#J�\���<�{����L����l"XL���_�됏�Ȓe��C׻��kl]i�G������M����V��"�r*[_����l3�yt$Iy�߲pBOG[��� -���I���ޙ[�/(��s�t���=1��ӝ�v�8��A����4쫙� eCw���w�9	n�$�=$��yk��RR�E���DL����s��la�f�JWG<}F!v��wެ�ςH��i�ھ�;o@*���r��Eq:����B�m��9���f,�#y ��"��V�Z�(l�:�$&<~�[@;�&g?����O��j7�;�Lⶩ(���U~�l�������J8�sb���EL�~賐�?�j�0�Ju������A�8�����o<�r%ȃ��A��8��� 8�A8!3<7����-���q	�"�PR��������3ɦ�	 ��!�6+OP]m��@��Q��|F.1� Gu���H�������v��`v���;����-wޙ��d`���΋���z�Z,��A@�SU�vLZ�8�*豲�%7&~�;W����{���hw�?��
4�K[��6�ԫOn&5�FQ�~3[��NәroW��M�fC'��Q��vތ���������c�l�>,	dh������ig#���}��>��y��� 7c
D�$A�k�Cb����>�?���vU��m~cg���@���be+!��P���r�Β���DWO�"��3(oN����2%t�̬���	�@nx�u7Vo7 �(9I#���e�� l�?ZAlƫ��I��Dʮ�h
ШQ��Frn���z�F	O���#�þ(�m�'�_x?���]8a�xO߱������ko6�--cݿ��MǼp?@e/� ���/,�>�C'Ik_�}9w޸�����P�ے���_���oRW�������B���}{���?����ЧJ_pc��KJnq��o"9�sq��[i�Z2u��������x��(��$͡��y�*񃇪z3?Z�D�Q���۳�D\�4^ha�R�����1��Rt��O��O���)*����|�Q~�YZª;9P9_|�t�a�HLM��R�����ҺzAG1�-
Y�h��:M���Œ��!�%_�ð�F��F����Z.���7�g�������`Uw3|��z�����nn������Ȏ�N}��3e,�ׯ-��J�����} �1_9a�T%�ЎB޴�X�z U��z��&Z��� ���m��F�������䔽~�u�W-�M�?�a9V&L�E�[��py�ǂ�<`Cg�~�;��r��Xw2'�b%���w��vuWO�W����6����!AI�P���Oo�ҟ>o���꽧���mNɖ8�S>��y�Z�q��x��nB^g�X��?�Иc�|)��#���,Y���!��������#��\��"���7����w��o�P�2�r՛rםz@͹�ξ�ξ�"I`$�&J��L�f}Zg�(���b��P�;��lfhzS��
}��y�@��c����;mǕuI�$�
��9}ٗD�P����Z�~8�< |�u������z[_�]���4�|�_�gb 01��G��>��!���+��ss�	������8�����@y���0(M��z���~K���B�MD���%��c80���3΅3O��;n� ,)X��e��?�ϨXRY$������^tI<
��n�H>p�U>�m��˻�7��Ų1m�A�ii�����U|�U�s(����ƪ�q���&A��j��ȵ�=�����2�5�ԓck�0�DP)��!���3�³��r齙|b
���0�X����J���}d����,��gߐ6"�$!��z�D�&�n��c����j�Px��"�P׊@z���W �u0�%�͒~{���*y����|n)����ye�q�_�C@��*(���ϓ��W�z,|�ϔ��إE���zrd�5�#���%�*�9˫˳�������M�� ��h!mh*��m\�B����l��O��9+;�'I��=7�ڹ�b�#��og�'ꦟ��s~j�j�q<�2�$�vu ��u��#�k$�&̉&*�x��M*̼sS����^/T�`&��u���mw�������x����jѮ�M@m5 >V���d��%�� q5q~����a�l��5��re/4���ss������1�n���5��kH?-����ؒd��9F|gd������ׇb�ѯ�k!�s�yv+		���RZL����n��c������5_�7��4;��O�h���o�����|�6I�I6
��O�-�$�Z�o%z��twd]����mk��.!nK7o˻�aD��Yxe
N�9����TD�Z l9�����4�/�y[��'���t[�����*�]#����0v�e�n���! ]�*?�R��(��/8���h̢��F5	��2eT����ۓ�ӓ�X�%eE��:�<U���l��LT��毁B[��%S䶳/9q�m��m��H46�4�1s<�ڭ��2�Y���Oz�|���x?.hh%@*}�Sz�K�	�w���9٧lIP3�ng�����8����b��:�JOW�&�*�{�$���R��\^gv��9nUʕ]�r�]ڥ�m�d��ˌ�:1����iX�%lw���>��a���r���a�𯘢`��;t�!m�g�.(�����,�iܣxP�F�r�|�QNW�I��
�&3zU��D�"]r��>g�5����v�^���=�w���1�~I%V�=�M/��{�����>_d�*�ZCx��BdB`����˝�����y�ň��w8�2x���4%���)Z�P�nV����dN@�,-��F�v%��c|'2΀����4Fj���PҒs�s�HǛ��	nt' �U}ᄑe�'�8v���XZ��[}s�����6��î�p�:N�ڂ�Ԡ�2t%3�z容᫳J�ɇx���������݅@��|��U���&���\�:Ǟ1��[�O��*߰_��	�[��Y-��3�2%�f[���zz@��9�LO��e�5�X秓!X�E軽ݯ8�t����'����[0� E:?!�nk{G��g{:[�x��1$Pʞ6�L!01�:����"i�ՓE���O�w�q>�OcNY�hj�gn�MY<�d^#�N��{w,��tn.��xiMrq�,�yˑD�s������e%��9���괞��7����j���Qd�ԃՄ�s�Y�N#�*�Lv[T��?
�Ny$A\�b�\�81����;f�����`���]4�|j��'n��y���Z���º�N�����A%#��W����Ky�h�d�z�����;?����kw�1��1Zg�OE7;��&�yy����>E�lT� �_��(J�?����wKB���$�V���)��������K
		}�h�(��$	Ey%u�Ji��c��T��^��O{V7�q���J�Ou��}��������u�,U�_t3T-�Rr��EL�;+K�g��''��Mb��L�Y�2��;~=Z��:cE]��)G\O�3Ͷ��+`�*K*%Ӝ�;��½���3��e)b 0m'e��J	�������$���/��FQ�-*���Cr.a�P����L�������ƚ`q�����~I�o=n������_���O֮C'�`��Zr)�:&IjQl��?w�i�c<HrP��&W!mJ��*�p��ݟ(e�[%U��U��]Ŀ����Ob�2G�"�rj a���ʏwp���HY��޹akf|�ػ�Hn~�x�]��l�5��3�L֏s�"*Ă5���I3��\|!�]=�n��n�=w��r�����9f�v�'����:�MK�n5�V٨E���V�Y��p�B}��5(��
��u�E ����J�$%,Z��+��x�������[����<����,���F��ح�@��ި]���ݵZ�vN���F,��m�b�j��D{ڍ�-OM��y:"�Ʒ�,?�.�BR��]���+��i�� �	��X��>L���c�R� ���9b��]�c��v� �2��8��͞�3FH�u�{�ȳ�`���x�Ku@�[�� p#���4�2�䅏Pm�M�?`n�=>���\�u,~i���y�__F`ܶ2S�
k��{�̠��KI`�+���ʌ�p���`�S`�����BX�z�Xw�`g8c���9��w\�!�YA���3�X�n�%bI�#�����V�(SJW������PQ��x��*�VQ&x#g9r�,-�z7�y�lgI�`�y��4���U�m1%ٺ�_K F3���V��7"�=
�dP|��;���9Ku�FDY�j[@������ƾ�&���
����n��h|����1�ed���Ϡ��"����\5ؽ����ϼP�V�s�f�5I�d�Ȣ�|S���R�d]%�T?�^���o�^��=��K���~��C�hbs��sx��폅�6lM�	��&�]�?#����'ሪV'EFYD�[�Xh ��~�e|��~*t@�,�-��Z����;��1;MZ,PP�I�Qx+)Χ��_w*��F����<�".�V�0�VI'�:E�:Ȣ;Lm�6���t3N�Y�Yv�w�.R��Oz�����Fh�b6��ez5�(�dҟF���O�٣�)^Ȥ]2�M�w��S���������\��dE�	�|v.V��^I�R���S�`�T��}��=�	��`��0���@��6����<�օ�2� �󎈥���! _Ԗ,����=��Qr��Bn~�)w-|�+%a"�/!�h#��<?F���c��I��lb�̱Me���f�E�w��k�_� ]�p]c�w����l���;�'$
p���`�G����G��# ��1��\[��V.��5�2����v&�h�|_�3�y��V��%i�����ܭ.sS���5`٢�j)&O-yƤbc��6^>�ƣ�J蟺R~n��Ͼ�*bZ�d�tA����j��&I����B�:���QZ�`K�ẗf���Ce.�Ub�CXf��Շ��i9ME�˱� �n�v�B�t�� 9���XTTI̳�6^�({�o�/��H�[\�X���;�Ê̋�w2�?'����Jq2��@G~?���j��}-�����t��3N�J�_B����;�D��-G��nȋ���Z�@

y�]:#��_
�(7�b�Z��ǡ�]��L����MB�P	^۵�����z�%t' � ���x�K���K�ǐI�´'�tޥ<�H�OI�}�Bhޜ�B�"G҆���]�ӊ٩���R�}�]��/��8}G�E�A>��+��R8�>����o����'#S�T�N�.홭�ߺ���%mHQ�(Gb��(N�J��^;��@A{i�tm%~�_���|C-Nk)~�6�Z��3r��>��R�-m�a\���$9;G�3����5@#x���q�*�&jc73�R+dy��@�`)�݀�f�y��V�$6ܵ?�y��6�����&X�`|no_X+G���Hzs.'��0ᐢ�ov��쎲˜�	~���M�����^Y[�&*���l%7ge�<�?J��H��Jv��c��Ί��q�i��[b%��v����ҽ��tqY��X�fPJT-��܄�.�a��
r�e���O�e��U4�]�%�6+�^/1������lY�k�����4"��?~������jbt�UyT���Iq����<2\���x��Lޠq��X������ӓ*z�K����� ���a��8�n���'s<���s웏��<�d�m��p�W�D-_}�.�S,��Q,왌g{{M4�_x��-p�5jS�y+M��g��u������1���1~�{Z����'��S��AF���ȧ��S�p=p&p��.�zy��>y�c��]��ZCB6�C%�����J Ko�r:��W���\bP���e�F�+qe�Zzs�W��f|Z�k��\���>o$֙�<L���_���Ѹ]��'7�J;���9I�6�ݐ�g��mV��S}�6��� \aX���h*��s���L��� ϚfK(���[��֯�ˉ}Mu(��+�!�֗�!i{������T�o�y�7m��CNR����9�ձ[��a��HT�i�8�s/M[��e��;�E�ք��_(W\�Vǟɲ}e�O���������Đ����ӂA�T��$��c�^��J�\����iJ_�`:��;�Yp�h��hvN����V�(A��5��W�pX0�\W��z���BP��y��Ǧ���5���V��#�8�D%���i��,�|����@���}�<��M,ɣ����|3�u#���� �3>���ު\Vܾ�yԞ��嚱�U�J)F������:e�$��?k��
~�-� ���iI����z��Vu{�(�1���daq����s��k�Ka5����<P�ة���r'��}���[���WʭU���RB����	��$O�m��r�?�?�X�B��`;2�_�P�Ǉ%�?��	�b�HRօ1��sUC��G�4���X끮��1NB�2w�5��'������q�I�/x�x�~:���o�Us��M_�BJ4�x�L��,:�Je��d��D��[,8ͩP��|�i�G�0����X��r��y�/ðh3��L��(Bj��r��Pծzc��%�/ߙ��^i���q)z�d[ݺ!3�X�(��?|i������v{��5���Է��V�f�9/Q�54BL����!P{P)��a�t!f��r�[΢=�`'����ߚYl�i��h���1M��ڢ �9�)H���Dz��-���Kne� ����>J��88~w��o����K�M��%w}�!� ���� ngy��߳�#{�:�c5���I_t��݊�	`BGdW	'��*��I��̋m�j���L���!5	]Ԓa]D����#-�;�Ķ�K�xp[|-H�ME�����!�֧�������c�Ƀ���M��ī�M����ߦ�B�A��`�?Ϋ�c����t�m��Ŗ��^���s�͖X�C���$r7lo{�Q���-L:���Cќ;Q�^�A.ڑ�:V�jAړ��TYABT�/�T�8�$�J�+�o�i���boܵ5�Pܨ����Ҫ=�����]T8�r�'B43ӧ��{�
߂�3y�{B�S%����15��y�η���[��ݴ
kA��0��ə�`H's5�E����d~xmq�Bm�r*�ƌ�	���U�%}Oҥe.�`�:H{PGF1�P�d{�9�4S�a*���tq?zI�u�)�I|�|���ҡ��Ү�/	�WIn�c��d�e��{7�}eڥJʴq.:���C�v:�ʭBwǃ�(�
���z{^YK����_4�M�b�L)�c8Ru; ��r��a����ۡ�lG$j�_��|w(�3#�?n�]��~��CPy�^;8�Js��溊ǄNb���Ǭ�T��sg�>����6z���׹%)ч�-������cZk�qQg�x��S�Pﻺ�:�l��RRu�Y��Y��M�b��X|�J6�hW�n-:����[Ndt����ߢ2m��)��*�IO�os����zF�S�����U�$��Ų��$�n� �䞍՘Y�~�e�Kc�����/f5t�Z��:q$��z�=:�َ�r��I:X]�߶/�a[7�P��,���}=�.��_��
�ڼ<L��u wz�Y�q�`� �G>z�HA��������ʇ}��vh�c�X_�"�8�sr��)��[���zm�4��u�x�W���6Iԩ�\o.Ә�]�<��ao�D���s�z��+��-�ĵ>�̑��D���#'�wI��6umy����K�5����.����
1Z�K�f,�J�7J#Z���P.׿�:� 9f��A�o8d��U,O�n�[���T�]�����$Z�{���K�G��>j�.0y�M���{��(
��������L��,�W�JRO!.��p.^���:�b+��$I�D�G��=J�����0�upo{T��;��>b��?+]i
�BZAYj~`��m.�'0d�����x(rWX�=�e3�a���?�b#�QJ�+���I�pu	��!:�Y4�l���8��bY��|x�1�ԁ������aEܾEdzHN��202Nd�`/�OQ��'��s+=�:� �яi���ۦ���I�Ũ�hd�9ګ]K[�s/~t�q��B?d�킗�G`�vܩs_[9���� ���f35Տm��CGNݿޙEu�2ԛqm¾�s=��YB�]�����	���J%)�)�<N�4��0����σ\����r<ʟ�!W;gÞ�ف)iZ���u��p9&$�D@�Qn�y5s��0����{%95�Հ6i��O*�a�i'lg�vV]iʔKd"{�F�>ߙ�E����[�8��Eq�x�eH�/������߽��"u>dfu�Ⱥ�T�o��c�7�Ht5�|1t�5W�m�׼�4�T+S�U�E�ojx���X�Y��b�U ;�5ݣƕ�̑���؏M��r���#�?U��v�-�Ę�j?}�Φ^]ZB%!��LMـ�.S���K�O��9�VYk�e��%9������5� TV��b:ͺ�<�A����M�4j<�������
8l���P2B:$}s�\�f���p���� �M?ڂ����S|�h_G���"3:?ny���&��1s��M�� [� ���ZT���/ېV���0���L�3{Y��!���b'�X	9��?�E����0|+�>��*}�L0=��x��pJMg�W�b�S�T������s�6[yT�cuJ�>';�� ��U�9��[[�8�Ki6M?�dHY��חv��Z���&�P�����p� �O9��ah�"0e�F�Z�B�����Xw�"Ɛ���e��JֳDLW4֍����QID��Q���4�X��i(�W��/ɿ�V+�J�Ȧ��] u)]9��/}YKus[�J���.5�%��X���K4	���6�ҟs�_���b��L��f�Ƹ��s�7%�3�\���-<3�Q7�g^w�Z��whx�'����>��/��L��Z8� �9U/vz�=;_ɼ��5=��a�g$~��k���yHPCN9Hb #���^��[��sM-TM�d@��*�:��S�b i�)�L+�lX6��eCv3
,y�����Ks1P�1 �<����1޿8E��~l��v�Z�ޫ�V�F���,���nn��XA	[���~P�EP��� "&Ɔ��)��v<�C��o�[�>�i��\�08s�Z�d0q�[���V��=��q�A�>��L~m�b@����0�h}@�!�{����>�?�q��V������?"�Z�]��.�|���*z)���<$g���}ڮn:1SWo�����h��D�X=e'�A2�`�`=�\}��0�Fu�D�n�W��❔ڻ���~I�,�k[5�
53g���C5� *���?��h�Dmӑ��مk�M��A>��π�6Z��	UӺdJb��!�~��7�O�d����sg�d/�HI$�C�y&Ѥ�0���0���&�ၣ
�)]�ʡO ��~|�|�lnhr7E#8�H��B���=���P��%P�Lf��?��`c߁7ڄ�_{
Ų^����%�&���k=���tʀ���G��!�Aq�����3ZJ׆�M�
�y��'�D���Mƪ�S�Qj*�D�8ev�F����c!?�2�z�)�H>a�co��:s��Mƌ����������V�}
R�sF���`�DW9�耿0i�a����9Et�50XDCmՍ�=�f@��k�*��Ƿ�:��;�����c���׋o�]|�<���M��i.ִN5=A��D����CRF��v_9d�(�V� �N��:��
���>���<�/�d�j��9{�����T�8��(��K���S_<�P��z��;L��}-����)�-k��I�-X��Qu�)�L/��g�^o]��7�\KtI�Ȑ7'�H6C>3�<|uTT��7ݥHJ�"����%ݝJ7H��tww�t��=� C|�{����b�u��O�b�g��na�C��ֿ����u���f�S����k�q�-��+S����cL�-�Ͻ�ou�03G�}d�A���
��������=2P-xG���=Z�qj��V�A�q�� [^����&xz�s��M�{��%b+!�,�y�)��73��?˶�L�����_�z�A�8�4�z�S~w[��wVnLȺPͬ���뤗�4"����ǲ_���{�h`UF���Ǻ_���t��c�%�9����p>���O���ވ�yH}�����Zle��h��݋�-��fUA�HFX�m�Đ�ZJZ����k����7c����X���`�)J���}��|��y�!ml]���}�dE5�����d9�~ܰ��Z��Q��0T	'�'��ū�Ќ��A��R�[�k�p�B����S5���<|u�}�c��KG\��q!o7�.�������%�D�j����� �6����o!��9{��?m�W�L6r`Yw^����G��w�PJ�dq�VR�w¯5�ߠ����ƶ�S�]���R�E����}��\�������������a^ iU4p�"*#��^�'*�C��P�{4��*��&�sPб�g,.��G���SI��o�\d~x�Y�Ѳ�ӷ@��u���u��t���6Љ���J��Ǧ��I�nnZv,��[z�t��O�!��m�����4��}w[Ւ���^������m+1����c��"���Y���H����[�X��u5GD�J�SW)v� �w�ġ�a�4��eB0q!}��׍�m� �fG���R��bV�.�2�:��N�{� �VЖK��WxN���H��������[�$���-�<;{<��})�^��*zt��ui�Z@7��cW�;��J }Ԃf��a�j?��p�q��~�/lS8ي�J�:���-�@WBZ���.>T>��|w;�<�xi��Q��7n�_�>�Y�P�������r��o셦�x̔Q��Q@r����cTg���Zk�N2D<9;�eI0x�������gr���C�H�Z��$�$�܊�{k�0솎e���@f�a�O/��Y�T�5���Ym�7ox�|�t)G�_wpm�`ۘ����j�e���1ӧI�KC)�o|�����vuI�D� �$
\�o�7����|�,�.�t�6^|��G�kya��K"4~9��"��b\3�nq8�k�w��F��y�����
F��je�W�TcYxyT��3�"o���6�+&T6-�����j�\f����$�q�=֐s./C�	�+��Y�1�S�����lj܎X���qj�F��0���q�rj�)}�҈�1@�	�x�l1x�
��6y����))�9��7u8�+Ø����'�h�Y����H&*���1cv�s���s^$ۉ}�M}�
��
���r�OIX
Qhl~�	Ǿ����I�ٺz����;OM$F���m������]0�C0)�, ���Ϊ$�:��� v+�y���\7���-��,V��0��N[�p܍�[g<1�`��/n����b��潁j�-��`6x��i���!��#��*�+�\�J����>_��i���_7ў�^�mXGѥ���(���ك��b�o���\�(I�+�W�U��4�٫�tNC�n�Z�}�����׊�N�M�A�z�w�����/7�	y��m:(g�$���,�'Yc�s��Jb�M]�R1m��A�f8"��Y�y���C~v��w?�*�M:һ�����3#�gk9�%S��L�`Hx{_��°����t��6���{�KV�"���,��e,@�m�f߁�s��(��_I���T=ED�N�a=<<0��>-ko��!JL�m�yB����-G>s��(Z�T@��T�:|)㼍Nϥ��<a�y�J�&���At�k�8��#hr����i�ݗ|݈Js��ё_u.j���aﳿ=���mO���fc!�i��+�.�X�{��W*3+����= ��sՌA2�	;��?�J��2���<�౐��wVM!x0�ܞ��|��U������}<��9�K�����MǲVX�ĨQ�>�ν?$������! �|M�ŏ�����߷>,��[�Zq����\g��J������(�;-��z� ��?y�u��"��z��
��:b�8����|���pf���mJT���9Nk�U�~}#1����������T�d�����b��<��>�=�%�Ɓ������T�`/���_a��EV�f��z�<�Z��uV�ҡw�lc)9��Q�Ol�?o�Ř4�3��|H�=И������3[WX�!J#��o��%K)Y%��OB�����z��͇�Y���ww��1Q�`�+3����򗔦�n	q�Lac:�d͕)ՙ��Ѣ��9>�fH3�y��S��W����h�nwh�7����M�x��t���g��T�n�j`(���n�t�3S��U m�:Yu��^��Vڣ1�8�F� �de�BlytC���NȬ���s�����M�]7d@v��6�>y���R�a^My&1�b��S5�k�魽u�&�g�^�p��L�ܣ�p2ѱ�ʵ|.�b���A3�;YE__�Z����V�7;�6�Q��y}Sd^�^�35'�F0:t<sf#��ْ�����]�s�B,��2c�h��B��}�K�s���̬J8|&�&z�d����ZYb,O,VЙ��RW*g��l�2�0����pԅ�:�DyV&aֿ�t2��$C������ό B�׷�L4{#�<�g��[Uu#'~�Y�;�N$$5Q�v�tߎrci^�k��XB	x~#����Ey���lsrjS% ���"Ñ!L�\�ŨRC��&�ź�֨�X�bY�?�u5zG>���L�Ͳ��rA7"n�̨m��}�k-)�z�ٌ�GN�tft�|�ћV�L>VZ��<I�Kw�33����ɒ�c�!��]���B�)����_��!v,���`#��ڮ�E��XZr���_�l	1j�+���eA���sZO�H" �XW��"�_��I��P�\��A*�Wգ�����J	JK7�x�!���wOu$�z4su4a'�ؼ�i��:J}����_�!���)�t]��$5qA��O~r��fܾ�5��
�l}~L�o�<lT;��+�t\/�0���t���t�����i���	D�[�����Ybs�+I�4����=vt_8����i�p�m��Q��B��b-E�')
����2s�����V���=��ϩ+lV��D�O�?n���ҫ�	���&��\<���?�b�Jß)����Ƭ85a P\�!O�O8]Kj�9�2s��6����E���M7���p�"�2|�W�h=w[��X֝�-ꠎ��葜��E�ne�W񶸜��sۨ^yⶐ(I�,�S~��9��z�, �����o=�߅�X��wXQ��I��f�b���0=w�	o��������2�l�>�WV�C4��3H؅��Sڱ*+GB+�� 9�|�-eL�����c��d��b���U�i|��ļ�ʏ_��m��Q��A{x����IBflS��8̓�k|C#(	[,��Mټq]�/;�P��қ�j ����Bf��Ժ��~��x-i��ͧp=���>9�◊'~�<L�6�1�(s>����R���+u2����S
�t��)����L����-�bH��:����+�QRWǮ���^������$aU��Rr�0Tk���2ʶ�r��d��d�8�i�������9�ҝ`��b��:����"J;q���(kszh��hy���!���[��]l��/C��X� ��*�V9ꗨ��rcy؍[����`����=2X�b���-���D!਒��߹�1q�I��h�X��/��a������}�j,+�mb��a� �9y�Vj��'�D�F�-)�xf[^&�����'�Zb,�bt�32��i��0֙z�]T@ފXZZ�:�aW�[�:��тo*p���*�*Wn�0�y�N]�K�:Ͼ��)�2m�W��o�f}�s���Z�w``���6��ɋo�v�hT=�n#�6����7W2S�@�@��p�z��	�{�v�}߮�'���ǩy>�����`� Z	����|Ӳ@̎��{�,^֢��?E4�ɐ���q ���')[Wm����#P�)�x��zG(j�lq�l�$�R1K@v��5���,@ar�??>�(���A6'����dJ:�A�jڔ� _԰��vg��Vj��R�A��篺���א���KK�儲�md.zS��#y�m+�O2D�#z>���UM��*DvA��j;�������X��w#ST�����]XU[�棦��`Z�����i1K��t�͛�'�E��w�K�ȓ꠯�ޜ�6����`���Aq�ρ_^烯<"�b�	ȻKr��)�ë��Z�j��ٚ�	`�F����o�U��p�m �m���Nչ�_�Y&�?���B�"���U���Wަ,H��`%����F->Y?]}�q��I
���U2A,��I�5��!���ӹk
��7<��a�#���cG9�4ķ��M�{�$>G���u#�Y<��w¶���h���BE}�J�B�Y�@��� ��cc~�U?D�ـƾ�Rb����CK�u��ۧ��-�^����V}��8$�C�����w��e50N��Xjdx+��v����9BB�/��&��,��?�]�����K"��Xqn�]'z}���,�[?<��"���^@S�r��n����{�`� r��� ՞:E�7�|Fs�˩���*��)��j�m�cw��?&���&�o��B?,�9�7�c��Mdۑ��\[��T9�Ü��+2��K���Vi�ݿ��{�NY[\cB��I,���c��ק3~��^_��vޗ5
��K��e��Gxٍ���߹���U䁯z�7��`��_t�1����Z�ɬɺfJ4-Y� �H�Lyb��3wE�t�k�-����A����{i�Ƶ΄��(3�TY9�Z�xN_�\}�Z���3�����F��C��̍���|W=m�'�V�<�oL�UR���A��}FqbV�I'�3(�y3�ti�c�u�v��GE	��8�G���}!ʖC����q�� >�>ltU�9g�N�{����<k�&����]���.w4��
���S�%�♻���܏��B|��\n؎�o�o$�O����!bz@>Cf���<��V�B�g�NHB)e!�g����/tpe�ylk�L�ȴ��;G���l`2�6-ޘC�1D��[�	�r�X4e�>{U�������E�sj\M45�k�KE�rk���������y�*MrD\�2����ه,1��A�X���kL{e/���9��8�E���T����4�tn���b�S3.lG��vH��q��ZDX77��Ʉ�I�ε�"(7wa��d�~���>��M�Q��y�!���`b���U)g�����7:�ܦ�)�K�@vgk�J�[FVo�=9^[!&�7�#b�Mn�G�pL��N����i�ʤuΞ��rJ��m/�,���9�A׈+	�D���Q�%�����W�ٿ�W~{=i���.m�o5���)y��xAڅ�+|����S�N��J}=*&���7+�yz�@����]V�~2��Q+����2H�P:�-9On���U�4�w�i�ǋJju^n�U�3���Ų��$�Λ#,W/��3B[Oy���$�������VC\�rJ���V��-tW -�ZGB��:�����!���t'{8Au��ߛ&��1����n*�Z	G����
x�����.؜���G%���b`	��9}����w��|r;��"��
�z�p^/�B���w�b���*�uN'a��IvM9c�;����SQ}C��f39�zƎ�I��_=����.	qD7Sպ�fTtUa������mU!|���Օ��a��3D��z緒T�TC��2�������P�����m��Iz�
俅�[��I4Y/(�ZE������Y�4*�=����4����f{�Dp�94Ց��{�ឮz���HG�����r�l�͉�G�o�\���1xm�^�]�MוɊ�2FS��"��7��qR}݌pX�ky���2�����X�G1���^[�'�f�7��V���W�����,,t;E���\��=-W��mmUk�P,}�Xv�y�*��RW�Y�����\��C��Eha�~6g��^�����3}�>�ȳ��Ķ�oR�f�}�9N �Ҁ}9k�lLk!�V�M�w$}�Ge�DF���J���L�G�k������C�FĶ`�:���[\<f�{&�ݨ��J۬Rך�~�^�~^�>ov��CURh?�ʽ�K6�Zz���e��M]�t���cǇ��+���&�$}b�ϼ?�?��c���\���&cFFG��Jp� 6&��/<�����O*��3u��Hő�|to�7РQ�]�767=����\[]KV�r��+_���qC��c�N�Yk��:��g�1F�ot��FY=����"�������)�Ji=0����LT	g��x���$���yyI��L��"04[�2W�?&vg-�(��T�֋���������N�R��Mۙ0}���؇ �i'\��P�a?\f;M�LkՉ�:�����
W}�qKh����67��R�������h"��p�X�����l�W���P=�n=�Rl�w�{oҿ�^B��q���G�����D�ܡ���n���u���vS
�ܕ��T=b�d�����2�,2^� �S��	0��@L���Z�6�*�/��tЬ�i��L���Qgi��f��`�����˾���0|Lf�Xl�uJl�X��7�:rs_�z8�&�|a�%�3�Ɗ �P��]Ӛ���;u�X�Ծ�d� ��;66׋(7Eϴ��b�����R�T�Ѷ7w�Fm�{�����n�|�`ٟY���aX�4]~��lv>`�B�7"�9��Sҷv[LU�N�<^j�r����wMn�F�cEm�:���B��Ac(_���n�����l����.!zC1_��a9���~��c�����ؒ�M9Ie�5WU�R���*)�󩆵�~��)�2u@�S����oR]-t8�kR%��t99&��7+/�U1�|UJ�Mҝ6���8\��7�!��z��5y����uU�|�g,�߹���2����!��x~��j᪻޻�ݱ��a �iU	4�}h~*�%��J�mQ�\�`Y@�f�α���E����y}*��BB花j6��R'���ܪnq_L��9����Z�ɴ�?��@*}
q�~}�GV�U3�]����/�{f��9v�al�tѳ���^R�qLM���v�p��.��,V�-.�ā�����g0�ʾ��c��w[���Ǹ"(�٭H��l5�\&\,��lj�*ƬW$���9Sŵ=!��{FO�jO���Cr�զ7�=v��B���d�����𳴏P#� v�+�md�e���v�l]�����}҃f�(�Icӑ�<��e�����4�����
,NQ^1����[34Ь�p����i �;��*oE�߼�o�*jV�~���ѐr����<Ő o)��k��}��L(}�@�n�h�yd�x��eB��!���S��I֗R#��O��O�p
g��So����s4'����Є����F�x�*�~�`��G*���.[��?q7�ى��t��h�lm���I���t�T$u��`^�Z�Z.,�|B�}k����$���p�������g�r��5@�msZc�L�Z�س4/��W����bD��f������`�)7�ps����.?�.�*���Gw�C�M���@)/K@)�4\R�ɺ'=���'<z��]��Q$���cȟ=��)�<
_��(��]7S�^>�k���$C�&0�"��V�彅N���2uGe1�~�����~�ƿ�9b<8�G��!����a�7F^�@��퓻h�̪�#]������� �S�)4�l��!�7����ޘe�j��̴K�xё�6?tK9�\��o����]߷�r@j��s�Z�!-�HHZLS
_+�U��UPjK�!��yr�A��}������SC]��Bk�[�-墟�p'_�J ,�;�{*����j�ϝ��ո{���h�g��1��S�G�9�D�~�����Gi����,x�k#zÆeǋ�|�Ǌ�w�)���Ǝ:ڐV�0`�JL_��H����k��?*��*�a)���
ۣ�+Uׇ�u�iX�!`�U��Ϯ�,l������Ks�{�V�&���oҋ!��vr��i=zE��M}����y �;�&U���N���2SeT��o�?R�$>ڸ�*�+�~ػ#$#����G'Ǔ�+�R���$X�������l�@/0Y�X;�\����4��_����.s�B��-��Wو2�?��RG6ɬ��K &@�����8�`���׍ ��pQ{5��u��\�xaň��pjj�n9d�ݮ���2����i��C�@Ð�+?�VՀ�Vyۣ�}䃳�u��8ڦ�oZ��o�<X���8�:���D��aF=3fѣ3�ch��R��I>o݌.�9�2���uq�a�44Y������ix��?�&m5O�;>��9!�A�7ԑ������ yzh���t� �xmɹ$
���PQZ�C�/6y�0�C�n��2�h� ���\��t�*G:a�.�4����^��IeO�}݋��y�%���g�4X!>�27����(i^՟�Z�zʯ�&?��z}�K����!4үpu����կ�����'�or�~�E������c�kfd(�A�ҕ<2!���HU�؅����w�3n�+�� ��;�;�n��n��m]O=C��k&��s��_�C]pOo���J�6���O�5ܺT'o8��3�#�!�T���qB�P�u		��#����7'ܑt��>�6��("�B]�&�K�������N���V�,����DFPo5�iŎ�q6�$:o���Z\��|�ȗ��E�vγ�@Mo \��k �$��n�F���0�w|�=��
�P���y�K�5�{R�>x�����D��������$���e�u'��ui9%~=�����@!l=�ޖu6=	E��*a��[�;`��!ˤ>��
K&ޚu��Щ���Ct��Ֆp����sj
8�h}7�!��V!�n���#��/r(��&㾿� 7Dz@Cu盞�b���Z�#�uhԼoW6���/� �&MiG��a��iJ�"��J��]�%�9Ƅ��р�ꆕB���*I� ���n��,��Ԍ(��)b�0��3�e+�$6��ꪡ3F��Oe�@Y(~����.�Τ�4��G�����d�f�p��i�0t盶|��n�=�luq�I��#��|E3د�6-���q6�׭�R�B�Z�¿0�G��n�+07x�Ϛ�)�Q�>#�&�Wŧ��
���m0>^h�v��z�����jn]6�.G}%"z��tH)=���uW���3Gr��W����}�)P_���پO�<��Zj(*%�����~%��q��f�T��Պ��K6�D�V���T:�F�O_��~�N�/2xcw�I��N@�E�*����}�ϛ��Θ��1[��(��̥@�?�nʑ!�j�3e�Pŗ�6���1M�D�s>*Y׿S��Ќ˸ǝsBnk�d{���gi�Y�1�������m[}�8i�v��ֹ{�p�^=F����\��AS�1o���4|������(M�*��ɧ��K)���N��b�d��!��ݔ�m0���*$v0�y������k�u/�h+���_�����]���ܗXWS�/Vy�K�,�`����>����q���ok�?q��5��XN;��7�hO�T���ؘ�5^c����ƽ���>&��+DIcΐg~u�Yӊ��)F��o�)�;���ߋf@�BK]� �&����˟I��Du����޹�������x-��.�Gkw�1��[�5?�Kգ�p1Y�"��V�΁�=I2꟡!r�
� `��[�(-oy�f�{����fߘ����0����j��AUkY�D���7;JH�<�?ǬH�R.x����g��o��t�8/x�C�= \#}O�wٍݹ��tǞ[�-���e��U$$�>�-�P��_L�Ú9�U�I~�����-�0#���jz�d����BJ亮��.Wj��:ϸi�ME��?D�M�N��^\m�����
qE��anR�q�Ck���Q�S����R�Hor4�C��&�[����~�hIq���
��]��Jo�/:|�߯׽��!��Y��>��OFUC�.V$~G7l�ձ��Ա[n�Y0���8����'e�I�TvS�M����/��w�]u�����Lfm��&7��%�mZ����L�!��焂�`-��Z�q�BKǣ젦��7�������;��I$fccs�&6s�&�QDr����G_f�f�;מ���@����Ws_������ø���[m ��v
�i��.2�:�e�T�q�b^�ͻ��3������� ����)wMW?ޡ!��鷼�/	"U����H0�e:*���u�T=�yP���d9&��!�C���:vKe�qJ��,�o(5x\���?%��] ���X4�\�`�mh��<�ջx�L[��g�[e�T�N��ko}��s�9�{2��t櫋��W��U����(��]���$V��٫x���]��s�����.44�hx@�E��ӕ��- ���X���4^
7���Jj~�?)9Y��Aܤ�}�K�`N=������Y]��*'� T�z珕�����U�CHd�d�߲���1��{#�M�7�(ޛ.u��<Ѿ%�6NRJ~w6^��s�Ln�1���7���G��?�������=���ƺ�/���2L�FԚ�n)= �m����Ȑ��&yU�d�[�:rt>�f��ԛ�@��i� �����;���Y�@�da�י���z� ��]��"�_���|V��C�06�yV��dg+��������'SEw�Ȏ��/������u��@�B�7IƌL�Og�;!Y������;�ԁ�ຎ o��7r�!=�=!pg�Ů:A�z��$������z�:�FJ}Kj�&! �0Wz����TX����Q�w�D*�u���!��Zuri8�!���P!�O��w<ˮ.2��(	�q�l?
.��/D1T�<�D�}QV-i���.ى$��^��Ǧ�T�Z���Z.̯��@����tN�U��ė�5N�}�>믢v�t��AtFϱj��/3���%O�b��1�����29�6�|�M�/��\�.��:�=��9�4��sPNiE��s�☉P��.~?��zg�==�y�׬���co��( Z}�Ch��F��t\�w�~���]V;u�����=!͓�<c��ŀ/��3*+` ������ю��Iz�]�r��M������u���(�e�3W�J,P2�pNq�MkȽc�2�v򺑝nZ�k�wA�Ԉj���,>���5���87��Cr\u��3���ORU�a�O3�3�U�qBqS���8��G�KԽ��[m|�̏�I����[䈃�� 
IR�e%�I[~<�H���~m�DU��:)�y.G�SY��]�<�ae��W������=:��G+>���.@C������6�����,���bN�[M*Gi���3��NV1���_��M�|�Ͳ3V{�W��ah��`��=��t�vz��"��m�&�.XX�ڟ>Q;���~2|�{�sc���kV�xEN���ߌ8�:�1+�}��<�����x���2��"�g��"?>+�u�����[��D<U�j�����TO�������}���#(n�{�S�l��A՝>����ۉ}���3}?�'Ӟ���l�����+�J��aL:
B���r�����=;��,h2���%|��4c�!#�$4�b��;�S�Qb������R$ݾ-���FX��Ƭ�s��#~@h�j*ղ�c�]g5y�F����N`a�����qq�w��>���G��y$�E�WVT��2o��5���z��<�[��C��� 
_�}R{
��̆�}ڍ	�b���D�|)>�k���=���X{��Y �3������P�A	_ś(>.v*<[��5&��v��i{���-_�|������S�Zh�������H�WfV�E��]�9����fC24�,��MG�s����U|�B�3fڿ�r���(�̇������G��OX��ή9/�Pi�!�mL��d�D������ŭ���Λ�=5�ytذl(�����q6�r����>�v���W�i�Gt��3�ٰ�ʺ	�Ńb��9���iJ����o�6��>Q&�2�#��z�6��4@�0��}(/�����_7?���з,m����o����'��p�|���iU�\�w���@%.�'�#�sf���.W����e�f���@�:.Zd��=J3V����y_�CC���m�[����9?�ϱ��t}+E�%��ۭ�'�8�㇄q�O�t����I���~7�]�,��$���PsO��MO9��E��#p��e5:O�#4j���z?$F�u7�����v���Q>&��{5��ݹfEߛ�5�J�-�;�ص�"]k����Yd�_�N��$�=�JH�Tp.�=�_���S'�'a�?_����T�,Uz���\Q;��g���`:TW��c�������kV��?߱�`%��Qb�:O��(`o�%�V��F���#������\<�ڮ�Bt��R:��8$����@�q�D �ف(p���Lus
N<��
��i��B���]k�P����}�Ni��M��!�RZ��j�⿧NL��טI:�63�lJ�����fL��'�h�p��~�E�>Hx�O{y��q�IO>��pE���>��,z�����0h_~�`v|"/Ò(�_I��	���qD.v0��y'%��@��.�	�iw)�U`��~��fQ�ݠ+Jح�U8�r"��i׌��I�!��P�1��ڷ�]�^!�bu���_ZV�"^�V5�\�5�]��[;�}tbX�����s�i�e,�\�7�������^h"������Ѩ!4Y֞��Y�3{7ӒC�_�Y#�uCd8��)l�cl/�wRm��p��G�}�\r(���@��r6V�:.ճ֑�X�`>fA��c�i7� Ӭ7R}�1n���b�9�U�V�q%�M�iY��/X򊭙E0���^�/.ֳw�^����<��>m�wr��Y�F�(Ge֬��q�'[��E��^z�R�w��|�ϝ[����t�jo��j���x@!�G� =��fڴË��{�5������Ê��G��l|U�Wus�ښ��!)e��T;��GX�d	a��ڮ9������9rg�P�1�6�dc�]ȕm�&or������]O�^;�p�6{��ߝ*���Kp�fZZ��b��<���D��v�M/���f�x1�x8��12��}5q��7�>��/,�/cr
5V������a�B��?<Z�G�h��z7���s��K��,�����"��Qg9G��c)'��,]�`�oۆ]���zY���,,MN^�K�n|�1g3h1�}t���e�M��҄��u,f����C�ˤ�����Ɉ��^Xp����j�Y�IK��;�V����Uޢ�`y���'�@�?K�m���9ks#����4�U���C�3����XV�B6��<e(&�x�[�G��c�k-����'��'���JEXT�?mx�]���|
��(>�W3�="NF����Zi��lnK	�	0�5�}p����G'�n�%��T^귅V���*ϡ��?m�괈�|�>0_җ���q�ƦV�{��u���z�CA�qc���#�A�\�߄x����o>��'Y �]��Z��3bw����IpGa����-d5e�o�Db�
���6�ԻZ;x����{9���ޖ�&7Ŭ�XDQo"Ӭrmܕ~�������}H: ݺ�N?���\ώQ-Xu�-�0��Dᘻz�V���G����9r���M�}�������pQ7((u @�fQ��qu�M F���(��l=6�ţ���2l����n�v�P���;��oP.n��L�5���=����ۘ��:n�nM�%-����^~������B�����r��z��h�}Nʡ)�\���J2�ܥf�%T_f��"��fܶ��N!���;�9AH�)�ز�,�Ah	'����q�2\����������sȁJy�� ?uݎK��i�
]K��hsyh��8�'�u�,]�SU[� PyNC�.�ʍO�TT#[��~�0
d���f�m��5uC	t��L���V�Q-�%�k���;�+_��D���
�sn�2EvV�f���!*�1���}FH���鏴j>u#� ���i������4��B\B;�<��8l��M��!]������S�<,%��-���J�	W��f'*�)\�G�/5��BR)�u������ְ���Z�{z�xu�-������y���� ^�ڻ����<nIś�ӈyMޗ#n6ns��iP�4BKR��	ɢ<q+����)$���`��Z��W�#��o��;����&^o$��su�,�7�?wm^����'�]�|�"h �F�0���巴{*����0�,�� �lzW�ts�d��U}�f��ɵ[p9�ڝ�W�T���R�I�Z9��p�v�;J�4Fa��7(J�r-@�킦v����yQ��̭��i�^F�j�!��G]���Sǥ--���pt=��Q�@!^��Xocsx��"V�Z���Z߶�}l��_����c����ռ+t���]���*5�z�~����,��>X��(�Bt�p����0 ,Y����j����!x�*~�/��������g�S�����m	ŏ;�Cł�] X�u.BQТ~����^�8���F��ӻѺ !׾huϢ��|YS��b��&sK��V3�[��y�m���m���2��s��䔋�B\"���\�w*?/'�>���%��NF�):<�#�7g�&e~H.��� �1f��^D�'5���I+��V�[]!7/ǵ�؎�pUj�G�I̠�*��:+���kk����爵��3����`l�@��e�|�B�2ItT_*wKnf9�j��l��&�֘��^Z�O�TDd:�R�����f��˼�|�J�@\|���wl61����}C��v�4F�J���p�E�9���	a^�yq���k�O������7K���j�˱9�3��zp�o�O	���J���|Q��M*���>-�{kĊ�ǘ�H��=�����6�O�GWHbu�ρ6K��}ar�6)�u��"���c��?WI�AE����索ŏ�v���`��XL�،O��ej7�译��/��5h>�`4�I���(�u�,�⨻���q�Jfd��x���jTc�О��}-:�o?n-�c�qf�ϸ�0z���git��]y𨺠����}����@�4K-4�*i���X~�f@5�m��_A�m�����ǘ�<���v@�S����7.���&`��i
��m�h�|�ߋ�|�:��g�9���(V�ȷYT��G��3q\�9n��B���q0����<�h���d�K
�������~���.`9#�)�yq5C��;�p�e��f��BAQ�~�����{�ޥȂcN��/4f��:�03_Ut��|�?����H�>d�@R�g萬�Ʉ-!8:����Wi �)p�ku�2V�`'���n���>�B��F$��jO��>W�_�
�ht�#��]�;�����؊���Ҥ��!B��uuʴ��s쵐#��f:UhL���*}cB���w��^aa��Se������}ȅ!_�a��@��M�G�(��F"��Q( ɒ�}�xB����Է������$Yk��Я��*�ߐ���&[es~8~��VT���VG�i�b�9�F�ƞO?/ǌ��R�^$@:j6�l#Q�?� k!�x�=׈��I�2	$�yW~)��hʌp[uTcW��<+�3JI!�������q�Tx���	MT�e�^抾�c>����/�#�D0��,�g_>�){��^���:�9�xD��F"�v�q���v Rs,x@���3I6��͆Wނy�@NA�[�=b;G��R�w��
����b��}����t�o�����.�J�0:y�0/cl̬�o~�*�ds{�+��X�����N��ȫ,����`�f�^
���N/u���{�z+U���)�1��ek:zS��Sk���'lW�sJҸ�RU�l����?�\6�{��V��%nh��f�:��9�����iQߚ#GO]���@K4BP��N�'褕o+���I�|�}5�̭�~�`'yy�������e�j�>�חM�����)�L���C+�yHD�FЃ��yY:ڄ#�bɿY�?!c�ڟ.�Iִ�emH_�������y����sm���G4v7�c���*(�; IE�5G�N-�����T��P.��=I�X�۬��p�l�W۠y����#TMi(�p������	WmY)%�L��>��D���=y9��_�2��! ��M�w���?5(�?�­�n����ND:�A鐐��Mw�H���Jwl:�E�s��}g�}�{��;����5k��/�zg&��#�ݠ�q�M�z_	��Ỽ���j���ӌ�[a��R���K�k��V2����ًޯ�BQة���{<���� �JB1BΗP��i��V�HN�k��S1Э�<)˯���s5�f���Zf�ܣg�A�b�E���
yȰ����mò�NZ�K�W�rBj_f��k��D\�:@#a͖��T������ ������7�YYF�:�)h��%�o|�e!����OV���*r�x5X��<����DɌ|��8�����L�a���9~�4�d =a]�Á��ʰ�B��}��]���ۇ�\k�3%�ݔ���(,Hf��Zm9�,b`��Ê�+|LO�UxMӥ$��=�[ko�u����L�$Aj���<���`�:
��*�����l�['�RLI8�AM�5��Zk	M\]s�����K{�N1�x�bC.�]�p�YDn��T��u�F������vF~Flt���g�|�d�L���Gˆ����B���P�r}�)�[�NH�懒C)��%)]R���L!�vɤ�����@�*��MS	ԉD|k��^#ͨf����a΄}F�1�n�/5��ҩ�gyJs����/*���Q��A�\@O�n'��}�7�1g����62iH�d��'x%�����$�_�3K%���Ґ�Eq2w�]2u��q��W7��&����+�J+��d���	Q]7Is+�lջ�}Tw�
I�Z��+����-��~�E�|�~@�׽�V�E���G�},2�Ȫ�Ԡ�yЉ�$�\���v��w�E?=��󪍏"�
��M�1��O���t�� !hp�5�g�.�i�S�Q�f�A~�����,ƅ�b���|�ݗ�M��ďc@a
���V��EVJ�Q3\��$����g�P�+ʞ�C��uK�fPm>ִ�J�GV��*3��n+*I?S}�D`j�ӕ����p8MSaFX/#ʱ���Z�X�r��cE�`��x��b=����Q�:�B/���0����>��p��SX굡0��&����QQC���t�9��$�+�7������^��![�	�����q���PO]}��y5��AM$�Z񖢗�*����Lη��tisg�H�nEI��y��� KH��p?�XH��M��φQ�J�>���q=��J�
;70��������;+��R���%TH�'��������ݣԫ0�(YocK�]���!v��;���@w��X�0`ԋ����:����u��gL ���`R���r�kD�����z}�(���A�aѷ��C��a~�p3!���1�g�mWM�L����|xJ����@}n:m����+)�����9T3�!_r��y)�L&����IU�,��{��|G~��؍�do�&)��ny��;��ߵح�1��a��%\J�;)���r�ٝD-�8�oĄbn��+��n�<�޴�����MӿZ[T�*�!�̝U�����m|Ȕw������L�B�K��r	ե���WO�.뽛���XC'�+D������|Dx!��5�S�m��>�{%��D։���C?�TDVJ$�/p`Q���oܐ��_�k�"�BeS4=�6߬����'v|څ(~����M���,�M�=������Q�S�٧YY�?�Ѷ�~�%:7�!��4=����,v����h������u��]��q_7����r���9��Td.�+��	%�6rm���\)���{	�b ۘ��U޾�����U�!O�9P+*�v1wm;IAP�۴�s�C,���79��q�Ť~���1�����g�4{d�=�0�d�Ҟx,�Op~GkϚ�}Qp�}�'}=���������TJ*I�42���0�����K�G��4u>�/�Ub���'vE�`�Q���"�֭G�gB�<�M������8���h~� #�W�5���j"`���	4Tw����<�A�d�����/]Ct�Zl�?zKM�,Q��,��^"��qҠC���,�tg��,���7c�ΌM�χ��๽	�K�fc�����$��?H��:��щ�� �vn��vT��>�����f(P�y{S
̉gk�߸��(u#���M?>_�`ֿ����׼]ݻj#����e�M~۸�������8���d��N�2�!�%�n|��X[1�1�B�0t3�I��>�%z�T�?n<0��R�T�u����N�{Ιu>V?R�|��Ob��f�ޗ�����c��e�#�X��R6�hN�H�COvJyR/�!Ov�5k1(����@ߊ>P۳B^��1��D:�.VF�����{����S��9�h����6w�@�,2D܍/"M%��3���?�|��!�(�KT�a��b�T�lX��t]���*�Ύ��������Ej"A`*07��Ι�C@9Vk��f�6�{k����*q*ߡQ�7�V�VK~��}�-LǸ��W�Fy��M:Om�u�Te�s�a���K�Cij��G�o�çɸ�S�-X�/e ���EQUB��st�P+T7Q,aRG�5���YӾ������ő�2�$<���x5P-��Z۬�mSӃ�r~����-���6T��Б�ߏ��.Pg�چ��7#��4�z L�6/|b�d�&p4�$�u$����3Y�͖3��ZB��mf�fO�7�Ē7"dL�GRjH-iG�Zs1�y���g����� ��	ex[����ȷ5#�S�W���%�'�J��:JV��PD��~�	V�Nb�U��	_2t�+�z���~��/��"�i�q�Ҷ��x�Q��h�����3Q@@�}r~QE�"O��0c�r�N�v��B9<��/��,r4.���j����{f��|��-�}��F|�E]]�{��8�x�0?~��$�>�_�I��/�� K��C���{��Q"�W�����p>>rpu�B\���p�_�6)�����`�z��0)�-����,�a~L/��g�{\�&`m��A��3r(���N�wl8����|.�IB:��]���x���~�GFRJ~.�jثP��٘��]��;#ÈN��Dd�@Z4:ّ5���r�H<[����N�e�>]�ΏHy����~S��t�}ez[a{���w�p7�X�5�u����ԟ�V��@�Pq'M 4w!\�F��8dp� h䶧H�¥�ޮ�;�jO.�D�$�^�F�(h�mt(��7M������85*��
bXۃ�j�����~A�L}{�2�@o	l��Lm�w@���4/�Ն� TQN��7�޸�� �j��+��g�v������p�H��vW����G�?<��0]�[h`�)��X4��:�U�bc��=������h�'\VtHF�17YS��
}� m2�����8|�Xlը�%�m� ���]���}�̦�(oz�fb�q��}K�"�"7<���	uaYQ�C.��WwnΥDjG[�B��.�vg�]!�	U6�>}M��Z g�Y���Q�F�Vb�*%]�F�!X9�!���&�.{�����t�y�����v_8�g}%P��eб��1�d�{�~�U��]b0�����_v�G�{� �0�Y��`�x��uH,�"܃���HQ3V�|�`�K͎�k@;��y���B�^��K��F�8�V�/~�p�ᅏ�"��H��/���}���)��e4#CTQ�׶��^ނ����j�D�d@�4f�$�a�1�H�*���Kբ.3C�n��92��§�L�A�.�>�3��@�Te����S�.��sT}�2O��N�,�X��#�m�]�SV�JkFR�"Y��-y���t�N ������%^� qS��c�5�e߾�&nȨQ�HG��~�bAb[��s�O�6g~B3y�W�����:��I9���?X3p8A�wFN�P8���A�L�9=�`#�I<gʄ��a�>���ݓ��J��0����+Q^��]0���LV�Ֆ�I0�����x�֧����/;5��!���{�2}�ޠF�\�m����I�Y/�Kaww_���7z4f�MbI�ϒ��/�]����09��OA��>"3S��}�>Ԍ�ᑣ0��Q�2����0��6�A;Ig�N8�?N�VA�=E�Ê�����].u����	;�����9-��wj�x�X�?x�8Z�&M�D�J��Δl
R�=0��X�"�}�ʫ ���d�JqY����)p�W����٥�{;Ԡ��Q}T�����H������t��~.5��_�0Ѧ�|��FK��y:����b��x���k9��h\R��*	�p<N��:##�
$�K�JI�W�I��o_���~B�%:�=����u���䭚c��~���`f��6ܯB��x�z|�������T8�cŗ@!��qmK�D�c)Ƴ��H";e������4��%�}`4�壳�o35�C���Sf�D��f�vp��h�d��=ktA��?a���/����"5�^-L��j{g�c߽/X������C0�4��8��G�TDav2�>�H!���W�FN�l2~�c��mT�P�z�BB�d7���K;���9�^�����W���b��H'>U��p�VJ�1v�K��{9l� W����I�%�XܼxI��l���Ҝ�w���ߜ'���v$%N�|���g/�?�h�a����i�yY���$�v0"�R����a��c���[�e�UӣE�ñ�R#����a�j���5�g!���G�6�%� 6��73�I��'6��ι��i���_�;FKG�\�� xB��DA��dࣉ�!��J��,�Ԝ&n����.OT3V�,����ٽ9*�+7���0\�%��9�{/�����'�o
=�{4�_/����}��<�	�O���Ϗ�ǌI�n��Ӯqc���^$h��6���!��:�h�d��Gk�5�"��S�;x���X�O����������Vt]�{s;/A���H���SJ�b��mK\l����ko���JOԪfL�
��nd_q),�<=�78��:�c���<��?<��Q9R�G@'�lC�$k�/���N�B.ڈ"�X�D��" W��]���n�.�c�p�9� A�Gt�HU\X�V��_�rLR�m����\�`�wk^^��_�c����{���&w��`X�;D�E�O_��?��U��U�WO���{�����1�5sR�9ޑ��n���L�ʿ'�����7@l�%�z/c��?�X��ټ��
o����A�(��Y&|�T�[3�/��0�~_5�;vHr�_�( `�l"��%�)^�K�Y���}�,�3ͨӭZ��ռr�����u��>��&Tq��*�p�� :���u��Ι���B98ŏHR�.ϣ:�2-�h��a�om�Ӝ�;�$���Q����E�l�ST�X�}B����y5���!�	w�(c<8�$|5OjNP�������px��E���>g�0{l���Ef���c?�[�ֽ]܉��y^�Ҽ�ˠL�*���4�3�p�C���([�v�2+Z4Nl��Y7!�7�5o%	>5s������A�~T��U��N��S=d���A6^<jÃV�
Uܤ̬=�XY�Bmm��cN	�ݓ�f���1��h�����{���%W��[���x�	��YB)3�����s�{��ӻ��n-�9Ss%�!�*�<����FF��8�?g�vg��8=j��v�w�\��������ƖH/,F�
�O��C�k-�P)���Nu���f!��c�m�O���xT�{7ڼG��
�c��77ݴ;:IS��k���2�r��m��5b�u��0�����������N]��(Tӳt�~��/_�?T;�8ncF; �v�%U����:�帨����q�y���#��J�&��DʙR&\�~\S��b:��$�~��� ��pU��R��m�:Z�LLصs�����;����qO�
�_���sm���6��|4�
�0��W��f:� �G��Ѐ$����X*����Dю�h-���툜r� �u���x�D&+�c���J�6���?A�`���x}�Y-�s����F��S��E��)5�ա,��\r	m��dA��V��ŉ��m����ˌX�M�X^����=/�n�iM���gX��Tt����K�pk�vf)9�|0�iZV�p��8,t�V#�rkܵT8G�G��T'���&�(F]��O6�>>���$n��Y�c�m� �4�c�W0�|��SP�Y�t2�?��4L�ޱ�������uW����|��Q����X/R<N7c��u�醶j����>ʡB���M���'���m-�4�V<�+�}�!��m|z��0:M-(z	3����n�9�bLO\N���?8�/K���.oU��e�Y�0���^`�f��3��V9%�_rk�Η��aI��z��[� �%�n7)����;ӳ���7��a�]��kIf��1�إڝb��ϦR��gr'�;��,���ݲb7�+pP)�'�y>�^�03JAU�f��S����p�Q�d��:V��o��~���c����V]��2L�F������9f�M���zp)�{FƉ��D�EI��a��ә�5��rM�EK�r���Qx��JD�#�+xA�N"e=�6�J�]&�,�#����߀��a�Ԗ�DM9P���j |�`v�Z6���N���k�Å�bE'\�W� 0>8/Zβc,uE�:'�&�G����5�����]��|Bz2dQ6��>�����\%{���1��ݓ������+ I��
O��C��z6`�N%н4��L\�m0���"CZ����Lx*i)�Tx]�z�6���[�="��j��a�0��� ;�7��䅤�g��AƙH��qYf���C��$������*'{Be�%"㰊PX���V+K.�Ԉ��@�ۈl��輓�=*k�K;Z�#8�y����%Ε��4�+f}�, G�|0�=�趍��4��yY��f;K��4�k�� g~fU,�����/!��zQ�z�8BK:��F��	 ������|�$y��-��j�E? 1ɦ�^V�Z�������9���
a��e�:����F�sC���[���K��s�L+���B�ɹ�N40wnvT����ܱ9��6�����/d�7�`MC-F�ͅ�N�$%��n�+�WvU�S
�M�g��~�4(��b���
�k��(5.�|��� �����JF�Ä*�t
9�V���z�1⋢�3J��J�f�t�� ��a�R�!x�	�O2�'�-���J��~�. 
Ք��f\$�Z�W���� ��F����A:�=d����6vU��_7�3;�f壝mt�;.� 
�R���]K3o�9W"��Ԭڄ�~��I�Ս,�M�R�:�([�6E�H�b�S��89=�t��Pez���m�,�w�-�� ��\^��lG�WCY���a��M�b�I<T7�k_��5tp_�.4%�8''������"X��cSc��e��n{%��?�l��n͹~���a%Y��N5��I��LG��\�J����96l�j�ӎ�|�=��͹|��N�rf<�7��",l~$��"%Y�b��~w[����u"� t{�0�����-�LR}bP׳d�"��M�� }�8u�=��/@?�Jq��]������N6X9^���yx���r\���|��y�EOL�q�.
�T�Ͽ�Ϋ|�ڎJqF,
5��oK��;�C���m�&"?ة#�t�p�6	O&�b������N}�)|�B�Dʽ�ޘ������8e�<g#h!�C`g嚫&@��2��� ��'���/C�5wu��٧CW�m-$�q�".�\¼�Ԏ`�_��ף�{7˨�@�bu���_W9
��uŒ���˾JT�3� �j�p�����}J�
�o> e68��k���#i�6f����+����Wg�CM琏���q�Cڭ����V�ھc�H���na�Zϒ$��n3��:D@��N@���_���6�5�r��b`Ԫ'�mO3C�͖R������yz��Ȣ�oZ4��'�:�斌�L@����o(��E���.=���͔�G��(�賟$9�	c}��*&��<���,�M)��U2��X�.�Cj�0����#%/�]��^0{vmo ��# ?�,��bw���yz��RO��̬ܧ���w�oL��a�c��2؊���TWu��8c2��]�Ҁ���FT1�=�~e�j���z��N��	���6�$�	6����jz�[��)<�t��ʹ��9�˿����z���𿵤{y�o���2g�_�2�o�]k|MǙ^��c� >eQk�m5��4x3�ESV?V��h��r&��)-�݉;-����hBI &΍���w����,�`x�Ю�>�!ʹt�[�����l�z�(�����cNo+I���rZ��"5�r�15���dYI>��������(L�|q���vB��I):KJ�Go[�����xh���P[Ӥy�pչ�����7�{�k]�J9K1
��2LQO��r� U�vN��k�k¬r`���v�_2
�o#J���@��F��Bo-� ]�!=�&��9��|��H�ł�$�-��Ձ=숰��O�L}��0�V�fV�a���4z~��7d\�������;��f�D6"�TV�A�VW3l ��@G�Z�$\2I���]�X�$h#ԙ�b���dA6܎�QH�8�?��6l�;��z�}⥗3��������U0�����r��9��0�=��jܸ� o�c(�I=(�Z��t
��I��R�����(b��m(h�&�ɛ=e������kږ����`9g��qە�]gG�J�4�)������K�v���dS�w貙���n?���7,�_<�-���^1/��R��לK��;�u錃���#Ԁ?������W�h)����5 ?�o���)��z�ׂ��th��u�F�j��̻������5\喉w��`��%�o	x��)��� 	o��TK.S)��_�7{�`L- 1U�6CWnO�Z�����OΟ ���7�ä�W��ًYi[����q���%���I��y�/(��%X"GB����k1�?`t�=���:n^�\kZ u|�̼+�����u�G��=��G�sX�6n��d�(�cN��G���,i�4�����:	�P3na'�������|�g .�~�hx��+�oDG��">��J���7�8,�[�
��>W_y.�}Ԅ���:�� <%PEe�xoZU婽^*ɫh�`�����8���4�/ɿw]8�;�.2�UY�P��r��/���&V�T`&U"z8hذ�s6,��+�i0~lTO?>ۮ��${�ͬP��H}�ԍ}���l�X>;ߩ��܉���y�w|iKi����'=n��)��M�0x��w�6:�֓�7{	�������	��� E;m�l�Y����� ����M�8S�8���6��M_��>��w�*�����]�ƕC���~�V����t]�#� A�g%*,A��z��C�e�Vfc*��VZ�{�w�g�A\U���O6��Y�;7y�Tы.hm��n������N_�|�\!!��o@e��d�Q���P-�:���V���;S���n�c�����2��jp��Q���$يU��O�WE���/��G��X���=�l>�è��ѷ�`ġ�mA�G.�H�}]�R�6�u�����htE�uN3fǢWcJ�;*{j��*��6���Cg�#�p���?\���P���?���rq�돫�ރK{��Y�92@�/��9��,��csW�V��_��e�!��C{�pP��b�o�x�e�}y��X�?��0`���t�n0���Tڨ�X���U�,�y`L��N� g���I﬛��qQ���d
B��˻��`�R}�s/�5�8rzvU��N���5��M*�Y�N�Pn®�'��vN1:�RI4��K�;X���Z�Y���1�iQo��T�����)#�w>N�Ո�jsX&��v��6>�4��t���f-���^D��黧a���̳�|�~M�CI�n�j�*	C��7����Z����'�S=.���2z���o�:M1p̸�@��1����q?�'�#褬���1��i1"�3�R�X٥� �s�f�������W��赗�GvןP3��F�\�*��\���JJ�*���bbd*�Z>斒e�()�,w#�
���K�K�|3�+�!`���4ܙ�̰�����0��&.�p�*Z�����k���2��_�O��Kh��%4��PB���kл��WDb���s6�|(?nlOzm/���kG�t���j��Jh���`��Wn� �"{�����C���#� ����Tz�>���-������[���z{"�t�R�rF�̀�h���5U�Ky(8Lyd>�gl�O�X���(���q�_�;f�Ty�>Tw+L�4�[u���Qũ=�d��}iW�m-�,���*��B��ùW%�!Z��F��Ԁ�(�51v�m�4�������J<"�uc18�.�Ŧ��c&u-���`t��[6��b�S�G���q�*��ࣝ����Gz�	v��-���-kz��c�寧�\ 1�t���a�{^���lB�@ɗr[�b��~�}��}8��6w��e��	�fzbm��h�� SŒ��@+#_��,r�'t,�����H2�ܓ���[�h�J�x`a�����+��6c�I+�n���Q���gO�2���5q��8֎RL-���
x��KU�ыr�����Y!Zơ��س��mmY �x���@�a��B$�)_C����T�4��fcR<:�-ӷ_�BM�p�Y��_�7 J�H�h�����-�b�7	�
H�[��B�Ϝ�Ư���%g5���̙�{��0�;��wU�7�[�n�ە�JZ1/�\M)'sShu͔�#}�`��}�7��/��K�,��!�.���O'�E�b�NJ�x�N3�XL��e��ZY���{%ֹ�Bsl��v&���fO�?���%��3(I��-��\�9���F-��6���o���v�	�~�;(�L=��I�"��I�aG���堝���q�+�bg��W�l_��͈���lQ�qPsȆ�ֻe�%7�w�>��D���R�&@�V;��Rut$*:���`�*����I]��ٝ��
�s���:t�䪙Pٿ�R��8.��qgV��v!����l�ґ���޺�_�Liĝã�s�U0��ӹ�A�%3�%��d��XP��S�����T�����M_}B=�����b�^MaI��D�gk��c�`�~]��a�&O��%�e�"T5n�Mx����<�>����Faa�T|}z��-.D`B/̘�6�JA*�}z��*�b�:�&�_'����R��_lT �������r��\������e|�~����m�3-���4}Y����0®��Kݣ&�_u~\��A[2
)\o�BJ�O����;V4����n~�;.���8,��(���L��Z�.���+X��b�U���R�?#e?a�5dڐZTK�>$4#�*덼��>y-K+��s���*��[s�Zƕ�@D�d���)��������yGP�uM�Y+vQ�\߭_	�/*��X�J�0�B�7�΁Q7I	�U�/��3	0��rpԟ�*ND[4"�4
��-6R�i�VY�+f���g��Fc��+$���c�H�����j����`(����ţm]�9��_�������kug�p��Q��v<I,���T6�R�OM�����bb�#�[~>��Gs��Y��O�FZp9%��Jc28k�-;o#���3���t݈+�/5�5��6��Z�D�v��<u���.��Q���+b$&x���v՗:"O�j'wBx���ęͭ����Tұjl�	��ڴ�$*���V~QUw��܍M�βl��^WC���)�GuZ�^�v��[멺�	�]��@%���T`m�B�KD�X8����s���{���[��q�+g����w��|��f�Q*{
i^2�"p;��s~4�}�i�z�p-SAO����bA
A.Yc�8��ӫ��U�X�ZEx����+���Yt]�\�ɛfj��k����.�6cw�5���R�gZ�!�@�J<§�J<�D��Yv'�:���W�M�R�o���_.¾e3)���Y�fY�̉
q%�uu��C�o�n�v�Lb��l�Tĝ���ZR��H��ⷯ,>� Z����TK�9�*�@�^��B*�]?���J@?)���b��T�|%�,䆣q���i�����}���,pG����X����ÈZg8�!���l^�C�X%D�?.�����'�����!�uΒNꩅ���ө2��u/���7s����Q��K����N�^��Y�\��3���8�#���ܐsz�'�}��a�Ь�@�i5��1S�P���*����#�6-5��m��^?�9�o=�;�
����`}�aE/<����*����]���7#6Ϥ�e�=~J���۞����[��n#@�������� �������N��P��ʔ��������৳�q�x��oj/]�?����������p�:yp�IG�+���5G��*���q��RP�QhsD'~�r�.�1s4ln7�JR`�}�F���-�^q��[T/-Ƙ���:'��2��Nr��@x�4{z�D��N=G��j+��p?���6�U{�v��m{ih4<~�U�^���\��(��(���jl��gG.=�=F�e)��r����)�ń�k�3A�W��aΈH@�B1���f��lN��B����A欠�g��/֍7_{rs�Hz�9��eo���������.�b�W��XM�����I�	K0�"���m
N26����BjZU�J��o�t����/�o��Y��9����Lx��p�{�*N���U���F6�]�.>��!���~7s$_�"�>9�w�V����$WvS�?�y�{���T&fbä����jγ��}q�*�Æ%�Ո�^����K�&#�h߆��dܿO��O�an�?�g�<B[���s�L�pM
w1�H��v�h�@+]V4�h^ʈ��H=t���dL�.M�j��ў�����zzr� ��[��vAшob `��)7�`F)H� ӕ~��Xػ2eOxϗ�iA�z���|Ǎ����=�F��c��.f�f�䍳 ����B��&�%dR�:�`E��o��83R*:[�o_��p��-�BW�?v�*ډ���?�Ϝ�� �6WE^����R��ȑze����5����P�SN<�5��v�~��7hȷ������	'�~
/��Z��I�y�0 d��[�&B��� }�,��e �sB�K��-C�^�)$|���x�o��/�_��eV>�7盷��o��ݥ�R�Q�h'&�=�1�f>E��3ߍ_�ъ�zX�r{�|IAJJ��p�n��8�;1�a�z�d��[�a���Ubb��'�(lc��j!��?�^�*$�hmΏ�	u`B!�,aQ�H�^nl���k�/�R�1�������6���/v��r��Wv�w�J�DY�{aĻ�Y��>OTo���J��� �t=ʴ�����9��*(f4N� ы���'-�"���2�uR� f�:�H�j�ʾl�bw��w��%5�n�]$G�� �����p���o-{�AM�o'�-sC�7�&��w�[@�%]��t��&���W$��j���@h�^�V��~-G���3�gy&W�o��ؠnĶ"��7����0<�ݿJ�;�=& Z�o���|��GF��N�f���O��k��OY��e��ښ���6؇\�s�����t��i���N���&�j��,py&Ψ���a.vr��-ZJY��I<J.�ѲvT���K�E���%�F���-"�0�^˪�9k��l�g�~��:_ӂ�Y���h���h�O�
'�-��Xs�����}����]
���
l@���^S>	B�;����e|�˛*�}���nF�g�TƨB���o����O�̄�r(qN��r<��$&K��yy�(K��e�[	�\� ����Y�B%��v��t�:���R�h�]��3����>�iw����wSl��&YƻK���Op�i�5u���b����o���dܪ�aFF��PD��j�	=q\\\���2S�(|h2H
�d����}��i"[�#�	k����F�{v��)�m��>}३�B���ݴk�I�͍���2�|���?�yK�����z�"Zs%��tg��!k�s%s�A$��܂54'������eM)�p�씩�J�H�$�ѷ#8�@��u�Vqq������N+�x���:3l�B�W��֦xO�׸QhוI��M�d܌���<L����ޠ'&ER�PD�c��o^�S���A�NT	R�T�@^��^���ԇ����p,L�۳Q/�i�}U���gM=Fb����V����i�������3��)�5��q}��;k^
 �E��Z����!��X�6�Ɛ���^�u-EZr����qS��r��^'U_{�������9Wr���Kv��f��I������y����I��O{g�	O�-S	ey�q��T'�^
8X�H㤔�����U�|]G&F�K��¾�ƣ(]�0*K�o��.vMzM�z/z�����V�w��c��?���\P�XxA�U��h���"Z�������>�-)�fu��%xxs_�R4��EE(�֔�8'�h��(�X�[�	����	 ��n���Դ�OI��O����	�3e�x;q	����&���b��]�cJc@m�H`lu�7J�Gf�2v���U�A#����&]zO�Z�&瓛���,�头
ǋt<�e�m4ژ�~=�j���c\q	�zA)�Y���k��YN&���sO��=���������	�Z���[�o=C�r�������wT���S�P�#��k�r"R�����b��x�J��u4"�=����x\�������E��kXLa���h���m"����=�ן�Ҷ�*|�pd}�+zl�t��`'^���G�k���6�@����ͯy8�9��>�2��&W'`��7���H��VI�U���(���ՙn�y��I
cj��&l��q_�S\`Ų_�J��}�0��K��1b��B��])��}�l/�3��D`���S��v��Qd�Q7�H���Vnd��� ���h�_�Kt@#�=��ߣDŪ�.����G��V�Ć/@��X�g�9E?�,LX������L���[)%�b������gnl��t��;a(�����p)E�ޗ�*�2-.ٺ����pV����F�}vg=�����['�k.�����L8�{�/���{.�g̶�?���*y>���TZ��$|��v{�����Lu%h7BjׂL�Ɵ��Me�t�I��h7J~K�8�P�1����,�S�t;-f����,%E��ED��jmD�ŷ~���5�wCT�Ѷ��� H]�^ƃ���*�8̓ۢ\�b.��]# @*@«�A~ӥ%O5p��߳Z�'��Œ���[Y?��*�<V�7��ړ�:QXׯ׃fמ��!D��:s�u͇d�w�au�αt� �׆�'�U;�Lw4���X�6
��- ^fr���[S�O�IW�ɕ�(<���*,���'b���H��a�a޽n�j���N��"@� �`�)s�1F9�͙���\T���h)*���w�iO��Oa󑑐0UȞ��Z߁�]�1��mZ��MZ�l(�޳k���Ue��7���~w���pr����F O���ff�d�b1��w�C�����_�`*��{�kt.,�T��q�mO�-طp����x��a���tہ^e���a�Q�EW����k�g�����#�|�=n�9]��|�Ht��%����$�t����j�y�n�����T�z2��`\r�K m��#I�έ/*�+���"������h�8���:��U(��̔0 ��G��k�!��*6�;�7k�({v�'j�s��(&"FԔ����$��Ŝ���{N[=Q������O��W��@� �#�^�Ǔ��;�\O ?j�J��T(�7YS��4����/怸)�v_G��G&�4��>u8+_6��;k��)cG�׶?%Iོ��U~ެv��^d{�Ҭ|u���2��5V��;�Ӈr����ު3 þ:m�|f@�9l?iV=�e�����y8G�D���8�"%Ն8��rc3��g��B�U{�K+̮��L♢�ï<�##������O�"P~;0\�}5�Zj��j(*v���v"`8�NX+z�Se��j���3����E��}|��(�[��z�2��#?��R�_+lb�k��Zu���<���%'#Do�Z��Io���_C��]f��@��7�$ �#���)�D_�N�o�~;+�%��Um
��,�\Ur}����x҂������S_bvB�݂�JJ֎n������ND���[��IrVpP1bG��q'��L���11�@>�޸�t46�VU4x{+�f��H�<�ؿ{(���G��p���+X���G����Ϋ�d���Px�Crn�v�Zh�:��*��Yr:�|���sj�ѫ����s�����fnEl|h�&^�=]���'G�G���q)���Lv��)��U9PA��7��!�`n�Vb@�K������T��ҫ ��eC�l�2�W
2ߒh�$�IB��Z0�Z`"��=cᏈJe��.^m��A�I.�I��Y��Ϡ��e<R[�����J�^&O�q��Ț��S�y��Ml�a�R�\#�~���.7BE ��w����:���7�7�r9�A)r�����.�̸�ݒU����M���������
���������q%��GF�(HH��F�@S�s2��r��$��'EV/ZC;�Y+�q���`��C�5 ��}���nl���ƶmۍm7�m�hl7v��������d2��ͻ�{΃��x�v<�v4��;�����	���'w�E�Ŝ�\�v�X�t��)�`��Qm����I/d́�/�SX���qj���?/�7u"����'u����Ȫ�öRb�ٹ��(j�W�O�E3�p�^)�Z�ߚԆN��W4�U��Ry�U;@�S;��+�ع��S8���L<S����_�s?�U�a�>N�eN�г�x
�0�����U�Vt*��:P���^2�/�����؄��n%*�u���pCb9O��K;�Q�y������yua�܆}���G��@�	��j`P�U#�$Ǔɍ��
�)1j*l�/�y�p�iwC����0Bŝte5��b�$'���/���sFE�?���AbQA_'��Z����!��H�D�Φ�񷢅��C@
��wղ8�7r����ִFW�Յ���c�LpR���H�8O%�VH��2W��)xhΪ��X�aHV���L��#OP]؟��������N(�ަX��+c	1v�F�ڈ^� ������D��@1�d�G4��C��-E�~����.�Qǵjl��ɟ�p�@$��b�
|��]&��9�ܺ9�C�M-��s"x��rU�4T��-p s���h���L�H8�r�����u��P�g������=��������y�����3M��&t�0]]qm�X]Ɔ.c��FTn��ȁ'!q�)V��>ɓ���{2�r a�کU���e-l �;��>�-]%"�×,�g���
���}��W��c���l�1���0`��ɕ��";�S*=P6��;ۿ=����K�& %�W�Ŋ��Z��w߀T�LL��aNH�M�x�����L�^���DT$����`y5�1�y�2ԊL�vE�I]m���]w�� Q|o(y�&�y7@?�+j�Q��O##�+f��)�"�*�,�빜U�gh�E��0��K�6É89�Wleu��A[��<f�Pɔэi�ܧN��5T���d�p,��o� ;1I��A�L(��V�uN�|���N
�E\2	�9�,hM�z�ΣC���M�J�7IZ���Z��n.C�l�W�Z@���P��w�*��n���Cm�lo�+�ŵ�t���A�;�J̯�7	@,�*��Y��P��n�U9:K?&���E .�R��� P=��m�C����f�'�S�8��	",S�1�l�������6�:����~PB�{MMQ#�	�}�;�k�e�>"�t�(H��;�%���>&��UqO�\���)���H�/��
��\n��.*N�t��VО�#���5=2�iNrLD 5�׼� ���աz���݊�����T*���h&Ct���`iy)q���G�j
����py������gC�s��!�#�P����k���D�:�-�C`n�����)�[�)�r����ܳ�K��L�����`
�OM����n�Era �ڦa��0I?��w���^W��;�z�-�f��1d$r�:N>��x��2I��͙1N	�;�.�֣�97�PooĮ�W�NV�?\�K���>@;w��Rx�{��[���
5�����	���#��ډ��9���%��p���]*|5��+9��Rg.T0.Z�Ob����6k;Į� 0�6i��F�@�W�2�'Ck@-�Xl��=�޽m�)H:|&X������[�n_Z��8΋�B@�#Z�x�0)��x!��ڕ}���r�vGm����qD��Ԫ�@K�J*g��o�,�����f���a�!����h��tK:1r��স���M��)d���������j����B�Z�ok�~C�����;���ҵaQ,���
S����6贽>�}>��型ގ���3�,��x�T�u#��@1�݉苔JE�i��o�Q��W*0���Խj��zb�3�/5;��%j{�B�Ϝ-�{1����E��$P�P�hvl`
6"~��:%C}n�T0j)j̢��8���Jj��ĵ�"V���g���{,
xB�Ȇ�N����pŅ,x��K�8o�K������¶[�1�@�Ƿ3{� �qJfK�G~��`EPG��N	8�tBq�;��dt�yW��F��J�5� ��0X�6,��H`u�6�m�Y��
c�,ת���7��LX��t�[����~)&՜�0 ���/���Eɨ%>���6&���<ŇKH�,N�[�b�. �>8[��sً�ԋ���Ѱ��T���4�o��q-���%X\/KfÁ���(�x�"�as`��͒�OD��]Զ�a@�V�ٟ�r�ő��'����f�׹|-ƋOBG
��D� �y�B�֏�����Ԃ�)�1�/���R�|mu��@g���S~}u��z��� ̀eVz�x�i��u��4��O�Bm>$��?�K	����(�Ti�y-���z/��J�Ė^����c�т�B�V|�}��ַ}Ц���xv ��
��F�&t0}�#\]z,��0;�y�X��BCK"nF>Fً�PA!9s_�{�G3���;��w>)Q�&���K�E���Y6���z(��_�0�R�#f�:���=b��a��'OD�J����R�W���8�#��a�P�c�rw:�����6�u�ݔ��2o������ͭŪ�S�2�Y�"���?&��~�*�
�i���wHKgփ�Å݃��C�HPe�E^+�I����{��;t�]��ɠS�6����/J�d�G`rP�f�RˎDvGN�F�=m�8��8�=�/�Pٲ�ӓ�Ls���G��]Fe囿�Cbe�r���<��8�v��x�
+VI���@>@Mj�p�!C-����Ӓy�qR���O2����$sj� P����ؠ����"�n��5�r5�*�.��߷�.�T����>q|-j\5�i���ҸS1�l��G�qo�Kā�:F�����Ԅ�g	��(
m�����������ئs�� �%�:,��ŧ8�����ǆ�����O:��m�q���ߍ��Lޜ��'��傀ԕ�]6H�OE	y-���-��b��W�П��]������l� H�Lc�M� {N��s�����-�~�.�v�e�H�6��ĲυEl7F�2�{�H��hu��)�9����j��h	��ЋR8W=d����40�M����j��gZ*n?��D��0���)���(��|�م��ѯ��]��:M�O��;y����=c�V�WEuT�T�|����6)����B�� �������L��\�c#�b�V6Q��pu.��8\��s���Mu�	���>M.�O��!�3��6�����6aXKo��cI�"�G��������
J91��N1%2_ɁiiF��q���~i%�)�`�<ɽ)��&��[�._}W	�(X����=]�j>��@��P7��^}��f(�� H���.�?��ٰ��̄0ɺu�P�[9�ho�׹��Y��@u���ա��*�L���S#��*�<��X"����s����]$W��π�ec��(�f�>.+�Z5I>A'�x�":v�2������^�:�*CO"e�5��y���,7�X2;T�>"��φ����,���=d휾���m�VWn�%J�a��5:���:����y)�%�/�	y��Q�R�V��{��w`;�f�r~�yr�?8�:c�k������8�c�S�Й�̝��*R�$H�.T� �lG݂�Ԏʯ��9�~/�܉��/F�p�h�4R�d�.l�.�oi�i��_�T�5��@����]� �ز�h��S�"w�2\0�H�!I�VEr��v���䛋K�.�l�:����2M����������'�2�N�q�/�م��#aϕ�i��Q��?WS�.e�wf���_���]�"i����|)����d�_2K���0	��L:���OM�c�N�g�����.B���q�Ώ?�x�T*���a���D�ӟ�J�_!���Ï{6�r[9��Ѯ�4 k(|م�#u�ak(�g�m�H���[�Y`Q�t�� u����6����"L_�6�� ]y3������q�	pPAU��@��WB�����g��Ńu��������ز���W��ۥ���~F��;/��T;r�>~���,0��F�T77�͖��S��e�!9���a~�iYe�}�L�֞2��?}t��;���(�1L�!5

�;ȞfI���Y�)�v��v����xt_�N�d��r�f�td������[ѩ�R6���ĈM�@�i/�Ԇ�s�l��FaBW��5L:��7T��b�C��r�p�/l>��b<&�J}{HV�P�o�myq�Av��#��f� kY���;�2��d넜�w�x]�����N��"4�cȝ>>V��k��TS�4��*_}%;.#z\"w��i�k��n��[leE�m�Wi�޲��t�����V~OK������鯁�g� ���&�Z�+T�{�'���n�]����U� ��BH�k9�j��;����zB6}���y\�z�p�h�W���y�`79�V�D�����t����.�lH ���$��ף� �;L�&�
�� ���C�������c�80��9��v"]���ۻ�z��9+�ȃ%��'���ma��o�؋[J�N21��W��#�N.-�����5��í|������c-yo��@�0��N^,��Py�����O��T����@ۿy���v�L�˂J�gf"�BL�@�C��O�;<�o�_�H_�D����[�>�����p!kx������n�������{v`�Ј�+�SZ6c5����}��M���F�n>�|�ϝV���1��1H8��2��(����K��Glb�-Ħ�}~�%+�M���S:�rzn��<�����]����Ci�����-e5��a��ն�߅���=�r�\4��J;+n5�����L�>����B�5T��;k��5߲H�=��`.�"FbK�U~{*�N:Qw��+c�֍��]޷�ʀ�I���ýGk�
fH\i>%*eV��_Ǡ�}�t�L^��5
��ne��Lk�h{�����M��d�t�WD0M8��7H�9$tQN/�]���cp�j�2)�6f���YB��d{��h���	g�B�W9k޻��[��ּ�c�:�fha�m5����*�m�H��*����O�ùgF��f�@���?_GR3�V���v�4`/2r�~am He�|:D}ia����8�<�����a���S�L�L�tT:v"k���{8P0�K�ƨ�����s��B�]$w�,����Qd�2��3�Ȝ�q�Hy���c&�)��#?J]^��]����p�hPx��s��u\7o+��o�s��tvm󱊷�T�r*��wOh7�q�r,�;�Ӂ��H�%�]�l��a"h����mm�D�?����'�[4.^$E�/���J�����kb����򠺬�H�� [�G����H��B��i���;a���ۤq�4�Wfy�r��~:�gF�f��jF�<�3O��R���L|�\#`��e������E���ĳ���W�e�� u!Z��&TS)��x�nu��4��B.XS�\�ͦ�'�Q�o�v�:N�-$N��fxF�n�<G�p|���f���h��'(!z~u�6���q�T�|e�_�T⏷Ԓg��>��cc���R,!\��Xu�6��]>Q�~��&y���S ve�a+.�d"�"B]a�:���K<�YJ�3G���$�e
��O-�㺫�p��v~�_\1��Ԡ|;gZ] �w����*j�k���mx ' �������U��Ӣiǘ಻x��6�6q��4��-�������jf3�o�"���Y���o���{�O~H�I@�(P������Ƨ�m�8E-Z��=��r\���L���IgG�N�����A+&���N�x��t˘���D�@��}��]�v�^�/.%���G���bE��ᕏ�!k������V
v�o�4���%,|�o9���O,�NT,����)�,�(��YK)/���9��R�O�����{]`�}��_yo�W��E|ۏ�I�����3;���+�4L�Ҋ���fl��t�Ǉ~y>}��+��PH��^�b�Pu�ҽYU�\���!�<LhB:>��ߎ�-Bҕ|%Jޛ(�R�Z�sOv�a�b�Nr#������ZJ��JG#`"��j�6h�e�'���Ϻ�F�W��D[c���ʲ�����32�_��zs�܁���"�ݥ�o'�VA@s�O���nVr١ى�Y\�~Z�֋�u5T�w̡ku-?��x1Y �m�S�}���/\����v��!KNˆZj>σ��J#.�9D&x�^D����A����X����`�����^>�=�ri�v����,���D��CV��H��2$�	�3�h��
����a����f@�uk�<d�Ϊ�P �\r�a&��5��Hn�&� ���ݑ�_�bI��/�+��w�I�өl	`k�W�fg��e�gks�A��C�k
�V���2�$�)I�6�-�R(D6ZJ�.jstVkSKl�6�#
gx��7��M	-�X�TJP�r�������\���m�f^~0�����Z2H�C@���g-��
�c���Է�֬�$�=�`)VY�2����X:��.f� ��=�-��T3�\=��>��a���/U�7[��{Y�Q a����5wI�i�����^��R�Z��_����i=�?�ܡ[wI�l��Y �BD��������a[�,�����dEI�i��)}�`�W%>�)�m�4U*Ρ���EJ
C
�q~��v����Pk���h�;}\�q��!`!o݇ˍ��'}�A|��LR�b���0Í�5�yݵXB��h��Uč���+v�]_+����2�L����d�Mz+_��u�'��4Y�\'�3�"�o�A�q�*� ��.yM/��7&�W�1�.���rrԖ�Z��j���*��K�I��y0F�.F��ʷ�ŧ˹.a�}���&��yJ����� )H���U�MN;���=fY��_W�\k	��I���q[{�=�kv@]�4k7�\#��l�8���O���*�Zsmp�9����@�S�0�33x����oz��r�\H�~��K`'��M����"z]=���ln�q��O����a�1s,#�d�3vjӬ m-
12�Ʊ��3%���~�B+��磳����+R,���C��D�_@ $�͗�(z�.o�������i�H�4�׷�QN8���A���E&��IyX�Qm��Ɣ2x[��6��n7؉��Pm�)r�x�߾>!�Q2���,-R�����|q�/�wM�H�b�V�Y�����1`�M�"�D�RJ��V�%C�1#��q����zD�[�}X-'A,�=���k���[����WX�g����v��ƒ2�ZlW�ty�����k�����P��L�vo����5�Zۊ�����o��D��V)��I@��8���[6�T� 
����|�3C��Aqx�*�ⲙ�t<�<���ɣ�1�vvP�U ��|,�+�U*���΄�-S)M�RHNzCA��fh�����>�����v�d#������>���ð?](��N�˯ǣ-F�����֎iw�*#�9�p�3Ξ�L�i����ؤj�Uq�Te�;�{�b�[B^�1��y���9���$s,��_�**X���d�i>�P,h�(N�b�\�^���XF�����%4�{�q���N�;�CV������\�T�]�9�}�G~���ѢjH�Z&�g(5��D%�~'����nm�;f�^�����������y8v	�V��m0���p��P�O��I�@�yqX����E��	��7�� x�R�#~��ա��k��A��m�:�@��k��?>N�A��\�W��<|_�&��I`��bk���hshF��_V�H��9�S q�����!o雍X�+���+>����i��.E0t³�s\Զ�wc��]1���(?�a��HY�s�n�a�F,P0j����EҿL���r����َ9;bHV�]�8�xhKU~q��J�&���s<�x�@^0����2�{�9�ƣE �K�J���6;k��yP>��LK�B�'�C�O��9�˃�-�R�Ѵ�0��Z%��Zl��:�ɗL��嶕���Z��rIiHO�wp�;R�=�)����_Z����p�ȳ�937��L�����r�0�:�o�C!{�#d�kG���Fy�����1�-v�6á)�e��D�P$.R��w��H�SO�n�&��T�:?�!?�m��?�� ������a+U�]f(9�Ffv3��x�����r�|T>�덈T�������AHa����$R)��@��q�D8US���qj.s���T q_mN����J���P(�5]�1\C�3�8Q�#�F^���/��+��1O&��~Tv/�5�j���.������)>͌e̕e���ZX�Y��S�i��>���9�@&��Kd��3I�,;�~����K���\��%�pa\����i\0�@j�c�'���׬�����|�
��7��_��am|<����S����K�(����8r�l+ĩ�T�Md�z�a��nm��S���QoeN�`�������U'�q��		X�����C�����t�۸��ӕ�����DU�o���V����j����c	vn���&��n, ���!J�x��5N�M��_Ž6>	�n
h	�3+;�ز��&�x�<)�a���E��F�@��K��&[���'=3��]x]pwj\bb�"ǩی��d���^�@�gZA�=�Z�ʉ�i�������)p8�F��x��"�ӣ�Q$���<�j{ݦK'MR�(�(�q���U~?���!��1�C3p^b]�<w�$c���j�]�iD� ?(l�AP/�規�$����A�j��!]f_���k>���j23#��������f�O#�?�b�~��n�f�`w7߯� ���#K����,�\HVyY���ù|\9���������*B��0^����j���]�ѹs�s���U�GBvC�n����4�r�M�M=X��-�ټ����������Yo8ӎ�v0@G��. �.Y ��^���,�/�ʁ`Y�4H����I���Б�W#Q;��ҏ>+�	F�*L���y���q�����/Ys��ʥ;�g��і����Y|鱗����Mu���h����=�ܪ����+<s(�D�H�h����Y`�Q�\��7:]��k_PX^"{/=��Y�W��'�z���򞠹h��1=�4fL��f�cjs�d�����rBJ� �b�~�)��0�� ,q�~���Z;���v.͠[�]H,r)���TwG�FH�*7�>V[��#�\躨�f�xk������iF����%�~����;5��d���=�##)�z�a�1��S C�h�+�������[���+U�[giآ�>��x7[��m/�*'�_v�Q�˽tܗ�N�5�!��o6�ep0�f��6�M��8vo1�����}�pW�t9���)4�-�pe��ۖp-������Z��tT����62F|�#~!�ݪ+��k����9��(��WG�c3�_�*5+]�tu�U����}k*̀�v6�\��}��+��,xl�xW�l�!~j��ie���t�Fe��Cj����B�'@�����86+S����J���/DZ�V?��N�XnV�<�bՌG�!+o^�r��"=#w��P�ȼG������O�������ܱ�b��C��� ���'���p��͋�)I�;�L��!�[g�F�)�O�vZoSk�ݣ����ƾ?=��ݞ���n���`�����B�w8�m���P��% �H��r&DxbE�U�0
���`RLLlS�*VO�����+��9f�G����L���4�7��
�rX��
���̀�c��'��CJʃ�NqRa,�9%����ǹ!�reX8�͛�򤺧H�^ �c�h��`1�O����͋������7\�IXl����3_bE4fzgLy�E��E�����sG9qH�k�ꔕtf�~)���GI�=.���gv(ԟ�5Q��K?�[�KJC�N��nb��'xف���R]F.�.L����\�vH�h��=��&n27=<��s���TOG-�2� X<ƓXj5GL�ֆ�{�װ6�$�|tG��@랃�����k���pW�G�@I��
�����Ldl8�X��&RM�U�Ӵ��h�kl�����T)�Ahx8����N�@a�����ݙ/���w��%��3k��!��`�.�`����cr��S-�q����x�|�D�,�
v�;A��tt��\��+Ǭ�?���o'�1�ǮV!�A��m&�єgQ�z�1�gl**m������^�`�9��f��c%�\�׼��|��I���lj�X�����H�� ���Mvn�R���I��9�z3ME�Vc/K�bwY���`���lF9��~^���@�-������믄Mq��|0�a���k�V�-m��g�/��^MZ��5A�*n]#��_)*�R��N���"┌=:����u_�C�u3B���l��TC MA.T�z�?�Q�!�{�W��W�"9`w��4���ߏ�(��]	S�� ��,{#�.<��I�c��."�WD���8��ȏvm��FW������+H��3��2}w�F�{�{,DE�yL={*̇�*�xhx������;�,8y.���H��O>��TI��FƦ`��"7�D�q��cɣ�w[�ldd/#4=5g�H.�r�ЯmG["�@�a]�.���jc�$�R?�e��F�=B��wN��}H(�5B*�v�}��p�5�p=˷�x'���\�YAg+K�CS�x�8(���I�$��&n,@W�����n=�K�>�m�{0jM% �,j��,����U�D���uP��Q�x��u-^��~��w��F��;��z�dh����<;��!�&�%;8��c���(z#� ��]TR�KXͰ�h�j��ڕMH'4�10���Edo�Ml��D6g@#Xؾp�YxHf�.ͺi�S_��e`�ׂD��,Xc�(����G���P��T+��`�� S�C=��TY�W��_�~��4�i���hX�|h*�4v2�?�?y�����r9>�nQ����ru�� cJ\o@�q�^OAV�l\]�q2xx|��q��#�׻
�!��q�����OT���ni��o6d����D��
������R�GN�m�:*=�ۍʎG`�|���i�R��f�V���d��$ڃ�,7!�7;��a�%�k6��Pc�E�6���{3�ߞh(B��k����>~�&���i�P��P"󼵮�;��/�����NR׵�ݎ�8�|��C�.Efz�O��h�'Lѳ�v��Ie~��z,ذ�g����T����"���C:�����1��,������:�ĵ�UzB��w˿����}���: �G�����}&�|�x��� C��5��r8�i~2�V�= �NT�b��Wq�@�x�(>t|h��o8��/%��8GW� ҽ��~߀��Ǣk'�=�`��3QC��@���]�H�8�L��5l9�?��'��wJ=��|<�5�ğ�˲��N5��D>��܌;l���IWs�@�K�e�ů��P�3J�gIjt���;a�3��䝅�)��m�`r+��k�߲��͛�E��f%���C4ێ��k����k���_c;IYI�>֒�:��-��G9��M��L��*�x#W�.tl�7�g�?�����-׵9b��y�o�nS\��^���C6�����'�_>�X<!�D�ȭ�t�1��@$hOO������j5�a��m� Kc��G�ͬw>�t��l��ǳ���z���Dv�pD�\����+�Ӂ�|�m�72����ݱ_QN���7(��u�gy����Mqt.���^��h#��:V`Hf&��l!kڔ�c��t)�'tcu��4�4!�aU�ko@��
/�j(�����hBz�����彣��a�u��WM
�:����U�����}jJ�`N�o�1'98�c߳�{�l(���hh���*��_�����J���w����GT�?���K���ҍr�v߶�f�8��1�	���<TyW8��QVϛ��[ר�n���,�Z�]�t����!aޯ��
.�m�X)���d_���a"�˨h���n%�XB�=�v[)A�f�H-ߥ(��G�{��fp�G��鉨��V&��n^�o̮[T��a(�R�D���0+sxa��$�ِI���0zzjQ�>���+���,���t«�D���~&$JZ�n�:�6EnOKoh���ë�w�D� m���/G?m1y���B��5��S���r���g���(���ń�[�����H��Ӏ�a3��#�Q�<�u�V�G���3so���%/�y[)q��.`�6�j�.i�a���mlG���������p}�O/��2��,��*�ʵS�f�A�Y-Z����î����&C���6/�W���ס}?���)|���=��!��]_"�-ٛ�6I>�`N����NS.		���5����� =U�t��,x�x�+��������u~M�2���X��ͮI�/�1R��W���W��Y^ \�S�z�L h��%�����p!�s�F���}�_���^���^�����^c'�;�ί�7R�¾bJ�ܛ6�
�O��,���Hz�/t��Q�3Yx�3��*$<}f�[8h�K9�h�;/�|\H���4���b^��~����O�&K��~}�D�3���q_+H�x���j�F�k������梨��oz�4 �NݠV�m`K��mo��o伺c&7G%�_��d��
�B�c�J%-���|�ӵS>4�뿣b[#�h��0}6Ȅ��,�T��q�+��]1L��q�_7�(�J���f�M1��`�A ��Q����K�v�MF�	�������"��=N7n�{w�Y5W5��M_���5���7g�v���2�!��r�b�'�kv8{7�K�V��jc��>`�H���])��&^�4� r��?���3;�|!&��coz�{�e(-�u��n�0l*+��֛[�I/�@����v`����y���|>d�R���9ۗ�l��,1 �2(��8�}�*7� ��e^  ���GAw�_%����+�JU�Lx�]��O��A�  �~ ��X�F�Fт!��c����|Q�(f S9�N���@�!Z��r1�e�����Y�B{qqu1uq��y�x�f<g�%ne���}ʕ����<�x������#����]�Cg��9@��2Dg��w؟�}�iQ���-(��>XpCf��=�)����jD�Fd�y&c�J�o�oק����,�0�݁
�����i�O�i"F�{w�����j����Qtʬk�x3l��~�?E���͊������czq1��'�z'o���ڗVS��0�e\&G�o���T������+������	���ƾ������q�w���xcI˖��zʂ*�2 �F�w���t�4'޵aS�R������s��d��/)�W�{ð~s|2~�h=\�^�
�����(���/|D�=����Gd�o�����2�<r5�a��('��.H�_�i�h9`ww΍nbc��b�����wL�}S�w�Gl���G����X��	�4��/�-DKsHw0f�"��6M/�~_]*:�8f�CwB��������:[ڎJIU�̵�-K�q��
���Mb�ĭ7�������I���}��k6:��g��xp8ׄ5��5����ǭB��hԬ0AV�?3J�~O�y
I�2�ՠ8�s���-8/���u$��LUS�CZ0��;�r˞^67�t4�4~���R���w��[�Toi����o��UH[cG`�,�f?��fO�ö%�X�����m�ۗ*�7Z�+�"��A�`;�3��WVJ��!�dc; Y�8�q���ӄ4W�Ұ��g��46B���7�a�:T��HW� ��䴀�]%��r�>�z�O�̈́�٥<����D��������Z��L��ټ�����1~��KO��#�f���e5���R.��_�xC��z�4]�b�䛇�d���?~�5��w�:we� еy
;<��F�����ZW�V)�s��_��k�;'L&Q�N�[oV7!��Aɇ�3�3�p��%*�7��F�x�����?=������k�����x�؝�$�K�;��<�{[9i��?� ��kK`>v-��QĀ�Q�+a�V�����]Ģm�N���|c6m����d=Bƒ�nf��a��z�>����	z͍�a�;�[�l����yS��l0?B��gs/�l�q�6�_������H���ݶ�n=JV�m�����X��$�=/Y�#Hz����0�<��{sŤԍ�����kU6ĬN[�����OR�6C�ASZ�S�x3����]��dFwO�1pC���';��aF�S�o��`�y#��yEk8�W�]v[���N޸��Q�$�*�a޷-���P�*ꉞmAa�vR�)�]?$���z�(m�e(�#��Xs��^\���2�1��Wݜ^nQG�L8�����`��?���/�+�,U���k�ԝ�0�h���i=5HdeN��S������k�(�{��
ۿ1��D��uo��x��q�mK��� ���
c^H��0�os��Xݳ�T�E\�����<ɋ~3A�mo��$C^����(L`]��B!�	��Z=\a���jС���s�+|�Q����$K�ro�C/�=ŽzQ�Q3��u	�cW���׽��� �RB5�f1����:�2ͧ~~�V}՟*�?�ٻl`�g{$`�u�)[&��3��[p^�9k�n]d�ZwH���O;���J߼h(k�J��5��u�ӌ8�&SЖ�MlZ@��5�\��'Pv��l?�����+Z�u��j�}nS�՟�
�(�4gW�O۩ca������8�N�u���Nf����j�ץ��%���B�+�84���i�V[a-:Az��k��;ߗ�%�!C�$�`IQq���>j]�f����K&�S�,��Yxp�i:�g�z ����o��5��m��ġ	��%��e�1t詠�cg6q���[���t�v.޷��6��#ͮ��K� e�7u��y\ę����E�,�ʑ�.�ĩ�R�(���RoZ���6�7F���ݫ��nBjo��_f+�W�x9�6<��1b���4}�f�`��ii��J���{��$[�����ڢ�[*f�26������Y?�5�4Z.�܏8n/c5l���7�_ʶxx6أ`��جw5GV,�~�!����~����v�Ř|q�=o��y�R��N1�:V	�y�������ø�$�:��;�of�5�,�^��-���փl����j������d��!'��#>nT�������p�K��/�Ly��ĳ@���-�6+#�j��u�0Dg�\�p��^����D��5�ٚ���*��C�;�,��>�|_��ڨw[�b���%ΝC7�fA>�����|rH��8�	�C�1�RŻz����r�9��n��+���QN���7��]q�$k�<u^Q�E�v'���]4ޞm�r���6` �ܒ�:�����IU���V�C�`���'�P����jXO���x8=`X�\��qO?�)"{�Ijv3�,�O�_�c�G_�]�x�X�|V����Ԧlf�.�oUn�\����',�r2"�Os�BZ��%�a��ȇ���] �������J�	"����C�
._+�":"�����u�[�R���K��,�r�?���.���]���L5`&�]��I��eW:��l�\�Y�V�5dKTߓa���BQ��Z�CU��$}L8�QK,��qEc����̋����T4�;fYs���z��=~8E�;a	1*.(��:p>�DF�)�vuʘ�8&X�~����)��F!j*LR�H�#���,N�Q��Fn�z�xx��5��zw���UN4�ߔÚY<7sֶ��4M����u>�p_�L�l�S�y4u����\ ��/;{��#\�1[�	�O��`]��0ZP�~��K�a,>����N�����N�
T�s����l���&J�����'J���E��}�O�+��� Y���{�"�A�۫�3��\�5��3�FI�����F�a+j��c�YC7*�<n����u���c�j>�m�@�k�y�[�$�j�wQ�U�%�����cBD4�,Id��I����	�d��N��J8��3���< ~�YDX�{�f�I@�nX�w�ׄ+s�֦��u���̨#;�_� `��\JQ�����O��;�G=dl3��r�R}٦�bi�{�u��0�ci7�
Ng�\�"r��_�(�#�=�o��r�O�����Nh������}�G^��u�U�^UU��rpv��^��U���z?*����w,/�̇�^Xֽ�Oo����D���C�$�b�ҊA�d��ڇs8�n�=N���6�����f��j���5�����K����)��������ܭ������������5֚r���{��E�#�L��?X�Ҭ��k��Ȇr���-=��ȭ�::L�,9�ϋ�fI!���F��i~Ξa:�'�Pռc��`BT�;O�%�����g�#�y����q�r��M�XqY��ͬ�cu:l�ޓ�r��H���L�0�d���@H���zPxsPh�0D��9F�S���a�m��?��ȁ�]�j9؝92��- z�� �fgk��q�s<Ij%�h��gDh�ѡ�6��4wN0Ee��'D��HV)�韊ټ��^���g�sv��?�D�u��O�U���	*�'�xf�,0V��O�l�/���?�^�_�@���@��r����{IÍ��T]�'	��w���Ɠ�	W�������G��EKdԉ�-�:������r���hb��ݟ��DÀ�)T�kL��4�m
���)]�L��HU0�4)=t�;5 ���z�3��l3B4nL��R���v~s�;�No��3�a�j����u�Ʋp��5�~�K���c����d"�ibe�rzhuk��q��-v�L!�t�����h[��c������4C^�Zm�)� �d��G#�B�Y	�O��p�{��KW�g�����Ɍ����,Sv^�)O��[�����V�����5�e������N?�"�8���WeJ
�H+�?�B���m9��խ�g���OS\|��|w��ߗ���C�Čn��J��jTJ0�� #.h>��p�,�X��B��� �ː�����b�V�]� �oK�?^ןrjf<#�4�������]:�ԣQs��ĭ b��pat�6��� JXj�s��eM׫���
�n�}�Л<EQƧ������w=}*��_m����ũd�	K��ւT-D�P����9�Ke��^-;�|C�ս�$�>�n�@dCt�&9��i�z�S���7��.뚦Jo(������u����mڳ�ː��w)c&�6����O�"W6�y�&1ڣ(DZ����	���?�+�ǀ���;1�}�λ�C�1ȏm�;��nч���g�m�k���c�U��X_��'P2	�'�����{�U@X �č�A�Zw>X���KS6�)^lI�*�@�;�D�� ��̫%�4����(�g%ܼK&����ekM�����B2��r��AGDNמ�8N�dGx�!��-��u���&ɓ���s����qO�i��R�#y[#��$Zh�Z&,�mσL;��E�{��B5v�h�VY��܋�^��ksnԻ���ґ�����t5�Q�?�"ǿ[�Var��fB�ٿ��o��{"2)��$���Cw?o�N��v��)|CC�Xr@)q%���5�\���9�q��h����^ҞFs�v8���`s'	���
�*� �ڝ,�vp� �ޥd��Ȏ�=�a���@U�R��p��O�i^����4��;>�8e\��Q���8�M�T����T0�_��9�O��;����,�v���PLȂi�%�7���1�Ҕb��������Ɵޭ�EUJ7���hGd˦���Y�s|u��E�n1�G%.,�b!QP��s��=0/�Zv�8�ͧ�*��6�ߥ$������l_#,��_Be��>����D`���Nο��b�ګu�o�PG�ɟ���!M�'�[۸[3��y6�a�1J�@��/��l��F���]���*5z�/����/�~�N�{��:�ӭ]ş�M�G�Qe��9B5})�F7yi��rb� %z6v륝wZ>@iKL���R��\pI�z%N��*D(C��%z�o�H˰��ie�?]_G�b=2�ņ���b�$7�\{�bb��3 c,�M(��m�pB��c���TT�z��pS!�8~���nƆ0W���U����OOĭ�����=g��߼��u/�d��_=3ω6,��-�`K��'�
҄�9����C�V=;�I����j�<��`��y�>Ӣ�,��%]_[��Y�i���1��b�h=�A��r�Q��#�Y�{����+��ӥ�A���������w�;I���C�����i(p���|��צ��G��~YN���̫eb�LN�LL���q72�ߚ�}���&�����m21A�;��	�y�ȷ��@���$[�Z�c�o���IK�>~S��o4C�7�_�/1�%��}$�w ���3R>�U�JC.�<9�ꈡ6��c�O&DD�ק)�����~��zݝĊ���Ap�\o�,��pt����rZ-�3Щ����\(�tZ�4�/,�Xj��u-��[�ȗ?�|2��i>U�*}��vr+�d��h��)�;@hD����5�B?4n��{I���x��QV������;	a�_�s���8�Y����
ڪ��b�o��j�>z�[ IƇ��Zg�g]�G4�p��o���{~!��t7��C�B��2Ks�m(H�p7� #�1�����.�\��_ҥ:�y� ��fO\.L�s��['��=ԮW��`t�A4�q�|�=B(*�N��z����D�Fd�����pZ褰�C�N��u�����,bgԿ�\f�LE�U���7u��X?���L����C��T������io׏�̩k�W#��w��@X_ �����6��Y��Z�v
�s4s�f�G7X{���Frt�S���	̉w(�Y����SuC{3�붶lu��i95O2��/�r�9�
�F��>zu���l�p���J�c'*�O���Qk3<�*$z��+j�������\����j��%.�n���Ѓ�@�֌Հ����} ��c�(��^�a�ۉ���G�>��˓�j�+��b�.�ݓ΃�7�@!���X�_���Pg��6�����U_�dD����� ����8<�|㌽��5]:� �q���'T�B�N9��^�T�JI��'�Ã/�;]���^UZ�Wg/:���奴�u(.Nd�OEh�W-�]��.=NY
�Y.�}tE�9����	A�	���#��i�����'�n{[#,*�l��mY}	��Sogp5b���7�p]���v�82�vVBw ϑ����ِ!^��b��D��w��p��^�fV<'���5��*KW+4�j5�N��N��OU��Ge�?� �F�O����x�᪺N�2�����!j���Sغ7�x?����k����a��
�i@zk����Hy���WA_L��/o���U�G����0��P�`y��0��Q�m�ӭ1��W�$�jtR]����E����V����G�:@���d����.ދ��w�,�}�� �*����r1�ڗ]�"��q�B��Tvm�5^r�l_e`��?��d��b�T�B��cdG���#8Tt��P԰���:�oJ��<M���O8?ݩX=�M"k��u�\U�g���2s>��L�y�����7"�k��~X�R��j����^��j9N�~��6�J�ƫ"S�ӍgS��;>�o��t�by�u9D��Q�鷖�q"��\�.V�����0|�.}�Q�&��V�Q�ʧ2/OpQ��w%�%iXt囡c�~<�=X@:	��Ց`�.[?��C$ �ۓ���_�Y~�®�SԮ��i��u���
�ŵUJ��2��O��I}Q$�e-�w�7�%�sg7���lE� ��N�i��~��7m���8ۖƬzE�~��Ɯ���^��eLx���z5q��a���\��9��ɐ�|.(k$Rݻ!�=e��ˆ�h�P�;��z���#�������yg��LƯ*	���7�����uE[�#��.P��ß��чg&�9�J�^�`��&���>(ʧa�Ȑ\�6O�w���/G�;���z����Qdʹs��5X¢»��0wj���@^c����^����z������#}d����ܰ�x�j||�F�=^r2�8��ߞ��F�?�͆�N
�gp �����wt�hW.�M^=R
�/�7��Z3e�+�����y���ݫ����F�D6�
���Ŗ	}W�ƚ1��J�6z{`g��'.�f�n��o*ǿ�� ����Dw��J��d(��'utA �e@v�I����1>����NR���]K�P��+}�z���QB=� �S`�uI�������1��K�N�������	��n���8Z�>tX�)�V������7Nͭ�vV��#^��nPj�J��D�a�O�E�	�g�KF�糇�y$%g/�9 dN�F� >�ad�������Ğ��R��RT5�ī�����~��f�|�k��/��F+�O�lF�P�D�V��6ț֢��q*���`�n��|F��ʥ�bO������{���Vyr�[�����Ŝ�6�U�7��I��܂D���B�e���6�gj���(�Ԣ�OC��8+ �p�!9���:�-���?��i<�R��u��iߥKE�E��nv�5�e-�e�����]z�ڣ�x��;�O��̯�/��-2{O��N�!m̖X�+�1Z���}pxN��8���ίbw��֠�e%X��ױ��#7�|�[�����To$4�(Yk���2h�w�.V�3�$�f	��D�r���k��-Z�����}�חV��l�f]� Y���v���w�R����Wޥ�D�AzRg�ugt��; 疵>�%�?S��F;���!��Ě�z�	�O�<�V���Q�g�(��^�����lB�R��o�RGp
A~�L_v�K��w�	��Fi��{�8����mk���i�9ѯp��md��3�W4��B��2Q,Qpp#Sl��!�D�)��l���8�d^@9!�;1���?��ZWr���]��IǶ���l�����s��HU7�c��|'M�k��:,�q��^!��ι���`�g�s¿lȗ�^�|�f�np�a�OݐP8��p5\�S/��H���v��ŦE�)1Lo��Ǆf��a�#ޝ��T���s��,��5,%	d�Md��>�Ev{�I̐�+�훀	�r?Rѷ�$2���7�*�Se�,�9dD2� 8�����{�(�]������?"��.pd�[�Em�G?.{?y�V������>�;�H��|���b���F'��,�7�m7���qD�����]�z��3x���� ���!��,�bF��z/�9�O�q�m�v��j�Һ��Ku�%�;���z%h�W�NV�x��2V��	�����SF2kPB�Z��84lz�Y�ǩ��=�0y9W�e2���}�j�k�n,T��U~X���q?�{R���u�'��O�;J�������/B� Zq	�\��WPֹF���{����%���w���E�����/�6&Ԛ�bK���sV7��ܧ@&�����_�%)
0��UÏ�v�\y���J+��4f'�xA}eB��n�k�!{&���}���s�G�[�!�/H#0̑ ����`�H�ݙbbV[*:O%�λ����>��7�E%�U�V�0o�9}�K�����w�%�NMo��������h䋭ݔI��1��*����Tm�|b��A�>��C*Ο��˪�Yv������؝>|�R\ �9�����j]�f�c��� ��~tһ�g���R�������~�<�Gr0��4�%�����H,%�� �3K����LQڴ<�l�@�旻�74�r�ٵ�)m��\���,�?[���U��-v��|�z��o4 �D��6���$�����s?|n�����u�+C��(}Wڞ��F;�Z�)������V��l/�rE��������t~�G>.���j���O��{q�bA� ;���P�78�bu)Ȉ���;��ļaA�$އ�a/�aJ�|�nu��-K*����r��e_�C���;���]6��쌡�/��'�T�Vh�L��w�f��B�hP
�Ֆh77A�y�/>�_~��~����V��i_�����Kj,��gf�|w#��B�0�Bև�q�)~�H��N �ƽE�B���Wݎt�A�D2幑��t��lx���U�.��a_mq;�9^�6��o0�NS8>��,�z����T�ik�]��C4�~����)xd�����~տ�+F�C��p4-��݋�x�)DrX���V���j�&��P�t�u2x<���8�^��ķ-��F-��i7�0���֡�����Ă�����y��ˀȉ��[ֈ!�F�j�I��TsB^���-S��q1�ޏ�q����5�@7Nq�F�s�	G�_UY����zoq�T�ë!*��')(olr5�I`��$?�'"Z��	MI���5�oTA���v�������E=�ƵF$��'J��ӎ.���HB�:f_�������o� �Ż�6�-ߘZ�Uie������o�������o{��1 g����>f6�[�빖�w*"�N3>N�g���`�yde�ƃuZ2�/\�!����r���?Sr`���ɿ�����Ҵ��o+���,_��)2�QM��ƚ���)Z\�0�j�j�;�k�Щ�alX��������2���r���P�q���!qW��U1�X�WЦݼ���mOrX -�^��ƕ�F^�0wW'���*U)2����Y'�I#yZ$�!�k�XJO��b��|���ы闡�juē���/�h-?�XC�2���Kj�ṋ�-5�Y�Tͩ��d�kQJ(ev�-L������E �'����}��L.��-��z��j��r�~A�w�P�H��tq���%�X��o���K�Al{�Z�5����l����Wr�a�d�2Kq�����L�?0�bz��[_�^��e�x'E�2�S�k����P����=��ok��P����tġ+��+��Qhqt�׍�Z�o��4$"�5d�:Mv�\Xa]"ݡ=����Ζ�V��(N���/���Ɏ�][)o�m|�p8X#���:� F�_nP��R�yn��
���F̢��z��>��U#?U���w���ն(wO���H��G���t�gs�@��	� 'GQ�F��$Adn����ա]�܅��V�x0Ľ�:q��I1ɮ�����,��W@�]o���X/�v�����}�r��~v3���_���ݳt�M0dA�W�5�
�f2Y�w|�Z����9�%�����!���ƚ���,SƯy��xZ�E���K31��}Z�[��1n�0�o4�h��%lZ�����0U����!�#?��샞O �Cn8j�]��s ���N<8*�ܣ[�3��z��Z���W��T���2��2�4^�X8,W$�����%��裎󟺗S�<�����X��)��[&�T=�2e�������������]�����d��O��P�s���i�Cx�)�;k�{�$HR�@C���4�1L�Sd	���yD�Q�Ř�g�11Ra�J�0B�])Z�/��*^��}Qm�1H�C-s�W{W�5u��=��5�3�*^=m�=��B$��������Y� �z����/F;Z�[?-�qy;����b��S�,�� ��Q�2<��z���S�>Էw���5��P�en�k�s�۪B�cLƸ�0w�(�v3��q�Q�V�|�o�i$0�3����,.Cl/F��oۿzf�k%��ᡟ6�w7�EC�lF�Vk�ng��%:����W�e݅ϝ���bzd�f�j����� 1ԧ�Ia&Sr3&w�?�nk��������X���
�溩V9?�S� ������G�F� B�+� w����,Y��x)+�Uf�1��)eS���i�_|����M,�����]f��f�������c���>�Ƞ�[��ۉo��dA�"�56��[|4��Q��o�qN��\o\��[�X|��ʌ�?���+A3~�L�xnEt��S�9�������q�/b�=��G6%Y�{��oHǠ�/F&m�uJ�F�we[��Ѩ>��>\㯰c�9i�
�̜�4T����T��c�t��ߒ�Ʀ��U8���O��Yk$��l�=����G��y/�Vt�����D�~�j|}g��%�K�t�7P6:w���f���@����8���m�|W8�/���Ig��� <�<�{;��7�/��P���F�=�����/�l���[W�?,�-��g��|�g�m����0�[���Q���*j-8��̒��D���=��o�u�č;Va��L�b�����FX��h��� ב��]O	���:
�׹5�ѤN[�;���r������9<u����(Ό�¬'Uj7D��<��Hw޻��ml��k�G�3�LHW#�(���0�4p �W�J<:y�Cvw$��2�Y���Hɠݱg!�m�[�
�A�gg���/)�����(B��{�C�P����l��%��cC�:µxy��{�@Q{��FsmhG�]T�{j�P&�=�ʅ��+]R^�u�DY��G wyI�����ew�sz�K����c�\#99g_0Pf��(0�oZ�t��5��3W�`$�w�k4�+U�4�J<	n7b�;���m�h����d@(WG��X��'�]����W�s����@�_�n[����y�˽g�{��RO��r�r�lM��k�Ǵ�p�HV [�k��D�2r'��m0S)Rච��[��[66et:QN��[�"���I�i
s9��4w���։v�2�,tO��\�	_}��c�_�:oKn?'N����A�P�n���'�\���S�8J�n5�v�ȅuģ�f�?�a�{��e��|��ԱO�N�u�V��o�o�	S�z�z~sU�č��t9u4K�N��ò�N[^A�a}ʿ�E�2ۛ7q����2�m��ԣ�Ig���j����"�gJ����L��ߍ�V�]j�[�{���'g�>OQd�4"���վ��pu��	��.�ck�����ϴ_��#Zo?U�ԯ\8��W�<��@Q`αW�L���w��'��aW��Z�=^�m'op��w���p��1�.�iv�|)�v4�k�,?�� �nԵM:�=Ƕ�^����W�y�-g��}��X�X���I�����3_RG��w)��<"R�9��>�%��1)B��3l�GI�K���L0t��>꠽����&m����d�kAI2�&}p��i�j�����VY�2:t�{���<l����p��u�|YIܢ�����*F)��(���ԛ�7���v������bY��
1��_���Y�����Q�ޫ39�_�K�q�������'��5=�E�k�&��0e��<E���;��3(~J�����p��5��I�j�n\��c(ϱm�9u�u�F�]��<v\�M1��������84~��efҠ�D���?�?�^��ꅈ�\m�6𒠙��XR�ec#�.�&�#y�+�Q�vaū�PY~�<�j����P�vʴh��?��K��A{J>d"e��g[EՁ&e�d�	�8:^g��2Hl����1͞�
�OQx�W�����w��A�g�^s��1X��2�"��w |��B��S��,����"���w��g���W~��hƳbx����R�����VVr~� õT�99P�Rw�p��@���+¶�k�ˌ�%e��F���[W��yL?{P��(��}�yC��>�z`<ତB#�.����):@�Ɋ�il,Ak٦X��㼙02�gߝ�3�?�+��띥���)'���WO؂X�ΤLF�}U?$J�H�L�����o|��v��6:�9�I�)e
�?��{3אKa�[��Pd�RZ	OHfI5�esv�6Gy��*g,�~���j��u�w8	K�x(�z��#���5:g�t�]1%Tޮ/�pC�a��5t�P�Xl`U���_T0e�����hU�?u̥�?c��ҧ0�i����^m�{���9�Hl|'�e��eeG{:ZS:���`�G3{Gޅ��?n�Y�d���,j=���*�����@"Rr��{Yg��c{I�/dܗ5�,L=e֦�6��Opԙ]�A��,T�ՂhV-��'|�I3���[���^�O5��P�om�=�wU��L����l�>��J��׫�7mrCH�x7��L���Ah�%.�%e����6" ����F�߃�|�4&�yt�x+��@-��+��e��W��:@�->bu������F���a��W��s\g_{߼jg�z�M������b�S@=���A.o��s2D&�-�{���ʿ��Aj��L��<���<E���d�j�&G=]��j�8Y�����!���4;[AT�n�����O�'
��Epc�\'���cQ�3?6Mg4��&�ʿ,�DH\�ywDb��봧:PH���3\��qлOJ
%�fc2s�~B�S���jE£�Rn�����F���[�yn��e�{q'8��+�1�����zg���V~��H��+{K�0
Š&{Q�0��v�U7/[]-�t����I���ۿ�K�7�r�#���㠩$��ӣx�xs�Ka�ɭ<%? 6���,���E��J����Ώ����z��_���^��{�)���"7������"1I��� )V-����j/%&�Z�N���h}���X콹:x��\��td���<~�Z�������3t{��̨��FjZ� ]�o/����x�@�60��	<2naG��Lu��;�����-��2㻲J9�cE�pʣ�hu�ʗ;$���d/���ZA���o�����/���C�f�H�^+��@,㯬��Ҧ@D�h����N~���A|�b/�񸭋% �'�*f��r�����c3���mrG5PV�DViO��H�h���Y6�sL*q#�Y�}_�u��y��g��}N��X
9���0}�9�9��թjC�3rӬ�u`y���H\v�!0�j;��I]�e�,�l��+�O�"��9�����y~��)3�T�&���5I��t�a�~XtѵM�S}N�dHB)���B�UEx����7 !�vq��9A��H8��asz9 �<dv�=yx�ا`�(;��מ�3s�k�A��x�uu�n;g��G��'���i��U8�u�����%��Vy����xH�,�����w���ޘho)��>�mc�����ڝu��T�1��`;�kX�ۧ��Uk�l�w~g�~����/;ڭ�n�m������mS�E[�9�O�D���t<b�H�x�I��Hmw�h�.P$����	3�����n���N"�:�Z��q��+���ծD��o��Rog�Z�Nj�
io�@�?wH��ƅ�\�F\��gݽ�ڏ`(a�/M��6���C�D�!=c�{�%�ĝ�fO*������K1��v��]�Ɗʀ~$��a���{ŀ��~Ϥ��bΈ�`ө[�jܑ�s�I��*�8zU1.��@Ɓ�M#�Y��^]ގ�?���3�7q�JK��E��PsX&�^.OCg�~1�^�����)a�w�I֑m���|G?�w�Â��R�Ws�
 ����r�#9�Փ1�?n���{�I���t�Š�}a�T��*�/��������j>�@Z/�y�t��S1^灊c ��X�f�Y-�����6�k�_5Ej�oe�T��ɰ�U�C��XO���ZS{K�h�
�����Ϸ�Zg��C?�m���*�E�22⣍�Y����$���kPz�u�_���+����O�j�%�^�h{AO�!̽�ߩ�aW�ԻG���0����l��?�q��$v��u��+2�1�߮<3f��Ľ	�����nR�``���L�m���~|��"��2I�QnU���P��
�`iީ�Z8w��A�g] �3��ߊ�	��/p�_o�e�h;MCF�K�C:6'\�i��'b�����#�8=����aHM�x�*ߛM��),%,t��#a8��:8�o������0�}�,��)@AP��(U�~s�?����������������"Кs��f��~NյR��g��A/+��<�M��W>S0mFlR�=FI�Fe��ϐ�ن�����J�>/���S ֚o�ǋ��l��mju�R��ZG��N���zօZ?n1��H�w\��C��*��>	�gNa���ڀZ�K9�dBWl��b@�y]Ox��v�	OS�l��" y�϶aX�VB����G����a�M .��ͨ�K���R�2
6�>!۽D���"$$�ݾ"F,�|�Ջ;�
���Z��혂�L�,F�>�!.@�
�=
Ss�~]�/r�w���m�w@Խ��r��ľ��6.��N2;Pf��
ʣx�Q�}n$5e�sG�U�{�R�<�f��Q�r�gHّA�ؾ-S�0^h�����ȣ��"�N��Y������nA�������j�B=�{L*�6�Ϟ��׋��k���݄$u��BmR$J֘UY�~�Eɫ}I���=��*So|�<F�gХ�rgl �B�*N��|2(��xי҇	�5�$���Q�E�;���_�3+:�]������*�p�8�,d�m����2h�U�3`)�V�B��a��E�50�a�hy�63�>����=�0�j�~b\s{�h&T�di��g�y�w,�����T�6O���-�Ҹ��]z�	�=��R�P�Yx�~&���f���PmF )�4��B�o3�$�s��ugx҄q�}!���Aꑐ�}/ fs_���� g}�n�~�ƺ�����wՖy�O��τ�0dи<74�t�@١�����|J�xwZj��^Xe��4��I����<M�N%�z:4����Vy^����D��1�YΦ+L��~�D�~Պ�8��g������M����u󷉼�^��=x�7'jj���hw�~CW��e�S��kQ�w{ae!�]���"��=M�{�����).�?l���;&��lOx�hO"��s/��m���I0���j'#��`�����C�f8)�<)_�.v�A*$�:u�=���^X��^sϦͭ<�JI���3��`�~�M'��s�nSݖ���E���3�8z���_��0��u��+�:ǼI�b���@��A��.���WHڝ	��6�B���ӿ����;s/%Xs�MY��lVA�S"5����L�k���<3�tuLD�9`�E�"#T��-v}��1�z�Hy�W��Cl"�c��g�����Eʹd��1�m6����L>�+�Rx��7�h�5hFp2�+(��<���|���X���O��Hk�̨����s	��[�"q��@F��|k��Bh��W�%��xk��O{���]3��4�V�B�1��.�X�n�lh-��cc�O��Kk���y/�cP���ݒ)v���]�mR7�����'uS�m��us]��4b���F;L.�d<�\ӻ���-�s/��,j��B[�D������i�� b�qs) J�C��Nl�����t��3� `����SP�m�g���i�9�W��fIb�z��I �۸��*L�hn��,�O�`��-YC}�4Ԙq��k�
�nv����`��>G���X�zy�?�>��lN�e�0I��-}���)zq�2:�BA�u�*���X���<��0m�دd�$�W���[u��5E<���A_�����>!�߬��
7q���!lD�}3��扖�zg�b�ֳݞD�w->a��;��z&�r~���#�˸��O�_V�k������k����<pg�j�N�*�{�-��\4C)����5��j��o�S�Tb%wF_�Μ���v�3!F��I� �����c-���(^*j�����B�D�r����j�Y����r����#���N��
�T��:<s�oZ����O.!:���C}QCSֲ.��8}ߴD������֦�qfy7��W�xOiV\{��� �JQ*���&�/�%�T�mBH�GXMb/Jm�g��M�䄇�W�QA݋u��/Z�2`��í����x2g��>��8Z�5K��L���&��������\�����R��J���t��?0[��.d�q��µ@�v�|�����8b����Fu�B��b?��W�u,@۲ٿ��	Bh��ܦ�;a�b���Q5��e�'�7��Ky�Z�_���zU|J�g��O��/X�:��<U������Cav�˛��榮��D�x��=�����T�	�я�y-^�HΔg0D�w�8������q�M��(�ᗻ�ZƲ b�N׊T�n���;�#�>����\q3��p9��L�ߛ�1p`&m�2J5G�[��i�/��9��Ja�Vӡ"@�D����'8��w�ۿF\�G�S���S9ӯv耑F��q�F�~��XR��u(�a�i|�%(pg,��w;��.����O�X�D}L|q�
�Ԍ������AC��LL-)u,�PM��ǧG���Mڮ��w
�xD�|�y*��h����\Q�!��y�VyA�~{2��h�rU�vt�L��^%��辐OZBS�Ӏ��󠤵��v`,��ha���wߧ`����8<d1��e�[��oS�U����G��{����^Ώ&}T��v ���K/�Oj.Z��{����c6�,d���ď��VyTT-�7�R�{�K�Z����1�=�s�H+���"���j<?�(fe�a�:��_�`nF$0����ba8�pS�i��fxOs�#,N[ش�!�����,+!bHL{z��py���.��j��x�T{�q�>?��6��H�"Nc���1��!xѢ�YVL���o1��J8�$z����U�E&��D����`aSl����� ��������O����A���6YB�}Rm�y�K���JXr*Y�-Ⱦ�:�C��=sX�9�`����&��r�*���K��8�S8G<[���L-*�N�)Vk�I�P�b�!��DO3�ybM�<�[�»����}M�h��+�[�,fc��j���RjLiX�5L�2��,�����nvY}<��E.�_&j�9���3��� ҷklvx�z��&I��_�22��C:�*Z�H�$��i���So��ǖ�y]�M��?�Y�����_�����߅��r�-C���YaD<k�lui�Uŀ�f������K��z�Ha��g[LD�c�?�F�Eͪ�ۅ-_=�ی�(�p�1`%��Ũ}��[\^��:�s�Ӓ �L�/�@��y���Ϣ���2}W����2�÷W�o�,M3r%7C�+k�5�b�Q�H]��۞@[��6Ș�� ��v����J���,�CU��k+.B��as�C�5��3��Əߐ�?�x�Ec���w4c^��J�ҡ!X���8_U6kF=B�9f�/n��7���4�~�vՅc����iA���`��7R�"��i�[�'��n`χZ����j�h�C�~��_��o�b�{�]�* �M.C<u����^�ma%0`���
뎰��c �B���r�K�뜱r^��7�R !TY�#( ��.C���9�\6���$�����u��k�ם~QC��Э�ZE<e�t2�p��l��\��E�����	"���yg�=����y����s����� �	$^�N;�%��ex�ܬa4	H��&��?�^i�>i�e�1�)<,;��}�i���Zp$ㅍYT6/�p`G�F�W��B��V��#��Y�ؾ����\ӷ�4^�1M1�w��R���z��9�Y���K�[^�u씐�F1Z�jM�Tk�V�$ ާ����*ʐm�|[�kq��?�u�i��s��b���1O0�����_���֗yI�W��B�;��fț�۶R�[Z�������1㟫���j��" ɥ p�N��
�^]��_��sٜ��,���TtҠ�� :�BM�;�;��kҨR�l���Z���z��N_���[s�k�ݮoX᭐�k��5�V�`0���:��o^U��o@�ң��h�%� |��@ҳ��
�.��W1��oi�����>A�$��:�ާ�fbE�0�Uk{��=a�Іҙ%�5����op!��a�S�wpD����qJT�$��z�+2ڹ��m	HGH9�����~�t�<
���.;������h9N��KQܒ'���J��Q�J�bQ@+m~�D�ĝC�U��CS���������x�����*o�J:eS��y�r��í�sY���Q���*x�� zM����1}�����b�,�~5qHH���2�(v����S)��A�Ѿ#-����섗-SG,cM 07��D���h[|OX�R�����3�c�"?��"3"��R���+���;�e����f@R�Ý��YIJ!��0Y����@���j�����.q���:�y��e������~٧$V�b���w~���S̨/������>=-���sqY��BZ�D�ԟ�u���M�Z�)�{���p�K�N���	)}u�λ��(��i��۷���{^Yn=���$��^���
��A3�F淪 �;�-%my�i���m�Q=i���"��#�^�I'��m?Ei���vYP��T��� &��� 9�
(�ow��ܔ$�EQw�(^X\7�?�O��K;�d��/e{��x���}��#l���s߅d%P� �vg�%�uCX�L �mY�r�xW0-�S���Q�QU�Q�(�t����y(�[��;]Jw�HsH��F�n�n�8�m������������g�9ל{o�+L�8�C�v��	��������6~{� �#��C�h����>Ko ��,����Ĺ�bR�n�Y��:,��l��A{m�`랃�K��Zx�Q+r������Ov�eH�{�B�bK��I��{J�NW�L�*e0ZAL�n�c�F���ֈo��{��q��V�2����DLLDjX��Zx��Ҫ�fd��N�����u�֥� X���t����;흣�pԸ�������G�$T�ܭ���6��aa�a?i���k�Uf����0�Vo� &�W�ܾ�e���]���?��}l��L	���i�����(v������1�Ol�т澒a�D����5	�t� iƲ��Ѹ]^'�&��:nco�o����h��hh��k)Ɯ�h�e�x��$��DJ,��̭3걗��K�@��K�"�}nk=1�Tֺy����Y4m�|fi��,v�'��N5)�����B���;U��e4l󙖪��}�|�X� ,�Wx&/�M��T^J�"�0�{�C��N��ڍ_m�j�s���pc�:�*���^CT�C��iW3M�'�J��V�1�:�^�a�oZ,�:��N�8aO@)cɾH��*Y��R�|[��^x`�^��@I�"oN��!�d�%�k�e�?�?��"w��ȿS\Aن��e�4*}G�Iu��L�:y!"H�X뽐;�Q4�@�D���(�7]ؑ�G�E�'r�,�t��CזXb���\�	�X8�.;���w��,�z����*�S�9P����3��%���K(9h��@V�]¯d9= ay���"���\ݒ*��]�K�ބ�q���#�*��i�D�7=Jȝ�|k�/�;b�>��^v6�s�_vf>�W�Q��˜�@ϩ�W3�E���]���`V��vr.����5&"�̠��W]V
�~і�aPѾ�y�Զd��i(�;�A*�Oߨ�+��[�苣��kW}k|i�b3��n""��߷ �1�s���/=��y91�#%X�B�H�Ґ$���`a~�U(�\��d���c����3>i�Ͽ��z��j�H����	�k�J	��k�H�����a[��jZd�!5��y�p|R�W,�c���2vїbP֣ bg]� @��N,ǚ�� �;�&_貺���%�iP5\��u'ta�$HzHp�f5�#-�������PN��S�G��T�
�_�E8y�9�D��-|�Iq4,Fxq��#_�s�u���c_�1
wM�&����ޗo��#L��َ�b�f`?�|Y)�W5P��S�	_��ΧY[���~|�H|�� �G�*c�K��K�&�A1�/?�Dj-�qlݮ>��]7��[�Y�!��С��N�m��T�E�S)	\��X���q�f7F(\ê�F�!�!��U�wì����{ �d}��Q�G����1v��l�zL#J��/��໛�I� ����j������s=ŎA�{(~�*c"�9e�r����D.^e��. ��:T��~@F	�ؿ
�Ɲ��ԝ��i��d�w��_�Ge0<�v�Qx~���a�Xf��@Q�Q���d(��T�\��z����OM���ZBE뱬��68ٙ`��i�.�K��6<'���Gf�ZCQ8���ES)ߺ	���Ճ����T���0!���]T�8���*>ؐ�V��bfo	.�J����j�S��S��"���./�\PԧB��L�.�Ujp({��9$6�^���wK�҉��-ݯ2�Ԝ`K�L��Z~N�Í�?���M��l���B���j߬��tDT���j��H�����8��9�"���}H"�]�{���몲Bر���=�� �h^d���3�|y��騽A�:��:`����}�H�'F��ߡ�b�A�Q����qZ���MZ)������/�0HB��hiF�5�����(�d��z�%(���£]j��B����N����(�9n���J��
��/]�B
�QLK�1���L�T�s7r�/�D�JǾYʇjr�b{�$�u7ٯ��3 .����$<L��&(��B)&p�clTL���ҩZ'�Y�H;��G�F&���H��FtK>�9���8J���d�̋%A�w�htk�<rf��wQ��)Bhɩ[{xr������Kӑ _+���"y��<:�(oVq����������2��[{�����^3��I�c�n
B�ۙc��\X��[n�m�cH�l����i5��� lL�h�g�&��a>�L��Asr&��vݺ��K���pZ�֣Kj����M���l���g�L&�GF����,�;��:M��m��)	�f�7ι{�7�q�9����II��t�_�\#K�ʺ傰C�)'Ν�O�������A��w�+0V�=9�ej_X��/f��|]����1�v�(�T�� 6�)��EDL����aA��,�Kk6<��kc@�=�y��`59�A�H�N�_#Q(�l���'�����ö��ޠ�mފ�D�O�.��zC�A��t�@��wH<�'���e�k3�ޒ����ဦ�d]xQ��U0>�؝���Ԡ�N��%�/�����~eN�r��h��V�ۭS�޸aB��EL��P��E���O�F�?W�N�]�z��ᩒ*���/�/�4P�۹-���c��}�)d�p
�k��f�R���;�U�a	/��6�>��g��X1E���+�K8�@J��W1�|���f�?sviET�%�F�ʛ	�K G�[
H� W�V"$INg��}'� ������,���G�Q��8��^U��<�'苮~���������ļ���F�",Xσ��<��1A��f��/�� ��Č/�����.ޯm$ya�S'���F{;ɷ�U��vQļ&�jȰ2�顩��PDC�T���	q��q���'��.�|[�Q�26vJ�h}KN~'�/W�gsvk%?���t8�S8��@80����C����_��u�!��gTw��Ʊ�����W�`C;�}�'QTX�nb՚ O�H��zV$[C{	����QO.x6P>�}��Xf�5ϨJ�k�@�4�11����U�Mh[����_d�r���]�1�}3a���������z�ްO�J��=0)P�',��2ͬ貕����
K����b���Iq��*�7�X�Is��EZg�z���W��ޒS":�����"��ΠwSؾ�ػb�H��A���"�a ��#:&�R��{5��j�x����GS�����H��QZ����mc��:`�~c����Y^�^��+^X�![�HD��� ����OȐQ2�n轎�]M-b#U �XrR�o'�����!`�y+�d���I�����,�-�K�	6���c�br�eK���Ui@K�����h�qL�U��]p	�Ϋ����X5���Ԛ��Nm��!ա<�FO�%
/i�os��G&NN@���Opi1�=��o��e%c�~-1�c��K���ob&k�+On�V8$vH�)��er��m�������-E0��ūA��M������J�1W/��K����!��I��J�� g�/�Q�R��m�#o��43��x�KttA�K`M��C�3�w��m� Xb�mv^	��*��	��{��%l|V45c�-
,��2OQ�O�Z{S�,�����4�4����_����[m��S���f�B߁��#�Ԙ�R�}I��l�T�c�./Uct糸�7Ϳ��ǇWI�������v+.���[��5���qN@_Ջm��?���S�P��@�X29����a�o	x�ɰH-z)A�6�2��8��K��OLnq��%U�J&V��y�K����e���}�<�/'?$Ƴ#E*���6$n�<\��|��z�[����� �������O��9iXs?u���O��{�;��}p��;JK�y-�8��χ�5Rc/$
gn��d���i8�m� Nl�)'��&6�g�}���NB�u��}�"R^:��,6��,��G�� �)�o��'�-,��E|�e�-󦟆�}I���s5�GH=��N��,F<�[�R����=�`�� �6y0Va> ���fp�oԚƙ�Ⴟ��%���E.CF����{ �����0���= �1������Z�D���o��1I�h�#߻������eQhrjG^�O0U�BL~�
�{�%ؿإ🝘�熥��=�H�|� ���|[�n^(��]�OU	��bR_~�>z��濵�ʷ��;ϥB*���j,�3����:�Jp�G0�������p8wr�^�eU8y�Z-��K�4u��Ƚ%���%�dt��0��}�8���0���֙{:�/�9�^�9��)�t�*>K&~$9.p���5����#��^���:/?[��O��,�H��{!Y�ҋ-�[�h<���=��,�9�c/��'��z<�c�Hy�����2L��!~B����ixS9kY���1l~��E� ���/�K��_r��LN �PR�K����7ٰ*Sg����$E�S���\�Չ�^p/.��,�����w���75��ˬ���ݏ���:}A��'m:,�A�
�t�ݻk�W?j��A�S32��n�SK,i�(z*e`l� ��<�h������r���t�%s�g&(1�Q��[Hi��7H��)���D>֎���P �(�^}�1�_*�<v#���8E
>oX>>*�,��� �g)x���8-��ZZL�v �(f�#[Lf�Sע򱲃���^�u"'{,a�k��O������gM�x�ld��U�ThK�Ġԡ#�dP~^���,m����4I
3	����ۊ�X<�K���}����=�F-jis�0)Xj�A�g��MRz�Qrm��?���T�� \b55���Y3'!=˦I�q�,�T��t3.j@h�^�KgSQ����=�Pes����%\rh3.^��#����Y��TY:�(�{���yo�jМ[�����ϋ$zߞ�?VS��H�K�E�)��nY`��_�蜭.N�(%��-����8�2��g�C}N%q�{���o+��Ì�:F��a7*P�4� j����K�8ɏ�l(txreq�-��Ik���F��3��~�6�ڃп�&�qdQ��������y��R�Q5���TO|�.J�������HJ<���"f�r�/좬��Z+�t�mK��;�	0��g�����-xW��R z���l�cv/���k��d���$�R6��E�#�����u$C�</����rV�W?jI���(Z�o�xs*��-j��(��\�:��>��Q[D��1�$&8i@��xj�far�'ؕ�o�Q�y�wR���~��ʭ��(Jz�/ȅ�=���#�x���q����Eri��\������0��J�Q�x���ⲏ4v���D�m��O<T�s��2��10�[^ˮ�j����t�d!M����_SQFrEҶ��+�J�]�=�Ӳ*|h��5���@<;L\U���ptY�K��F�<p�c��B�P�����2(����F;���#��Tٻ�#,�B}̪�Ўr�_��~�G"�r����������xvԭ��@�Hmr\��BY��iT[�M�5�����dA�ڊ⺢�<ӌa�>���Q�����T�#Fy�ߘ"2�^󒏐�8.����$�q��B�(ff�Tl���v��.�;�D��f���G��YC�{YlS�.�8��U| ���4�{��1��7J������4�y�+5h�#�&j��OetĶ��am����d��L��'���ՙ1�9���,y󟧡��%(;�P���?|����)�l*����?9�Y�a������d-
��iix�&�������F�3�]Y�M~�1Ռe�3 E�<('�4���-B)آ$�J�����^���Ӏ$�'5bH��X�o��r$Z�H4���}'� 5	��m5�51��`���Z��&�x��)�75^��eSh<܎��H^�o�P�%H�-��?7�|���Uҥ��Ɍ�@/�n�w�'l���i�w��]p��1�)_�_"���ʷ�9<5IM�]˭��H�uwI7� ���7r�Cv�t��>�����4�U?�<�)Mc��9b�5�����m�����Xt��X�L[�؁���Z�*��˻��@}��sX_��KҤ�}J2)�\i~/�>i�δ�MlAtϗ>���.���-����1<���R�5����X���H�MB&��J��؈�Gy��� *�K~)���@�F�2D��������E�t!���ܫ�}��)��s�ZV���L��χ�ȖΤz�$~Ш�j�Ą��ߟ#���!�(��-�WI�z�\���?�I�iy����}&��C��W�3��X�����| �ox\�=}�L�4���]$0L���A
6����.��r��^O_����5�k+�͢�m���Mլe�t/��H1�_ 5%�������z	D�f�8�{(#؀��g�[vx�)�SM@�d����兹�"�n����{�؈cҴ �X�DU�y��x~ҾVQwp>^ծ���1���Ϧ�.V8���W�c����@�F��|�H4w��%���$�Enɉ(_�3ı#�~4����;�W�T����!���*u�#�� c��Z���Ѥ<@3�P.�H�.B�z'WS'����U.]�5]�����>����Q=8�ȵΨ����e��>��Q��#���Ii��|�m�ϫ��|Y?�W!�0�b��}�VW`�Ʉ��M�$�ُ~�]Ľ�wv�%�*+!��?�˶��it-u���)�?}�k��U��K�a��@Z"=/(l-u����Z7�y�|p4?���:` A�ȧ�����<S�>}M��Ƈd�x$� �(��`�j|�L�7�j
o	wTO��a#�+{ �
q�M���ʟ�0��X�#�@�.K��HS�ջ���x� �y��&	r�g�eKu0���eJ�a�����̆������d778$���u�5=��^����� �0����ݘT�8K�.Q�'�3�;���o��i���$6@E�<��T�p���{�o���"�hG���,��?�ݸU^?�� ����`Ȧa�b��1e	0�S������YmEeft�P�m��o�X�}�V�(��s�_�붂�F�[��2�(�.˥�!��@E��:�^�Y���_�sZT�)�d��v�k]�R;�\�3�f�����F5;��z1n�
�A3���/�b0��$�p��N����43��	^Z"\0 I7#c����cȯЧF6�R6�ȳ��nDd�4,p������A�Ÿm�^{(���&(l�]��$��
ik�����:X�^�;�Ϟ�r�~����u����C��*T��5�f�N:������������@3}�,���i�^f0�NR�ȵt<��q}�o�l�Gә���	mY��#��ׁT�jܟ\�� +���g�{�Z���N�������T1�6��x3�"iQ��!w	3Hz�>B�;h%�-��<	/��z�b��d��7�J�H���j����m�A�����b |w�OO�U������A���(�v�YϘ&����b�K�SZ����ϼ@>�-sv�-��j��$�����P�'#U0���<\O�؎����pH��q�eJ��(Eɘ�|U[?�kQY���3���%��E�z�Y�`�-lLߌ!,Q�ߨqQ��'X�u�~�z��}�&D~z�����΁񆗭v�(*����8�:���=H:�p"��� ��+�a��k+�@#���Qv��۟n�]#��$ئ	����P]OU4�ƿ�k8���ebY��3�9����5�	�01I�������D�4�~�!��aT5;-��f��%�A�ָX�g����q�Kkܗ���3�x��f�RR,�Fm ����LIfW�ܔQ���b�׎�&��h�M��/����K�16�t�Jy��G�6���P�ZK'D!½��EX������\�F��<��}A�i��h{U�	�����.��wЊ[�cX`H*�#�S���ᓢ���cmS��L�4e���!��?�%͋��rB���$��C�������'/X�������,��x  B���i>�h�iҘ����#�.�.���mDuEa�� ��.�4rW�&��v�{��I$��-0�_���t�v)�U�ϴ�۷� i� pYh�e�(�2���×����w�h�"����A�����F}�y-�wb_��)�M/p�xg�%4�K�z�Q	���]Z�^E �|� !���-}ƻ���*ߺ۬�������f"�Fb�V"�V�X�E��z	����v�c�$�����_���X��;����/�U��Ù�v8:~��ܜJ����9Sa�q�/����C�E"0����2���ā�[OK&W�����R��}�̊�3�:t��|c+_�'�+���'P��z��A>Nj\�"�-��*EP��Q��ʱ󥴽���
��7�!,x
n	�9�b�aLL�̉��7���7�1q��i.iؼ�Hhf6�1���z����O�����o��>�1Ǝ��=�O�ԡ����또�dL��7��968#\p%�.3N[����*{��b����ݪ����4��#�)��~��=�Z��������(|IºQ���y.Xp����[����)�O,*���/�������3���!lV�)�+�(I﷉>Zu	��]�g����&��|.{�ڲ���գ4/���Y�+KB9�k�NZU�Θ3ǲ�.6ߏ���E�w1 3�,�Są7G$���xt��]K�Y�ߐ~��f�,���m��Vj}�Ҏ��A7��'����;}5��Ծ{��ҡg�3_�D�=�cץV۸eW�\��}���91�'��N� B�oZ��B���VsF(���Jݧ��L�p�v�Vl�<�U&=(T�N�{[��fJ뼞@���݌:`	�Ϳ\�����q��jej��m��T�c߃z�$�!�)�^��6�� ԒRօ���$�U0�`ۮ����K�����rX��R�wvp��`|�j�3�4�8�y��篦,Ğ�F2���S+��_��-�[�(�V�E���|���V��.3��O���َ��n���5�����O��'bo/W�)#=;s���I?����.4�'aa`+΄��޿bݴX�#�������a�g��,�����Mڪh�l�����y)/8(T�E�=lǨ���j̙����8M}�����^�k����yq�=c�N����Z2�T�&�+n�6��r��=Mvg�_8Q1�@��c �Jf���Ӟ`K���S�7�!�(�ey��U˻G"A�F�Zb����8N���N���I�u_,U{�2g���-"��d�����h.��D��,���Ȭy���G\j�C�N�A�]�O�l���Y�8mn��q�$7��qm�����	@�6�����͇�6邢E��lx�>T�#1����&Yl�x��R��8��o��댋�~�#n3��K�Q�q�B���� ?�A�Ck�![��n�{��aB)1����ث��/hFOs
{wS�A$&T(�yO|a�����f\ԗׄH��ۀ��+e��#����#X�C+�b!t�
�99D]6�׏��
���彤������ݤA1��:����7�e$M��B��>��]�5��(l�p���T�N-�����`�ϕ*ygI{��@�,K��
6�Bt�%�" 5�X�&����f`l2��Kwb��/}��L����|PUU#	N�0f�w�Hj�Y�8r�>���ؤ��d2�=\������1��U�),L
��D)~7��3���D�x�5��	JF�P0�Lq�i�r�Be���^G��}kw�����Fl�x4`\v�#��,ab�PY�0��G�@�?\���j��u`Z
ò��S���Ќ;�>g�]춺o��qwhQT*��,��m(4Fā�bV�u�m6l�C~A�C�}��}7��uw�������?oD[���V�͐<��s�}��i�<򬉱���Xi�}Y;�?�0ۄҟʟ7c۰M��+�٫�*Ȁ%�>F��#�JZQ@}�T
HJ�:I^�?�[�+k�/Ŵ�o�c@_��&��K(�DJ;'��3�Gx�
�IP�(�?'���죙������!*
./Wy�͓��b�<Ut���\xz�i4E2�gcX���`#��T��6[�ӳ�aO�o������o��dR�Ϣ���د��t�6�z�*�a��LY�������3��)7'����gl2a:��˥��*�{���-�q�l�z��a���vvI�Y=ߢ!w�9Ї����{V��R��2x<y%�,#y.cв .L��,����Lr��xB��e����.�7���\�#b���_O��T
r-�)u�FB0[l\��P�P"M�L}��3�W�A2�}��*��.��"�j;�rs�oq~OALL����z���o���?�$V#�l!��pBK��G	4�.�\W��j���܂�9�nH]M>R�8�BL�*��<���bٖ�#��5�A�;�'	>]���9��T��#3x;�յALƅ��-��	}��U��r�&����2x���5MW'i?`"�i��Y 6�H8���PJV�T1�RN����ǭ�w�X���� ђH0�qZ�f�	Y��>����h����kᮿ��=z�3�� R���ϣ��ו�{�,9~.�E#a���eo�:��ڱ�g��:5*4��ف
��6����F6�kv���<��Jl9�hf;�Ԅ�;�zt�yB��YА�~]�"�d��6L�S��ߦ]m�{@�ݫ��u8�u���vD�(�LiG�f����؀N�y���ۼ/Xb����A�J ��{��R{�w.շF48	i�Cћ�����$-�հ9�>������"�����.�&��1�(F����R6:R���ʕ�Qw0*�!&��fn�@|9���B�CbZq��P�r5^�
��Oـ$�H���2Hl����������-2���9J� ��rd����EB�~J�vQ��R`��-ծek��}>���b�vї�[{-J;�#4��c�����c���
�F�36�	�/�0r�(�W���_"G?\HW�3�G�S�B�+�ES��vc��@i$�~e���?�����JS���Rx����Q��x�jW�[s�����_m4g�M~�|j�Ǝm�HƳ."��i��9?mQ�����ݍcJ�5�A|��{ֳ�_�ɻ�>j�h�|;1���m{�M,W?Qfnr�Wj��a0H�Sq�(Ի��ˏ�7b9����Fug��,�(�D�4�-$�o9���w��q"p����@��=Q� ڛ����n��y:���8]��׾�Ȟ��Mb\��60�{鲤iO��}�D��Ѧ�>��s�I����C9����>6#��,E5�ߵ[��9&��z���D��Db��<~}�w��s������f	� �;o0��l�
��L_�t���4(�\k�;H�ۧr�f}'Y��3��$�W>��v��R��z�oJ�z]�Y�@�:+2s{�K��K�øٸQ��Y�����Z�������5+F�,xs#�ד|�v���҇(�I�ă�D��G��2��Y�o��|��ԟ
�� ���i�I@��)Z�^�{�J����]�IQ��Y�3��'&՚h�X�#�}[h���7�i�[͏�s��'oCQsV����x�Jrp�����5�:��a`>R�O�2���w�<u�3}"�q�a� >F�+���K�?P:"�%���HR�����ƭ�P&5�'��~��Î��@r0���mx��"/g��)�k�N�~.���g��]�����}��sŖ��g���	6��͹k��IB�yޭb;o��v2W��6Z��hL��+{� 0�90cu�D�k��V����!H�n�2OgY��3GN@8����}'~�C�����.Z��s�ܸ�\���f�=��h�K�p�|����o��������HN�"&�#��n�&K�ǭ�;Y���t\Ԫ�rYMC�<](܈��u��:��}1� ���|2�����\�����$��y��ۯ2OC�?��{���� 8]O��2x\\Y�=X�o�c$���{�va��,�B�l�MHy��0eY.n|U�k�����H--&�eسD0�u�F���MQ�ڎ��lOzV}V���l�0=��I	㛶�Q\ک�(��_�_}U��gᮽ���E�W�hL_��.BGK�u<�J�k3��dT�3�7�W�~W\��F}�!z4����G����u�:^�߼���N��&���s5�y�%[�? �Т}�9��W�dDiuࡹXf��_=L�<�7��|B�ˣ�4ݧm������E��p�����C�VzE!&>��T�z��ݶ����Ǔ.����?�D��т7yVY]|�&W����P�&qI�e�%Ԅ(� M�'�E��	j�|��������Ox
�]��SĎ�=�-b�v{3Z�|��(.	�����K��+�����F��gz�$��Q'��0fW�'���	�qyV��柼ȷ�Z�}�M"��,&D�>���|����B�"�ݟ}���ݏ5A�U��Ǐ���f��^Aec�mj��Ai-}|�,���W�!Pe,Ί�j~�/G!����ʢ�|�Da/��	֪�7LJc9�@c��.9��҃����
6����۽J�.�:h���J>��v(���2b4dj�L�r������8Z0����D�<�P�g�ѧ��[*k;�l��4��.�B�i>�4����ɂ�J>�t_���~���������͚<s$_C�0�C�/�[�ʷ�7�t��s���Vj��������65�h�(|2?��8'UHyHH;�:fв掾|s {��z��ܿͦ��A�>���>�'f �g��L��RTo����9���c{Y�U�fB4p�?+q=e�e��I��Z`<*�V�-N�kA��bω�؆ў�G��1D˥�[�����kj���w�Rt�._(	xXtc�E:�,"G'bD��nC��C�-r�.���Aq_[�=jOh�9{�#��i�hm��Pu[�����?c*����-\ty^c`�[c���25�eKd��3��?��ӂ"����?� 	��<������M��^t�xJ8S[(=O�+ٮ}W��}�'�/\�sh0cB��l9�R;�-��o�֮�����)N���RV0�$]F�7]dKpH(����yĕ>3-N�D)�A�wz�I6��#���Q��]Ֆ�@��L�+g����i=� �)�`�+,Ӏ���~bq_�tԂ���t�I`��O#�V7���U�ށ��F}����w+��O�L�
������K��2Xg̶"z �Qɳ���ϋ��n�G�P6��&�C��!�J11��1��C��"��a� �6�4���U$��Xd��-YI=�2���T����˨�=�W�qΚ�����&e��e���taS�9�)�*����:G��-�~�v�<-́����d�Y��mɥXZ�vk�J��u����L�uA�������O���Iu��gFF��q������
����a�ȕ���R�n��o���M��'��6>��7�3'�%a�jS��B��{:W
Z~��yV������Z�ZK�4΍���l2��$�TP��D��C��f_��"`?�l�*1a1g�G/��&����?�@��o����F��HCrs���W:!��HG|@QN�ނՆ�(B����u�R�C�㷼y��?�	���!��?�aא?��j�'�Z���`:V�dטw��B�V��&�����OoRo��l�h���&6p6KnG�B�h��]a���4A7���<~{��Oʋ�}��G$�e��!&f>��\��tXfE�dy�.4(�+te5��}	s���lID1�p�Ƭ@Q��rY�*N��O�i�yx�\7v����W�2�8J�"�i�1�6Q�?se�_���X�q�$�X��r��0�D���ѭ��#ߋ��#Hm��g�� �
ء����"G���@r�캾�`Buo��'�
汙��0P�(t�@N��1���Qr��d`p�Ɲc���B=)�+��vD$&c"��i�H��]�2����{��z�:��s��>t�.�#PS�������ĝD\�<��4�\�=Q�y+�EA<|���9Vt%7�(�������h�ŉ�P��r��~X�%]ٛ����̘ju���W8f�:}&p����}<��1?G����kF�)�}3ǵ˧�J��$��E,������>��:����,��Y�zv�R���!�Һ V=%���~_2ßm_����}�7��d�x�GB��j7/�|��c*\�h��e�I�qQ|��c�M1�R09���4�gB�~����n-�
-ЬE��8���.�	����c�ëdZ��c6�q�=ɗ���/��%!��P[|�37�b'Ih�3(���H�<�M�V�'h$�voR�k�,|=��>� �I�Z^c�"����&�0y���~���.I��:h�:�V=���wZ��$��]脎���`�Y��q\)}�h�����D�E���d(�6W��J�z�qӈӾ��55���W9�F���t��m��������H�.�ʲO�ɕ�ay��U�� x̵���6S��碈��QeK[j�C�:�"�J�uHK�*;�x�9_}�2
�8��^5�(:�
��GW7i��\����\<�b�:/�5Kz�M�D��\v����0������I2�Vѭ����cr�����٭v�ZH��wkz�mZ��8�c]��* �)��==J6ƥ�]D�������갔�7����H|�|g�;-ޥ�wu1���������e)��v{���,��FCE�;�;��!P��P�{֤��3<յ�ۭ�X�)����AI���TNN|4!���
��Q��-��L�t-�r:]n�	�	�̄�KI��:��1[�Gp�@Z�'���ظ��&�u
��y��b]Y��:�/�I�pU���q�#u� �Xf�4�0��\S�`���K:�����B*�L����w� y�6�C�&}3s�z?8R~r����� ~Ѫ/pv�O梛�����]ʙض���c�j;��ݕY��h+���O�,ٹZ1��!�_P[O��ɫc*�W�W":����ߧ��(�5��"J��%��1 Gڣ�D�i�.R�l�{����<�ɽ�d�b0g����'�ڴc�}�6���e� �����	Έ�ii!$~��S�=��� p�ƺ���]a\sj'H�x�f�P��re�.S�
7��ѧ�c���ڪ���~��l6�^Ԍ/�;����YN�҅��vj��[¯i{y���8@o.��7=�xץÂ�|�x������ba?
����X��%����:�۟OO�V�Ģn+��#�.{�n�8�(j��q�7d0B�Ex�q{?WLd�'Ϛ���.[����xr�:�D��C&E9r�+r��v!x���ͲE�ؽ �%'����|P�a��f�y�,eJ�Ӫ�7�.��tƑgu���	���@�?M0�`�Ê�ND��S�w�m��5��da�T���B��H����%�OS���]0㯐2͇��&�����h�I�ku_9 ��"�T8��
o	?����J��@�~U��6����$f����~�^�"3��uZ���d5���/����=��E�fc�G���ӝ��;�)�Z��"C�{4H4�j�K���k@�����G�<��"�<5����n�x4ҝ�S���g��N^�xr���Nӟ�C��}<v��k���i�CŐc�n�fxC�њYB� {�M#<B����ە���u�<����[����>׈�e�C��G�<��)3hO|�w�����Y	�8׾9r�I_��YO�Y=N���F�f���j�C��1胾�vR�t���f�� ���&�1|��.���6%l4Q�!k%��,�r�bvd�l.K�g��?>�U�i�c�s��._�ȩ�z��t��᫓#�^����z��+��G#�6���EΊ�0�7�4���~7���`�q&�?Qđ���%���.��E=��5r$�WCS�]TT���l4b��{�)E�9�3���蜛�+"�ӣ�]��_��+���s�z��w����+�L�s�9�|�7�@vZ��~�� w�rv0X�ÿ�������RA��z�0�!�WG����֡o[ڽ�����Q�~�&��=�E1ԙ�&$p������F4����GU*J��3o5a�S��7Q[&�l����a��I�'�[��ʤ۴��^��	���j,l�3�]��`�Zo�~��y��ͼlyD�3i7*2�����W.�z	��l�I۵焖�����m�q�*��M ��V!���F�C���ڠV��힁����F7!r�-T{]OuAf�jx�����T��v�7�:GWPf�ͯ�~N�H���g:�?�W��,j?��ԅ_��|9ن�Y$�ɇLϚ7ʵ}~h���4s���Pg����'h��b�Z��$���+���-w��̯Mx6>���0�rX�&O�^���DN�Y�V����h<��v::���/�$�!�o1{�;�]m�`�m�k3;�,��~ё���˄/��E�kNI�޷�	^��#��#�כ=9.;�}�R����i XK��0 &G;���#��#{!�h�Xu�.��>�l�lSEq_�n��Xl>�u<�76;B�H+��Vq����͕jq�"Ci�DMHoh(��훐!foe�ը=l����+{��Z�Ȑ���h��y³�[�����7�:�f����ru/����#��7��6�"��8"��O5�h��dh;�u�ec�k���q��9J?��<�d�L�]m�����l��[p�io�4�uLMš8w������^���ݡ��X)��V�������˛|	��&;��s����d��6|�H?�<����K_nʝ#�������_������w��v:���4,8<&Ahu�X��vX��B�9K$�b& At���fJ|I��h�q��������R���UQ���`$��YȜ_�����ڏE��k�0v����O�Mq�ڊ_��O�`�(� ��&QtS2�@���tMXS��xϲ����H)�r�NY�����(��Ƽ-tֱ˲�b�n�p��Vy_+�N�n#������I�LJB7X��B4[�lĥ� �-��0�j,��J���|XG������D�b�7zܨQ^^fy�M��X
,�8�/�j���i֛֋�bM2�V;��UH炵X,�m6�q�.3@�N�����x�7���R�AE���� ��HC�h}i��a��h(���^��5`�K���2��E�uM���i���cݲ��@���:�i5�����'�lʴ�y�_]H�qq��Ì��YoֱT+Mp����S}A�!��%�`���TP8Y`ye��?Fۯ��(Z�-����]�F���+Q�:�Hەhw4��@V��+��H^z{י*]�O�|�����6DN<ߍ��w�&�Ɠ���~�Q���@�H\8�~�Yޠr�9%���	tW�{�����t+5�h���4��������ߑ��X\��J�_QO�������+|OA|��mѣ^:�x��%�0?�P������|�«��.��[棟����^���@�4	71�?r�zY9��f
�;�|�o9�z�j�9�v�5?��qC�(c�0hUs�QYy~8�����e�|��M1�ٵ�綏V�
��Z{�s��m��M����/~�K'+/�b<!+=i*�ۈ����b���f�&���J���:ϲ�嶧wԧ��x3!�`�I�(�0��q��u{h�V�L�.��1��a�9�K!ʐ�	����>�b��<�4p�Fƃ���Ej�[��L��j�i}I3Y^Zxp�W��vZ�f$:2�p��-ۍ$����M9b��߼�(z�|~�_P�`�9� ��fF�Y����}�¥�Dl��%_��׼��7��0\V��v+iQF��M�;q2S6�wu�H �ڹ4��'2eL���:J�Al��+L��(V���U[���R}��B�\}�n+p�)]u���!;�$o������x�(����=�`$8b�>�5��C�;^5[�m��4���ܻV�^D1/]R�4�z��Z��Hץ�3����I�����\�DJ�I�j*M��f
�����:��.���Pj{5*�U%`���ʦ�0�0g���x;b=��F����^:���C7�T�o�$�j���.t�'���g�q>�z_z^Ѡv��Ǿ�K�m<�H��!�
��V�5e}�s@0I����|E������Ӿ������(��i�+O�Y���Qc�X�y�������Ƙ,���\�̗�pM�g����"��BU�ڗ���O�氿	�j�{��n	NwI��E���5OJ�̵��:�c��K%cϊ8�f"y[x^/�`���`�o��N?�f���V�Zm��o,j$9�Sv2���v�K��ȄO��wa��2Tr�GB4}����7�ϵ�X�tb��;�����電�L�ۖ9�;]x}���ֱw9�C�?��7P+j�.�ZS�"�>���鄠ߘ8'J�)?_^���x+v�.�S�Y��#�$*�e�K5���g�q�B[`t>p���.Ƈq�s�p�-�Qm��(���EK�%8�r�Ma�;��|��(��&�d8�o���,�ۛƮ�?[�����b��Q���6����u߅34h�i1�3+���wG/����?�!�6R�}Q+�H'w�BM�$�>�6[5��6Ι��Q�[�Rk݇�8s��z�Ke�.�X�\rv?4���-t.���:n�3c��<����Uճ�Z��l�&
Zw����a�/`Z�OY�E���7/o0���^ܨ�%�����\�g3�ɾ�N/6�K���������R�.�[t�snE#nb�N�+>�͚�ǯZ��S�K�ͫ�<� ���9X���#D�ӷ̂����w6�۱`�I8��������>�Ѹ{F��`\�c/�Rz|��1_~ܴ�KFڡ���W�ޣ���u�ү ��%x_T6��cIx�P�ҷ�XΚ3����,�R_�k�a fB�҈��3��{��kJ��eӁO���Sr)�I���!�m��B���"�_��NKw�CBls����~��?��*IG�JA
�j�rrEp�]s�H��_w�2w�_�E&�1����e)r��^:e��ʀ��E�x�� *���+�LyZ��qyc�5�p~hަ(�����X9��۲��j$�c��V����)[��B'�5�f(ʛ�7*��Q=�3�w�j�s�p���:���@�����%�!M������,XM<����jxT�
iעC0��@0�щ
R��K�|���� V@zj�P��F�$y��P�"G��ܶ�0.��L������2�Y�k匜b�ʀ3Y�V�K�ֽGI~9}�3�|٣���k` ܬ�'g����@���Q�H�ٖ�4��/=ѹ�6����5 j��H7[��;�x�c�u�C���q����q(����<�2é���Pt1��T9���pfדۧV@���h0�z�k�ɔ4P~2�Կ�C��/�w.M���uP���4�0ڨ���?�yv/B�B�5Q3��c�<�"Щ�n�x6bw�	��:�ۡ��WF���dø�ʘn�HL��7_�_t-��~I�i�ބ�Tpe����A��Ñl���)A�1�������s���z�wuf����A�I�f��k��=
4�N9i2���n0��A�mA���e�p��&:v����ë��G��e�W*N���z�x�Q#y�O/
H?�"N���ԏ��4�,�-��fS1X��v.��m���1�l��JK교�0Vnâz	䯅�)�>��%�H fCW�ܑiV��<�N��կ%��?��xR&Đ����r����)F>��,�����ya�+	���|\p5�����(�N/a�"(����7��88���ЙFY�b���1�)]��`I��K��i�<�PjW��F�#�+�=��������&H�o�r*��K�' ��	�m��p&uru��2�a�g�r���L� ���͘/\�����E�H�x�y�ό�}^��XM�ʖmx.���� ����F�f-�j�C�|�C�{�{�����X���=\��Ֆؚ01�}�����1�aV�+�x�y�_|�vgWa�a��ڧ�Mʈ�i(��M�\�����ɘu͵�{��O(��po��"�~�CP����z����2�c��� ��,ݥCo��hHI*�~B�<�����x��L
v'���ӱ�S�%C@f��)���2�����c�
Bt��R��2R�=�=�N�j��`�\,v���9tBc�}uj1�m�#?&���������F�-�5.��U)P1�P �"�<i_��l�0]���+�R�U.KS4�}�n@4�W�o���#�[��`n�% ��?��M��$U��L�eA���/���*sg��x��&�T��p5F�f��*d��'�4R��������gr���?�&�=�@�ݏ�i�k���(��90f?q�u�7��a�YJe�k2tS+����ė0�pЬ0
�!8O�%n���]�u-T�&$����O>���(�����5�>?��~��o�ktD�D����?/A�� ���e}d�D�l>^�T����쬞T�dz������S��f=Y���O0|�t�W�jd�S�B��󳃜�V䎽�NI_5��O[�)�j����T��բ��	y�kO��Ԝ�.5Q�wb�������L���.��C�����R�����eoj|y5��[�΢+.y��N~�����k��υ`3s�S���#D)VU���4����*���ձc�1[{��2�:Τٍ��;����u��?x:�s�9�k�]���lY5M��M�-l������z��J��ĉ&K_t�/�9�p9������tKF�R�B3�5��$V��MS�8�p��8b�������>�K�	qE���/�W�%ݻy��ɗ�%#���A�}��^W
�ð:���;ܒ�N�l��J���S��KiZ�+��xU�R�nv��lQ�sph1����J���\���M�ʞ���*rݲ��;�aB����&��(q�T8��Z��E#/��񠦧�d�x��g��iE���Ng��I��v}����S�z�I+�N+gN|J!!	����w����b��(%��.�?(��3YK����q�C y����S\U�>G���	/�n$lO��Ũ���E+�<{p���b����������]iK��W��IWL҂��"ѷ,H4(��Fc��e������cI"�K��!Yf�y���=�'��:M�C",�y���o���gξ��!�cvJ��k\�{��O�$0B�r"�c/oQ�5k<�0p���իX��L�l{����s!o�F��s��5� 1�JAE�jϺ�m:�]���N&�x��D$줞�3-�8�o�Ֆ�!�-��$����f��J岝=����C��}k��L[UB~�o�IW��_,�����D|��d����4����v�y\��SU�S��}^�*�^܎A�͚x��s�%e���ONÚs�r.'��k-�}��U���`�ax��4���d0�-'�	gn���M��A�Gp�c���6f����˺O�����O_ٙ�l��Ё���0��=2G������sa���M:^+k����R!j�����ڧ�X��'Y��v����ɚo�����|�ЛJ�#��N�tG-�R��e@��Х\?��H�A�X���B}�d(��Р�s� gX��B�]�1^Y�[��o0$._���������0iR�^��q��~���f�/ӟ��9��۪�����2+^.���\nmnspWؙ�F�"sou/��_��a�$�I*An�C��_��\�Jw��^W�D��-�bYsN��]}�U�����#�)}����=��a�|^�[xX07�x�.Qey���x'���p��78�;9����n�����0�tu�ss�ʫ�N�E.�C���á�h�Z��E"�_�i}xR�j�D2���QzP�*�L�CPc�[n[A��ͫ|[?l����:9y12��cU���'_v�ք|��3�^%���,��O�4*3���Q����n��ª���,t�O�c��I��1M����~�:x]G��Xz���C����UU� ��m?�fLѧ�xƾq��V�	Yd���6u/y�R02�)����
�9i��/�+��
fD�)["��A���b�0�f�qւ�����a%^��g+�Kzo�l�Ʒ�0�lB��Πq�lK`�NVl��� �����J��X�E��6�.���HI�P��AzB=}���t�}k��ᓗ0���4=�?��/� n�����8aͩI��n�	K;G���{�Nu�-���[`��U�Ȉ>�{O�)iAv�֬M��#��:�gGAw=��7U1 Ra��S���xz↊X�7Q&@�S���NSbCo8�63�c�Pټ�����ؾ��4������k[�C֊�]�����5��)��<�k7n�,;��r�}�k��LaC�c.�Hd�5j��S��F�`u�k��yћ�����څe��f�׳�����q*�b������չ��bYU��P���z�k��y�ʡ������ȶ���MٷKB����
�j=�s?���-�vF����%�Kc�*�YK���Wq�{��}Ba��m�)DC
Xd��cG��_�҆�9n�t���<aw����+(��8�׷�B���~3	��s��¶��W�0[�P�mz��H�ÚI�����	?(1z�AG����7!8֪v���������[(V�@�1ֈ`�$�&Bz�6P�g��%�5k�S��dݪ2�v8ۂ��b�7��S�u^$v�#�(GP�Ǎ����_!�`��<�.*T����)$���z����'���b�S#�僗2������4pȢP˧l_��&�b �	c��~�T�.c��-�7^o:���"�F��Fv��:�Q_/�q9W���8+jӝ[v��J�1_��ˁ�|�al�ZV���Fæ<f��]�M����\��?��skǬÏH\p�xQ���r1y&�9��_z�E�S���RX��� �['��ڬpk�/�pY��l�B���I����={�A�Z���5�}�;Q9C-]G)��Y��(	�Ԉ���}<�0�߻�B�!���j�	&��Ҍ�m��j�(o,��2ʴ��}�T�UuW��^x���Q�v��#c�Ұ���#�&y�]v�<y�ċ=(pN�$���QX�ꯖ��[��}�D�(x�g��ԋ�h�N����v�4�L����.�_����C�N�?�;���xlNd����­���O2Z��,~�Ȑ,��E,�ۘ͌+�Ho�g&�f:�&�!��bv���]V��K�R��j5wc�c����m�M���k��!�q<.i���2�k��GWM�Yڷ
?��Jsa㍥��R�5��Q��Pa���뎣�H�� BZ�����FE���Z������Z�V��?g��yR�A���Vp��2L�ESZ�fB�'�։��2�4�c�4�&�Q����vi
��o�E<!��o���G���;�J
ڄR6��?mV^
�"��l�jpg+�k`Yf�S� (A����Y)��{����jh���"5W`a����T}0#K,`ɇ��s=B�& |1~���l>�c�	��E$� ���jQ���g��
H��@�����,���n�]��_T/��[����y�\o�P�qp"oV���_p����:�Gg��eUQAv�0^��i�S)����a�%/�8�\w�Y6h,���ֳ��cՐj��u����Lo��_~|���^��y����6���屷����`ts�gc0r=pa�a6���]�@�у�<<1<:��n�s}����P�K,@�>lsa�J�~� �4�|縟L�!�S��z�J�������eh;�0��Xе
N:�u�8}T>i��z�7�k�~��o� ���[sw;�MT�����=���%�ք�/�tFK�������(nٕ}��>�`�N�4�b-�t�A�霼�	��#�&U�B�B)�K��lp�Z&�pG��3��ZKpѥe��B'G*r#�}�Oy�~Ғ��B�e��&��d�l�yˬ��O�خ��ܭ�gE��c�.��>f�0f+Ek��I<K����l����a$���#0v��gJ�7�Ç\�Jg�Go�M�ի ���6;�t�lؤ�_2���>}��s����c0��7�s
Q���S���~�<��A��H������~�����_ t[��[�U6����t}���D������qV침��/2��+Zt�5�&�S�=MD�M\?e��?ON+��R��5�U����%��h9�}.�q��3ǀm7��f��^��:��T=փ��L)t���#?�(F�(�Y��|2x]G�CO_˓E�B!rw����p�����M���ubhW����S�|b3K =$G���y�p���+�ZR	���X18P@'�{�}����O*� �	n�5��5�T�0
'�i����m����M����np�c��& ��{p�//9�n�$�� G|�4��V���}�"
u51��(�yR��+lȭi���� �z���ʃ�޳�~�I�E�h.�^^)��ز598ط��P#�m��/@.֪�����H	�6����9��s�}�܀����'𓜰i6�S�I�'�<��i�K:�؏'�/�]��7�����p�j$�� L�����<��KM��	s�U�<�0̓A>g�f�*#� �騘�b��G�0����"o�a�䍗���ӟ���^�@<����D�jʖ+O��e��:�2�3ј]��'����Ϙ�έ��]mb㐰)��F��<��E�kZ��>���l�=��K�]1h��o�[�!��8��pqC(:m����
Z��S��C L�=%�f3�O�*���%̷3KfM���Q?�ja��pb֌҂�3��7`�
қ;�\	= ���w�#�>
�����zq���\i_t��lqy^n=ʭ�eu�<���l"�1�ǜU��/,[�w�����u�F�P.-�QtK��-�y�7�HR�����rO-ʜz
�C\���w��n�/��T��KS�M.vqX�]㎱��7����k��������
|���LM5k��qQ����0ܽ��/m��/��f���&�|݇0 �Nf]���vQoN?�쭒�>�d��nk?t��H��Ǽy6Y��CW�W�����W���Tcp�L��=�<W*�Ԩ���>���:�G?Ԗ�8Q�O��^ӏ�|R���_��W	'���K����#�u|���b�+��֕�wEqy�����A�`R/��wy��2����4s�Y���,�ދX�8TH�R��ZP4��S�֜�Mw
3Z�B����/�A
�&�>�5�<y��f���y	S���@y���L5�����L��l��8+&���o�T�������Mx}$i���`���4!J�YP�Z{���gY��7*su+����-�{y�: ��BI!�dιzy���}b��h<q���j�ʾ"�Y��$�N�<��M7��bU��'�e�dLN/4#��8CL�C�j��ZU�����-����`�\��I��A�����ˈ���?ü�� 7"�{���[�)eG
.��X����?6wVĔ��/Mț���$�����<ɫ��S�u�.V��S�� �>Z�Y���5�Xٹ�tn,�״�]%�TpCdRE����ܸ2���D%*�a��G��� AM�ZG�z�H�Cums�{BD�����OP�?��Q@-=��mR���{��~x�!]�����G�K� �<��x�o?�(f�-��$2�-�o���&=VF�'�#�Q0�m_>ϐ�z�#2�%T�4S��𡕃(PЉˢ����JL�WG�cc���C����"/����8u9�zC}.K[�=�*5��?e{��؄��^������掱a�q�X�T��Db��>U��#�z�f���הG��笤/�<��|��sFj��4a=�[ ��o�]��x��2�����%���jυ�d�G��Ӣ���������wa�d��=�H;_%�Z,f*���<��<�M1P���>���RI󻻝8Ę�;բ���wP�A���ӫ���?(���VEO���c�ld}���(�y���[��t�W0�,V
"��Ţ'x|�AT%�'a�:��(�[n2%�N�7��"��JvR(	�~��,/�)��=��Զ��צ��׿��t�~��
_���gI�m������b��q���gPf�G�=I+��TX����NM���\���̚.|��~T�����, ȥ����^�Y���iKSz�T��$���Z8�zP���}"D���'Cd�@��]�����Ֆ�'���?]N���Y��?g�����<��#�޷損>�4��X¢.�*��Ŀ1�~{o}R����ูE>��L�e9�k^��9�]�S��v˃AꇆB�{�w��H"�5B��r�o�=�,M;p���sHT`Y^֑��}'R>SR�]�]5�u?��Qd@Zbi��ن���t �S�]Zι�%���6�Ԡ�t	��j��t*��Ĝ�.i�]������4��b��[U3���0A�h��8 ��Y�
��݌��v@��������4�򾆥�e�_���_~6���(+��wH���hd%�]p�b��yS��r���Ɉϙ��D�jӴ�Z6/w��(����S|��vo���j�,o�Z#�5`{����<�N�29S�V�#
i}_�E�Bp���;��Gֶ*�tî)�A�̤��p�{j�$-��7�Yi�/�uc2vG��Wpك���h����*��BC��
;B�� x��y��3�G�BI��rQ��:q���+�<�)�$k�9R��	 �\�MC��$!�c!W�b����'�`dW�ċ�^������O̧�[�ە��A�����.I�U���IS������B�RF����W�l/8��!��?�-1Mg]�(�,�F�t�*���(�,�<=�{����l	~�S�tݹ�	��I��^�=��yk�`E\:�QZ��+\�UnE��;̍���p�Gc��u�rQ� '�i�Hw�4(I�gɖ`�Y0�]���c���?������C��'��&l^�g�6r����
V9�cA�Ka��9䠺����6ј���r�^����L�`��]>]�Ĥqi���ul�{Խ�d��=yի��6j�+��;��[ ��X�\��B�p:7��5�T+69��/����Q���
�N��Bu�0���g�1ڱ~v[	<-<wB�b^���y�:xR|,�w�ԣ��w�M�U����L��ցò����"��i�^o/�c�h{�38�~�8�ir-;��H8y�\2d�����Ie�`��wB2f�<���9�(�ؑ�,������� ��pnLH�"e���7�J̩�u������`1r���s��>w�������K�Xٍ��r�땠�Q(�\Ƞ02��w��67K�N��e<��FY�E�*
�;����w�8����z����0��g��>pUyf�Vj��l�|Y�'��0_�>���dR�&[��(��Ix�7_{��z�evAyb� �&Vl<���y�?`:+^u��� �gn��;�}w��e�[M������x�fkg�}hn���9�Vn��Z8�� ;��l�4���=��ue��tv�<_���(7�Wlu�P�e]��s��C��J�m��>v�r'��!��g�]4R��ƝO��V�g8�[��H��Q�}ڦ~k���O���2[	/X�a)��i-��.=�ɛ�Oc�y<РW���fH�m�&^��B� y�Ky��~%0���L#�"���9}�4��8`ۡ�~���`��v�C�����#>�*���1[���l��E��Qp�Ӿ8K+��|g����
�݋c�����y���ðA�kPS�Nן����Hk>��M�̊R�&5a�q�u8�m?s�B��2p����>�o4��<wĴ�y�X� He9��~�j=%*C��o�>�^��.t�]$���ۛ�6ؗ_���}R4.�5Il� �=1�k�,�d:���%�WO�~�o�3s��o�m��ðZ�Z|�����!�8�hFmj�-�,�_B�
��|j$�B����7�1�
j�&�#�ˈ6���(xۂ5�;�ɓ&f�i�8_j(�;����O:EE���~N�!��AnO	�s(W1�'.������<zW�O!6��򻁿Y��#�UUk^��uX�8�
�7'DU^0�޻F��_��j��ՠ>vݮ	�~��*����7��Sv׳T�_RUu�,�j��n):�(S�o�N"���+�w�/i�]<��U�6�p`���+>Z�HK��7�E�%KgXɣ�	?b��N��˯o
�^���[�r�cbJ��ht&�,&Xz�wğ7Q50\X-A��/���*�wg���}�Ĝ��Ɋ�[;t��D�&�Jٙq�SM��U��k|���1�ɏ����Z�
=�S~%Q\Z��V�A�$x��7u14�6�?�\L���hH�]�(K�F��E� ��k�.Q��N���NT�����:��X�xB��z>c�A�K�����TtA+���X�!��S���ax�Y�y�뽘�͆oL]��F��޳�ʅ�/H3.m�����(�#[Z]x<�n��p�g�63	�L���H�r��^���'�k���@�,�m	.�&��'��B�q���X��������+�{���盢���;��6b��͵E~��l%���_�7��A�փ�����5���B���:�[��e�u�H�(M��(�����)C�C���і����Jq�M�/�/#���o���?��/�s�����\z0�>6�],��\�)B'?߳�4��ҺԽ	HA
�yZ8��;}cO0[r��F���Z	��5�H6aS^R�y�����fRh%h�,ss�N7=5���|�v�A�ԭ[��l�OY���.���p>Y��P��%��7��i�σ(�,G�"Qz8ݮ��d&_t��Cֽ�hE���CM��Ü��9P6�u~�c�UD>2�њ��U]�L��Ɋl}�5J��-+��o`��_�����\A���9�ܫ��\��xU�+SW���K.��[c;߉�]<&�Tb����'������~p��)���a>)�z��I`�u[أ0K ����)M�(�t��1��}�I���a��s�gt\�� �+� 
N�ԁ�=�s!E����긫���<_A<=u�,�,�7�%��*Ge��(��!f�Sb0�i(�~b�X�~���Y�J�����q����z�)>��w�q)����?6(���ނH���@�%+��U]�.�ddnR��]�t�[�	̧�Rj�� ��"����/>�xv��w"�r�
���`�3��b����j���١�������?z�������K�*�fc�9򏿜)�%,��,�#��W�e�"XB�e0��|���GLV��?��˃��\~H$�YQ���2�?j�_Z�"�L(�4��#��+xؕV�=M�3��'���_�%�Q6��jޕ���N�(�����Qr�"�m�N(��.#
֑c:Ґ��R)w����[��j`���^(��=�F��6٨/� ˻�_��#�[���XD�+m�נ��	����RB��BL�˓��ݸ_PgC~*�����Ap"6PW�Ɉ�:�	N�P��ԝrF&��n�yiIw^-���z�]f�HAbFIpMjE�9��A��Ϗ9���.�������o�=	D�uT��AR�ߒtų�LB�T�h�=P�ߎ�we�o��(� ���2j>Y���y@k�7��뽰��h;�;�bW�̚b���M�Wi ǰ����Y��� ���l�㴔b�y�B`�
zq�g�ƫ*b!�]����!���2��_�(��(Ȃ'����/����v��Y��&��@��\����ROj��+n쑆���c��&m��5�e�s�L	v�^�����9j�_���9���+��2����y/U�%�o������ͺ��n�v_�8�����T�%#C����0��Z��F<��?��\<\)���c@���`R�����N!Ǚ��!\k|�;�Z���p�bCK��8��Ђ"�@��?�qp��%�P�\}�>�D��'�}AAO	�>j2u%c�nGђk�x�� "�	\�!�������Dꝧ[���0�!�C�2��E&kj��ҖMԠ��|�t�p>?C�ы�In�),�K�*��h�ʴbh@m��@���� ƸO����i�O?��re �CQ�պ�r��{: ;�z�ul`���;oN%(�:��(�E �Xb���[��6�u���jz������#f�9�����n�}ˊx��ͱ���K�1��
_�q!ck�)A����%DcA^]8F�pQ.������ax%KY���iʪ�.�lJ-�ح��,K݈i��:kl��4O�ؤ��&3�����Tw���p��1� ��[�/�����}��Gp;�ČL�#��;⍪�X�|��Lx�] ��VU�eRh�}����ŧ�l�E�DHN�?ĎV���3nW>6b��c�*{�91�I�2�ë��M���u�:�S�i��(4<��Խ��Q�M^jW��������A����P}M5k�@�2��ƪdX�E˕L�{:��`�v�˵����K2t�3��-�e�ݯ�v��n�	�^���,����:Ro�O3���g��j��.i�DNu+�J�����i;�>l&^��"�$-4uv1�ૈ�>�t�>�%��['ˊ�/�d���d�PaD�gz���w�nF��7~T����DeQ��UE����}_+�~��p׋<��2EU,���UTi� z�Y����5�����}�C��Q'ۢ*�0��'��i9
��u|y�-D0��Lݠ�08J-4h�F�k�ِ��>���Ɩn�5����_�B�D�Vϻ��a���sN}�v�N���3/��д�� c�n%��A
�~��x|��\V��x����=�ބ�2�v{c����bI3��m�Ds"X���z�PC����>0Q_�����7Qf68i���S����TG9g_��_s���i�ǃ�Q��8��x�l��c@�7`���a���˜ݗ�/��s���P��,LnD�4pi��_�%[r��zę����IL���Y���:E{HG~��P���D��cOӷ��/tv���Ӧ�3#�Qf{2�_���ӱNk��#�~�y��~�*z
�w��w�Q��2�-��{�v8SW�
�>�s1���4�l���b��g�����K+�[��,��Z�4Ĥ��T������TI��B�52��*��J��j��m^\pOd*��t�!�w���(\���t ��+�~;GM��-ک:o��{��|�a<�rB ���hE�U(�q�0� brn2g��b�_e���}-�Q�\���Ub�w�n���������b��e��N���wy�����!��&��:?� ���l?Ġ��������V�@�c��Ȅ�T쵍?}xd�B��RK�3��垸G
�H\G%0�(���|����2#o��n�\�2�}�U�KX�%�&��7Yk7��9�`�!:�DgE��ڌ�J�w9H��_�%�Cj��=N��}6��E�Y��>�vV�p����\�e��͛\�e�q
nk����t���&�1Z �a��u ��g�D��cn���Tח����G��S�_��<���&w���"�oz��FBXI��3Ol� }BH��xw��i�J��?�#���$�y���=���h��3�l�	Û�62b����xD�y��)l�v' ę
Y�~��*S�,�GZ���(yΓ���l�c&!T笧�y��a�N �f���[�Dc�I�$.�*��6�GN�?0��۵��"��[qog=.���}q��"_��@;��"x�i �Q1�u�{�*]���E�ʔc��jw[d�#�:�}p�.�*�V�\R�����������iq� ��N����4�\l`��8�Ӥ�/6�3�7��<G�w�$uKuk-��R��I�U���bюl}�e>SB�ڸoo�oc<��m"c�����/�z ><l��W�߾wc���o۷�Z�'�n����[���y�Z���h|th�����	`P�}Z�����Ak��n}Z'S*��F����6�覮� �ߋ׎�e�Up�m��x�Xq��m-�k��"�?*�S�ګ�ζ����z�G�!�����G���W%B�����ː[	����'X{q$0�#mA�I/��8|�S/�������IA8- ;�Χ�4�aj�x`�1��=�`�h�;�Ӵ숊A'h_J��Rc��9��ԙF�I�"L_� �r#
�tH
��D[.��h�B*nI���������0YV
�t������]�]h6'�?����"z6�9�ȓ�=7Jp8�~Q��9x|�����dNx�D�x�=鈿������ݼ>Y��,f�rJ���tL�lI?�h����w�4��^ ���*!���h}G���2�z޽��/�/[�Z8�����*;�
��:V��ܲ�U�l��vj\_��辎Sf=[0H/�-N-�n���*�fj沺8у1�ʓD|�?�p.	��0�muM��A��%0!�⩑De�V���������Og~�D2�0�E67�,y/3'�"��Է�����nV����~������?0l�k9L��b!��
g��yu����� EOT!O>{��i�2�&2�I��PY
%Р�5?�Ş�&_�g1���z���D2�Dsᝠ��񓰢�c�t�V�z@6��Icih@-|-�,�Цl�
ǡ]ml6�.�/I�׃��f`r����U�B�8��-�l��F6����t#="'T"W3k�$q�����œ[�׋��s�vZ�I� ��RG1�x#pa��x�|��еszv.�Y�n�u@_�F�Z�� �0�����~?���f˳+�gI���
�Lי0�y"�J���w�R�{Y�0�lFY��P'1n@\n��a�6�p�Ŏ6N����&��=�؋7�'��J��x�s��v�ټ���F���Ǳ����0Mq�q+!�����I��`�TZ3�%�y��k�1'S�G�8���O�� n��Nr����[D�r���;q�vy��8��õJz����� ��k8�sV�'��7,��׾W�E����" -�HRJ�JK�t�4�=�R")�5�C)H���%�Đ���y��\�8��|�k���k����/��S���2{9�k��}'n"?�m��֟za쐆�Y��]�}r��p���e��I���4koV�"	u��,�`�C�Dh�M�\8}��K���V�N�� ��<,Y����,2�Z��y59>�4���e`���N;G�-Yރ�W�VZ��"ѱW��F���9;���Ц pT��G�ү�gs��h\����O� F~�0J,Γ�"�V[a}�![UI��,ֲ��f�1t*�+j&��=&cݳV�I�1�9%-3�	WeR���_hܰ_1A���.+wl�e�N[�]ɥ�dՔ-��Y�r��~�<��!'4;�Q?҆ȇD���������U�+� K}w���\�!�̮�-��9Ӝ���a�x�LP�iw��@7I�:��a�4ܤb�B�Ss�uF��_"!:^Z�R|�x�� �O}3X@wƫ"��_Y�m@Y��^N���!���ݽ���P��_z���� _�㣌��"U?a�.?�F�������2��)>��/bo&|���Kms&�יج���Z�YP��J;�qF�f�DM����Ėէ�l�@�pH�,ѫy-D�[SN�o����J͕R�Õ<���YJn��z��������ڈ�e���`�ϵ�n/��pmŏv�XG���M�*{+���	�y|F�vO/��DoA�IB5�Ob�JLM)���8��r����ɮ�����@��`[��Z�~e���XO���B���^�Y���ڻa�h�`��I���8���?��Kd�j �_O��Aj�d-�� ��rҲEri��� �y��O�Y�mo\���:g��3~A���L~��F^�Xњr���τkͷ�b��'�hh }�f�M����@����i�T��)��;���,�=�a�ۣ�#��V��Ia1��.��M��.�C�8T��\i3����8����f����f�Xu�~�s_���[�ƌ`���u���kr[K�z92�fo�e	XX�Hb9
'�O�.��?�͓_�k�##&>R�J��� $0�e3�Hp��K���缽k�+�@��w��eM��Y��9��e+�v�M�W⍬�̹!Tfsx4�hw�p�5M@�[�^��J���8;�o��8}���-�h�+�%�J�&��O6��%竃���;w�/�
�5e�m:y�/oAg[�f_űL�&��������������adݹ��\m-4�ݹ��AQ����da=��;޵~�uZ�S�ء�V�Eo�>�+��J~�G����kx4�.,�M����)B���˦6��j��O�~C\��2U�Ω	���p�&�) ��YhT��'⯸X�F9�+��ڃno�آ[Be�s������\7t
����k;�b(��]�e����e��f����=IF�m_PjL �l�5�����.i������l��_�~��$nKF
�@�]�I&F���OǄV����0��T�ѵ�z��®�;�����eb�M��� ������o��w47�태��H_B�}:A�#_>oU�_Ah��
�l�J�=�"8_j�p�/��|��U�:t[�M���U:�yڥ x��R�r_����y�}��筝�C�zlZ�s���&�γ��<��\�/IC���w�v�� �[�|�v��2��e���k<b#�z���YJ˕Ru�%ʪ���3� �?N�w�)�=��#�u,A���P`��U�ݏ�6M���yfa5�de���=�H���u,�9���o�tֺ�3�إ�uxЪ�������:.��$�~ǖ�{f)�����J�uo��Dj9�ɮRr�
;@��C ڍ�](f�Q�߯�+7�@[����#���~��ֿU� j��T}��O��ڈ~�$\�=�
0K0J�XQ��/ 2�Q�2uJK[�����íG�NlEE��n~_ ��j�s-k��E9��ۗ.�hU�c!?�k�5f��H�݀Z�<v�����{Qy��V}\JW6I<��Q@���qd�XR>/A�c,�u��?z�Hv�i~�kA`�Ȁ�`�5����Q=����U{���LC`e��BL����|�����>�-԰=�c$GK���	J�,	���:�/=�J�}Y����4K�;'�Crg��/��{Y)i��u����Ѝl�B���8����>��i�~��GS���Qďt��]�A�����|��^x���;����$���i>�tO�����$�h���̱��A���#F���
�j�d�$қu���-��,J{���4^����~���pW�_��	���r�l��Y�l�
���=I;���+k?~>"M��]s�������u�-`�D܀/Iοٴ�X�C��`�A�/s�WJar�16D<T��XdK�Qͭ���Z�Y���5�Ko�a�83��b�uB�Me{(N��K��٩�sXv����[s��$N�8�s��������R�������+7�ړjV�(��ڃ�g��?e�}%�\;�����ɑF6���hXh�Ƌ��D���p��a��5"c���fߵv��`�xG�ȩ~��<�����f�-���~^�?%� 4H߇/���b��?V(a}�>�<�v��9b��AW��s}�F�=9'���j)oO�;=��a�=MLˉy���	�R����&�Ӧ��`��0����.�������a�%���:���{�5����!���w�����޻b�b_��-Z:n������@|]�`"N
_��/�� Y�%Q���%ā���Q�D��*< Cφ�fg��ФvK�̵�M���bn�W;W�WQe�ؕ�?��jk�d����8�։�UAk�M���%�t���z>H�u�ܻ{������WӮJ 9��9,�C9�VBf����銝�q���?=r�L����8�}mĸ�%z(=ĝ[��f���t�Q٤�zD������L�^��3��!����.JINV����_P�I�!l,�(��G$|�W��-��!��+��ǖ�1]�û�uP����La��<b+"�ғ$8�*��>2vX#y4�K]�8���e�+��S�M=�Z���P_U���Tn�:7L��(q��a�l�zw曃wZ".�,.z<Q�N4�3bf�cfH�Y$N�,�1_�i���[�]
�h����imQ"i�l���'݁��=�b�8Lز�tXC{������.wI�gs��o�Rə�yAv?K�Al�xE��q�Zt8�"��w|�.��.���KU+}wD�f�=�9��]�?e����}�S�[�V-h�~��Y24y�!]����/�`J>#��z9�h��ǝ(c1�ޘK;�����UlC�!����Ў㾿�O�q��ݟ8��.���j�^{;�p��7_�9���q�Y6�f=�?)ތ�V��Œ8FH;�>�-��yy�����`����Xzr$tc�<r�ر6�%��s�&-�"�|�J��F�ӣ���j�J�T��������Y��N0�<t2�Vȥ^&DAw��}�.5Oh�,9Sy6��!̖by>��.�d��^X�O�}x?9���A�voQȞ��26�z��;�;�g��v��Jm�m��S"�J76�'�G��ױ���~��|�?�j*�~�;���]�����W��Bt_���w}������!�F���>g�@�[q�m�ʖ��e��'��Sx�R=�AJ�p���v�͡�ͅ��F��.���%��ʂ��JB�b�\w������n�m�xɚb3_���$��!��P����?��EO�,�tV�#K�w��_4M�G�}��>����翮�?�i�K�Z�y=� ������J��� �0�z���%��Ӭﱻ3�ڤ�Թ���a���I�'Y��j����?�5>��0�n�`�T�K=�aR i��A�=�u/���I��^�Q()aOҨ<�4{�Nd0q�V�nT"<&���k7�S��Cg}#�<#�iu����a���yߺ�>�r}����(B��򧋬�n�߽�m���-9��c��Vti	��H&�ͮ�X����6�}{7�<�@Y�t�O
�yݔ�_���Ҽvo����O�/��`;���tt�6&ۗ�����ըB������Mт�����Ј�ɝ�nm��_����+�:����^��5�`��GU��Wԝ�E�1&H?A�H�ɾ���r��	�$��YԽќ'"�wu�<��'\��m�-s�[Κ���q}g�(a�����A哟*adOܡ{ǻ��R_[�X��Mֿ�\B>9�|��-9�����3��t��/�S]���z����1KM`c��ȏ�PY������s��~�w�e�H��
�no�~�cҴ^e��)q�[�)��C7!�pM��GJ@C���t��$_S�'B��w�b������!]�Ǘ_y��+��wmj�T�Ζ��ΰ�����SAX��e��ߡc1�h!���z5�_+��Х�ݜ�%�M���<\P-nk��N"?�1y8ҩ�O�9\?�K�F����6z!���z����Þ\��I+�-)�������߯u���� ���[Ue0�󓂏��6�Y�]��4įn��Y�'q�d�<�\����; ��&��-���i��A�+�0 Mu*hy9�ݘJ�ۦ�v����	�?,��Gߤ�JVL6Ӆw����m�"�h����J��E�}0U-mU����ͣ��~��E�=ŋx��N��T� ַ=�*u��l1��O����O@g�q��.m�6�@�%�4�Tr��EE���a$�3uo�۸`������W6��	^��w�?g$Z������5����٤R�eq�b����~�0�O���9X�Eg����<c�CQ�}v�ج}�X��~�X�շ^�9�}c@��6�z��D��%<#,�~�� ٦��$��>�t���Yh�o��-�7�
�H*�E���9��k�p�/q]p9���o&�#QlAZ#K4�Y'a�G����c�3���SS��%X�WvB���X��/1$��'0�A0�ozSk�[��x�>j�hzT�s�y����f��Siғ}�&΍��� O�y�!�:]mg�aQ0B{a�����&���uH���2!��Qo|�t��d�
��]B����o��c�UD��[J��i<��1ڕQ�Ȏ���5�gD6����8�zl|�x��Zߞ��aWN�h͝-d����5� U�oUw�p��^��J�y��Z��hf֦�I�JY\6�?E�Y� myu�l�����e]L�~��b�Z I~Er�3�;��CL>�F/T׬�@ެ�3�)��	��ścI��f�6=���(�߭�A΂+�?I=Xl|��\[t��)�l�tB���a:(�30�C<�j��Z۬��y�Yږ?���)����<��b�=�
 (�����c���Q���~�����L��6���QG��*�w�� w�Q'{}���@uN��r(�[σ�7,��%r!L+�)<���Mˆ�a�)��W�X�nfZ�o;Q)9�d�W��������1��7{�Fe�T?Y��vZ*�b��|[�=��[υ�	�Ź�,vii4���>�2�R�%_}y<SʍAM�E�j_V8+U��������/�,J�%<�<��~|���/9���f��QfD� <��1�c���ҐA�Ѵ���|�����)�������#��D=��:���N�L�]q1h��nlڿ���s���!Wy�`���ϲݳ�F����~,B����[rg��cq�X�9���	����ҫI~M���j����$�V{�}����s�\�w�Q�O:F(h��I�������*y�_Ƒ�K�y����F�XiQx���ojnN��x$�m���t,��k�m:3V����EW��o��v��o��8\�8�E�H��j ��Ȏ�N��y+_���V�U��ݭi-��j�kuor�%�rJ��P�{?pv�i����j�gi��k��cN1#��Sis��F)����l2�K�/;Lc����z�q)�R#�J����&�B|J��2��_+V��h/1ǝ#.B�E�>���e6J��Z'�*�k�]��[��P�/�=�#7K�(�:�VK=���O>��2�OI:���]��Iϵ��C �XK���$����K�'�5�LRL9N��8 ��y�ܕ'
w��x���Q؊��MML�HDYj������ ��%6�>�����!fS1̬��دI����u���`���N�%<��(g�m�2)��X}�]���ܦ�_\�6/_[h��k�#�󺤴�o\Xxd�G��gS{k�x�u�zT�Ԯ�X>��j=�����2�x@|��o��4���G�p�F�Җx/4���V!��$4.�>4���(�	/aN��j����ō1�0M2f�1�#���T�����ښ�MҺ�{����ehcY���^Z`���篪ҳ�,�^�ѽ����ܝ��z1�F�.�Rfj]/_�@+C(]ۭ%�4��ƞq%@��F��L#��;�a��w��I��H���a?M�8QS�*�QW{UK5\�풸.����p�K2&�ce[,��;�ꥩ+������d��!��/io|��hΞ�IN�Mo��V���R}�����Oon�� Gl~�F�.��b�{���[ә�Ո8+G�����).��¨ant�N��4�f��L���E��:c3��ZP��nO�-.�8|�� by���O�s�.
J���4)|�B����J|��� �b��Bw���@�sW��֕��YZ�-~���-Ѹ��"�4��j�����<���ޯ��N E.gh5�5��5�8z�Ym�0��Lf���+Q���8������QSO\�a ����+��
nk�£D���]���f���:%�u���*F����q@ �2�����<-/S]�xK��ŗ?[�х������ňl�8 �����+���^�B����&�n�I��n\�3p�]uդM���圛2(`'���p���u����cz �F/���[ZFC0'+����Ӥ�~��@nb�DM�t�&��we�l��>��)-{0Gh����>���/�����ΗYR����"y�1�@��><�xQ
FXΖ�[퉌� "f��}ӺP��uV��!����t��0k�0������2�D�e5c�r�J����0ϯ�i7"���k杸-�͌�_�T��#}��N�]�3� �q�-v�!����T��.�.&-f�� q?uzL�u�y([�"�{o,Q����'K]_��?\N���B-�$^%j����Ep?WR���\E�v�J�'�)�K_9~ �)���Mg��d���Ǻ�S_O�܈�RO���6y7��vs?�YOg/�_x�.@���x�.k���B�L=��,��ת2��ɸ �����
3��(� x��&��+M��0��kB{9�K�$��	)0��	���M�l�:��3����:��b�<��Ǎٝ-8���؁:�+\�����1�\�/� �y�W���IC�
mI[a�7s�1�f7���r��e�|�`V���Q��9���!�����ɷy��^ ��_�����=�By�؇S��̠L�
���͸��|#稗�򕳱~��Æ�O�><�x/7@�.3꼫ќK�Q��U��P�갮oq��&��zx���l�1O7Y�vh�b/<X�d	�խ̐=� �+V��u>ߧxy�ו	 ^�6!e!�<�Q���Sn��|��L�Q��+�{�,f���������+g1���׬��:�t�_y�����GcW$��{yUgI) �1�,'2��iN&m���kd)��\^&�;�l]�!O��L�]8�hoS�јؤPۆ������H׵^os���?�2��x���_�H'��<˳�Ƴ�Uc�*��/��/�}��X� ��iq�a��1r��R'���1����6����Ӓˁ����� �Z����!6��X��Ӑ]_�s��k�ӻ_R�w���{����J��kk�(=07ڞ�E 9J���HH@ ><oc�r	v}G�����YS�C�.BȲ��Q�����;�S=�˅K�[��@��j�.Y�61ԝ+nj����a�'�v��g� +<1њcvS�|'��[4��@��B�ѕu�-�B�ȣ�C�B�� YÜm��=�o���2Y����'Oz��_� SE ���tN0 ���RI/�(�\��(�$�̰��%MhR �����8)����ثL� ~N��HZ�z!���{M�����I5��u�2��r�4I�}�}���U4iй@œa)��'�=�� 9j�L'5���� ��v}��G�����b;V���*[��(��q��^��ӻ"fGٺ��	>>x54o����au� Q�������lR\v��" K��������C�:�j���l�9K^O����{���ʂ�OiH\����擛�@팛p��eX�3�8ds"
�>Ű�8��l�4���p�F$=�*��g�~�dmi��07�uW|z�@��%#Z%{�	R��[�4 eYw� _U�Է�Qc�0�s�J? ���@h�og`����2�1�[�����+'��y��I�,���g)A�_Ip�E2҉+m�Fq��^6MS%MS��k�ǶU�tY�@I|�'�a�Y�ׄ� F��؈wrz]����2^�|�#a����_�B˵>B� ���a3j˫�᳣�!)����BD!q���f7s27W+�%B�'���m�3��&ʐ���ޅ�����W������3>L���E���b����tSE���T�I��,��\�o=&�	ş߫T���Ժ�8�k?�cv���ˀ�|����p��V����o������O,L�ש������+7xʑq]F-�5��Jrj�oͿ�PK   yX�_B�   #  /   images/6c59188e-af72-47f9-a95b-923959af310f.jpg�teT\��mC��Ҹ�Fmܽ�	4.	�N���.��K�7.��� !	$9����wǽ����ػ��Zs͹V�Q��H4 �  �v� ~� " �X��dd�$ddTT��44��T��44Ԕ�+5��������@M�"����+" @�$*)�/��/�����GDH"!��`bz������/������W��_�?��]�z �8�Q���N�$E�5 ��׈��[�?&6:�ޫC@Cb ��p01�����=)&9��%�����m����Whjz�4��wC�(XQ	ֈ�~�<s�^�Ǯlw���	�����ĺ�I�ޯ�q��@tL��H1��)X��S�0)m�B�E�XE�zQ[`��ƾ_� �,R )�`�g�j�%��;>�;ص�
0oSP�{�NV���S_�/�&�tCMk���UOj��P�!+4��z�_+��	��c����AӶڿhɃ:�+�o!x�Q!Ʊ�&�;�3U��͋$.��k�}������vl�~���·bl�� 50!0A}�觮t~J�#0%k��!�D*�P\pej)����3���FOuE�'�XԵ�T |����?9mP?~��׸3���tLƚ���ߟ�D8e�㴽/0VB�{���Rv���l���B�}�S��n��jyHdl�m� �����<j"�M���t�<v�u���R�*�bF�E3������H�t�0�CG� ���<L�yy�VV���ìXk��O�?�/��B��v�uW$�ɷ�|Bx/>�EůM��ڬߟ�<�+����Y�������u:��r?��e�"��d�o�B#�8@�i(�)�Z+�NDg���3KHg%�UKaK�$��x���R��VX�@��6���������P���R���]�����h�M�3;cch͗E_���.刦�L�������qڣ�@�m�[M�{.��h��֢OgB�g=��vB�K�A��6����J�����Q�q����r�l��QT흜klq��jsYf��ɩ�����F�OHa��¦Io�h��,���y6}h}�?b� ���D�[��W;5������i4=�)~S����;���(��ߣ��;����
��Q(���D0�)�"&}�w�2�Ϸ^��m�L�.�B"��'g���0�e�8�{�v�=N��lj����1r'ޭ7u�9_ЌQp�P���=�yҙ��S�x6\5�����)z}Hli������Ȫ�_�I�
�MR+���V�	K�+���
�)��a(�gr�9Ğ���F�D���� ��E�A����ߗ�X����pU�C�=K�U�R��&6@�Y����V�}��6%�_h�L����7������-`̌ �C<�5+�aO�^���,�L�����k ��by.�Qu�8g��:�8ি����:���=�gqp�����UQ�������7�?Qx�b=bSK��F$}��\��UV8����U�P"˼�a��]�:
�D�/5W�њ�ڷ�o唕�]z�^�]4��Y�n��d%�J����d��4�-~�r��,�E�"�8׏3=CQ��m���ߌ���6&1J6���@,�,��a���)	��P���� �����߲�����&��w��G��LW5aw-�@d�����U��"֚N��Ә�!(QU��̐| o����P{r��K-aܰ��)��c�U~��N���!��b}2�<T�,�ݩ���.ϐ!��ׂ�g/#�����TC��EȄ1h+S�X��WR���li�1��y(��x����j0���@D�j��&��\g�%�)��ڂ_a.�es\�y
�Y�C\����
��z�^Tȿ(�`A; N�e1x��Co�?��C ٷ�������#aD�E��3 WLxmF��s3c��ф_߼.S��5���@k�c���O�#s �0�m`��M��']fl�՚��<��{�{]�je|��iG�_�,������4OgN�۞�ڴpd�k�;�B���[v�� ��l%�汚����rvs֤����v�ǭQ@e�;��ǲ���,�oLThL��"��p��7�h�.ζj�3ZI��5�y�<��%?P8��R����$6Z�f�c��H"�̸U&tf�=��)Ƅj�R���F�-7�E��f�dй֕Q"2���9��G����i���CrG�R����=�����_�&��d'Z���
�$������c����*ݷ�U��c{�<"&S�Old�ր�^��-��^��G����TlEI��,#d��p�ǜ�]L�Kx����=Jй)!����|24��Y�t>։��?\h��~$�)��3��ϗU���nMS��bմr!�y5���1�!E$�@M�l�ǀ;q&�i��@q��>7���2$�`�qY�Pb��R�67���s8������i?�ѧ{����;���1Q,��Z8܎���[?1$� B0{.���yAw����%�t�3��J)��ګ��!BO�����%�o�c�R/��FG�Q��T�E�]<����WB���v�Q�2x�be��u�M�f{LK�h�-5j��[���p���0| ��9�D���OSy=�>{-�y�U}�N��&L9%�Jt�xX��|����6ۋ��)��D�"+G F���$�f�	!X�[�ᩭ9B5O5(脉X�m��`��jj^����Xt��ae�(4�̧��N�SH"Rj��G��l�"��pSŤ�����rc�H�,�	�rKǬ4�K�g��ڕ\�bui��k����aE���(�ƇJ:�ܮ��u��g�*g뚶��MeWU�&��+�b�\W�[��:@���w���%V�mM��L9�M"_F��M���
L(�>5N<iz�U�a-?\��X�����]6w��}��T�N.	1�ȣb�Y��D�(��N�+6J�	��Xz�,zb����t���ܮV/e�/�Di8�.��yw�p����<�z�h���3E����n�[Q[�����,͓_�M�+7�Ɔe���5m���vswъ�8��l�D����S��}�(�>7�V%8�͓�I�S�"$��GcV\�@Vi��U�{+�Y,:$\'���ɐR�dI�B���M�Md�΋�є1�,�<�5.��DU�~�_d ���R���H	����;��e�<�ˈ����t�k�jX�a�+�%�,Յ0�48��٬��{]��Tҳi������P������W�!Ji�az��G�q(L,li�5ދ�d��t���|m��q߽����)|(�P��|��^�$߻!G�z��y�d�ŻF�H�C��꤫*i��/g�9ڸ(Z'�c������C���km8&�!���$�Ѧ��֗)-wE�S��_ZQ�ɯ�M<k#�M�[�xv�$$-��s��j�>1U�p����)%����>�Wք ��ܵ�
���(��d�D�㒙��']��$,��:
���p9�L28���Ͼ�ys]�m^#Dx)����ʘ0�ܴ�qs��s�_|l
ۊ�������e�����Nmw������hJo�΅S'�����U�sHWJ eF�Z�i�iID����1./��Я��ysGC&���#�aq��w���E�j:��*����Z�^ ԙ�7R*���K�f��8 ͻh����^��0n�`��A��"�P�Ƌ	�m܈!��̮ZW���ζ0����m(&W��\���vC�1�.-��N�@�o]zg��J�+��_��VCv��yG![�z�Pچ�����*�z��p��YfM���
�d������|��唶�,/m�N�b��>+��q�%��T�BR�@u�N@N����'6<���N)�1�b���R��J$��_'Km��?i~�H��о�m�ʥ��,,0^P��I6*�1J���>���u����^P�t�ɟխ)����%(U3��]��63r�U��'*ah����^�f�1#��=xӤ�[?���4����b����y���E{T��0�K��I��6,(�#O����Nչ��t� {���疐��پ��`2�^1l+1Fe.�����n���Y�X��]x8/7�*"��_������b�A�O��֎���p�j)Né�ܶ�H� ����TM'��-]}���)�(wp�N,����@~$kg˔�����u0�櫊4�A�K~�T ��}K8"�,g�?����
�t�������2G�^*G��4�~u��w{-j����� R��c�!���70f%A'� Դ���ug(���3��ɲ\#��Ъ���:	۪,����ӥ+ͫ�b�%����wCs���O ~��6(V�[�ҴX�R�6��gR�d|���^ިGN=�e�E�5 Z�U�-��"��Ǩ��L)Fd95;��s<$?#-��g��G�������$���|�Q�wk�QU�"ba��1�b��0�>���&m|M17�{߯RX�><�M���&D�xn���5��I���w�=���T�'X���d�f�	f3�\8�����X�0'�;��8���zG/���X��"Y��~=[�5�1/O���N�\�9�? �l*��k�r��^�:�p" #H��^c�B'�9���}����"��ƭu�<r�]���=UH@�L`k��'�!YԬ�Vs	Ư 2w��W����/��D�S9��߭���^�C%�H�0�+�jy�
��rlП����.�[	0�(�"�y*j�ئԵ��i*���6�[<@+cr�+M����,H�"%��og��,\T��dB(��Xj ׉c"������n�#j71�]�����_ <�K���S�����o��\7��o.4���<��ҡ��^�D;c!�fb����4)4��� f�5�@��ɋ�D�M�h���NXQ�{��Gґh�k���V:�wSmY���r�g�	x|�`�� �6�y��u���@�ol=�į-�@�?�}�d�Ⱦ��౻#��,��˳��c�ʘ��q�-��?eI�sH���n ֠�� \����7��ɱ+��!Hh,ս�Js~�xHE�i��L|���KPQFҬ���۬�!����(k��&�V�g��g�~N̺�~�r�i�'�����Toy�g\LZ��*��"[�R�]�r9bIdZS���Zw+�b\�AK��ĸ����7�����I���-�28���A?�7�#�Zv���u�y����md�,GOԑ�.屏<ƽ}m��Jw;�
:De:YL���e��}�MX��j���k*
X�h�u�a #17���?�hm�%Xj4�����
y!���ͮ �LT�;B�!S�����C[�)rnO��	Vf#U*bM ����D��h^t�f�*��D�����)�	�C�Kf���p��s����M���.1n��J�#!͆~-����Ж���ic��%"w�,^�/pj�a^��n?{�j{�Y�_s���	B�Q��@F�@�s^����yb1U�B�=�HF�6��[�i�	Q5Q58���`���a�����&���i(�>;`3��Ht`C[���w�3���?��vT�lI�� k�b@�/�Ǎ[`o�x֢xj���Gh���{�咎{������)\B��҇��r�G��R�ˈ����n?�o���/3臖��]о���z\���A��t{y(��4;	hCP,ב�=l$���e�� ��I�t������b��B���R�b]49���Ѳ$�@6�f����}{Y�-;ӽ�=zg�r�wh���[(��u��H���le�	��yyU�uO#>��d���F>�Zҿ�:����V�_ t��/� �#��/d���|����� ؛"��wE�ߋ�9oƃOko=ߧ�.-�, ��7 ���τtxT
?9'���~ڒ���䏻���}�Ww���T�b�s�q��-j	��C��>�!��_��ys*t8�]^�_�O�\W*�i�ߍr@AC����W�깜��m��4w��벓!�8HuR'�������˼ĸ��F�����G��^G��AB��1�=�wh	��S�����r}]��(0��b��ԢeU����wLm.꿺q�/��[xJ5O�T��F۲���c6��Vt�6V���w���YlK,'�u�+���CU�p�h�-�������֌�z��Lt�d'������n�~����#�#ׄ��c���^�:7���|zմ1�$�՛%����0�t��d��<(5M5y�;rБ���yBl0�'Ie#��/�W�����{Џ���jD._x�~s�!O�6�*��h~6�p���_���:j�gl+���Tj�d��Z���KWv�u�;�~w�̌���(5�P�3���Dt�$/nZA>R���/;5��:���(5�w�����=p"�t�.�f�ol�⠜t�|u�f� �����L��Q�ql�g�2d.�P�j�~�uF-�\ov��S��J����̾Q��q�.m�FGg�E���Û�3�%o}���q/�������6(޼3��k{/���}M���y�p� !�}K�G�4�����%0�����}��i�?Ϻ��2
�h�gy�5"BYX"�ó(P�OG��嘽��&d%1��`�@�����U5#�e���@m�̽C���2bw3��/�d��q��J|��%�<�
�E��c�=1\֫����d:�l�_���ʰ�!Y��wzYS/��z��E�E$А,�KHg��d�����|��	�d&��c�,�Wc�R4{y�LFn/��Xk�4-y���ٶc��y.G��X���D~���HM���+>�O0�Z�Ҭ�(��Dx�_�p�?�����c��h���+��|���=U����{UI��
>��w*�w����攓�x8�ѽ��_) �˖�+�%��������]s\s�q��';�����Xؒ8��k�TqXTUj�qɔ�`�j�^ �7,z�������swu)��%�1�-�̀�V�N� YH9�B�oT+UK�V�V)���hhlG�/���AKq�-Ӛwۗ��+�����+(ރ+����b�P)��SE\���g�g-��x��?��ucZ5��]mOn��>�Q�{KA�:�|�ִE�\?}a55� ?�A���4(>	��D�Ƿ܌�x��${�,(}~���Gܻ��*����S�O�_*?�]|�i�cY4��=śSȂ� Y�ɖBj9��sC��`Q��@�� (,�/6l�]��� B��@�����J�����h@J�-.~��p�v�j���RxU;}:��=�3Q��dw�\����SXX��Ľ����B���R�`e�����ќ�(hsI�=���a�8.b�
�>*�u��~������4Zl��F6S�3(M����3��jϐY��)Z��eCE�Ow�ut8�~)�۱n��j��Q]$�BѦ����q��gȏ���
.;�;_[���T]�^��������i-�o�:-��H8FE��?�XX���.-	j������6�=�`���/����>��~�7��`���L8��ɕ�U�_"������5cTH�~�k�筂����}\$q1q$�Ix�<����
Iv�P���𯭸��:�->�����E0^��Lt�����V:��U�©|���PU����@0�yg�d�����tP�@��cOx�V�|}���$}�[��|���Q�,J^��N�(���!�����f�\v�%��C���ޓR�����drt0��@����7�����A�T�L�w:�BofO���}��g�)�]�	0gNF����	��yt�w4Nf?�Qm�F��/��aLf��|��y\�C�]`��᳎Ԉ��.�j��{l�����}��6�*�O!���kw���Ge�[�/�����|��S�-�w�6�?�?��w���@C�85�u�����F��L�N�^`Z���`�w��2Ǐ�l����-�	V�6��A1٦���o	_�F���Q�ˊ���O�v��6x���р*Y�*��Gi��'knYv\x���Q̸ƫͯ,�Q:����[�o�n�г!;+5�syK��@���w�idd��n���b$��³|���d��g�t����(�t��2C�=X K'�Vċ1�[�"V'D�.oQ������B/}�����5"�,����uN������5�������Lm�ẘx�Nd���I\[��(�L.I����s�*�"ЋXI�"b�"b���\���6�`�Urhs֤��wA�:��v��U<B\!(wzU�� �� �m���*��{�x���n��;�]�����2�MKF���� PK   � yX��{	  -  /   images/84b7793a-00b6-41f6-9ec0-c4aab3fc9029.png�XwXSM�MD��DJ("���"�H!b�RBo
W� ���D�	(H��"DA�J/�K(	����~������?;�s��3�wΜ��sga|F��w/�����1a���t=K��a�R��6=����,����D4 0�k�Ƈ�y[��aaޞ^�Uꒂ���TwH����m�����$�?�3M����s�C�G��j��j6.���رc��+iJBg�޾/���%f�jO���R�^1�:�$A���)���V�n!�C�ip�2L{[T������ktdP���j.���}��z��������U���x&�R���7���ae�>E[,~_��q7�L�5M�((�l�x��T/~��r���Ou�	b-�䶅T}������'�[�8TW�X�����k`r�ȵrq����=%�s��W>w�_����stt�r1:��3���VJM��0+ӎ���������=ƞ(��=��[�p��[%�W<P�3��sQ^ieG[�y�VX���V�ݩ��H�g\�맕��R����|�t����9���0���X��x�Y�`0|Bk�����bj�kixG �+��/9(�{b��Q(�ӎ���+v����CCb��,!�b�!a�j�h������p.��)!ؕ�n/i�ı�;�ډ��y��5$���c�k�X	�? ����^�Y�i�����	���bj�
�_rPW�SVTV�*)c�T啕pʪ8%U�?�k<o{G����?Gciξ��8,6  @!@E���URWW�**c���Yy� _�@y��t|�.��.D�5����WCB��$�=�r����B��h�URP�����y�y��1�=����������*���t&�}�����^�� �H�y,���}|O���s��i��������Mp8��
Sr�����`�K�6%�~���wLb�*
�b��.k=2���A��hH��,��"��b�t���S>,�x���7�!���1�?CY�U�))��E{;_��lO�9���XSvq�sr�zz8I����8m�ћ5�?\��=||�<�:�{�"�^��N�E8E;%���T���Ԕ���j�Cj��TT~��	~k��mo��7�va�.;���ڞ�Ó��+]A2���ן����<�����!A�#K�v���+�7� g����|���v�ǝX��_
�
��3���$���ow�����u���U�<X�˛U����`���q��Ω�����\�mt������F}���/~,\X~3��hr�פ)g��:<�!9��q�����+��<g]#z�P�'I�Mt�O ��r�U�,���N��[0�^sz�L'c��9�ws3g������ژ�6�(}#��a�.�����m��Q�g� �2/�A��+��z��[H�=�"#NGH,�����c�_��֑�L�;��/j>����^,i�dߛ3�Z��$O�9WWq�� �/�����ad�S���A/7�
64��E��?�=��E�y�3���)!�>Su2�u�����@�f����4�k����H�{θI?�A�̟aQ��	�6X6�ڸ���"W�]�?T��f<5.�}'~���k�Z	��P��ظj/ЄRo�E't~�FS`�|��O����K�h��S6d�ʢ��&����e�t���&���˗��Zd��~�a�͝��K�P#�ENC�V��Cd���;��� ]�7�vrx����Y�{����~:� }LN1���KZvrP�Jo�Փe��]����ʏ�ކ4���5�З�N7�[���2F����B;Q��@=Ѓ?�>�b�"��l�L@�h�M��\�-c��^a��嚂s;���y����3�,V}���j�.�df�>���[���F!md�+�^��q�������,�/�h3�d�x����߻-�^Eӣr�3i#�Q���A]#�<~�#sq%qr�S9]�=�˅��m��e)	^�+�~eDL���U�Nh3��p=0�h���<�<��pD`��+�-'��Fg�0���G�,t��� �V����1���V$�<�����t���b��5Jf_�\ӣ��zRZAn���
�e����&��x�����O��Y�9�F��wߑ?Q�>5�5�׌3��>6o�eL"nm-:g��2ѣ���O��$������gg%%��U�^P���8B-�,mH#Z�8��$�
b�}�go�g{��Et�/�A^c��������kg��Er;��U��	���j୽ɓ�iVV�]$��C̷oA�C���l=Z�8.
>�N�Ș8���9�ԏ��l�QF?5[*5t�j�B������mȝW�����F��?	<���g�|�Y95$����9��%�A2L���IM��J����;�E� ]�+I�M��F��l��2��+�1g8�a��+�g���Lzx�g���4o��|z�)bq�ˎ� ��>��n�\E�[m��"d�4zr�k��W�������
^��X�!՛���EUbԕP�̳�����k1Uy���W:���*σG�c���W���gF�_��8j2��`�����o�{A��"tӗ������uÝg��p��$�=���JN��7�`y��JLoƍ�s�S{�w��������V��;��C	c���N(I�+m�	�9���;�7�%�]M�OM��;t�y��*�u����1@�iS�yT��f.�@h����fY��$%߈�&ײ��Z���������6a�W�� 9��l�1]"]c��,�?j�#r]ԪiuOV��Q؜a�*������U�7=�C�;�b���e�I�'Б�tkZ޷3���Ei��H�ڞ�u$;�h&��ǉE�gUT*���Ǉ_l�iVh��AnE�#A�3P�NZ��l���	����oF-N���yC�v?�5ߴS�Eƒ	��ӷ�ْ�ZV.�[�Q����V�}�ܛ�{&vv�A�C����o�A�BY�Z���s> �R>�2c3g��<�"��V�׭�y���e�`�AM�5�x=:�L�L�4�4�>�=E�u_ Z,��Z]l$����0w�(-���1��-X�mkWQ��T�s���eXDm{��^(ѾVQ��R��	c��S`b�*N%J��ݿ9YO�й�όb�eO�\���ba���Vd �k�%s�{3c?��^n�]+� �l����Yn�����n���Fjh�ٷҏS�����0�O��T9�@M}K���%㴞h��,G��F	wT�x��Ǉ2~!F:�F�s�ř%����`�'�W�~+;_�d2!��e��h�eV���@�@ޡՋ� l&�޳5�@��IHg����o���^�2L�9��*��8�6T�(;������ 1��a�5Ő;�y �	��h4πg?x����[?ؗKSIK�gP�+ǅ�^"{�uE��p.oN���p�5������04�32��?�/bP�ka�W�0�?�~r3���\%j��m8�ِ���Z�8����Ѽ�}[�Ե@Z����`�ٰ,��d�xDï^�W-Y����=��o��bn�բ	Qݠ�ˇ�R;ܭ�:(�L�3j����O��\ [��*Ћfx"���(LPa�#�"兏��-�Z`��կ��(��"��4�q�'l3�bJ/��V *:�sS��hō����|e�S
:�gO'��HG�;�h`U��J��Z:3A�2A�ܘ��{+�]�#�e�BْFԙAhf7z���ɽWS���N2�:��}�&�!����������7A������>�hMT�#�q3F�[;��#��6�ѠR�}�i�d3�r7ڙ�C����G���y�ҋ�$Ԣ����h�_���{wυ>N[4��h�Y�#�.p{��D[��<��eBg{�" � =�`n�k	�4b3
��P����}��	/$�|���PJ��]���F�����
(5|�<�i6��;}�=3$��ϵ�Ȇ���vd��S�����!��O��ڱ�k��޽ �-%_�G]r�l����\ۇ�l��'vj�b\�1c��gD�o+��B����F�i��F#�(���;�%CiD!�)2��t�[s[�:��ī��NoKY���2o�#�B9��6
�W%c�������\d�t9Y�c�(J���UZCsz$P�|F�{���ާ>�¬�(p�CGO[���>(=�NO�7-��_�i���6H�z��\�N�Ci-���io�ѠOp��Ew*�c�;d�	�q�����
~_��SΖzx��z�z�K{����� X�e0��<��U�,ު�����f�����n>�GL�T�5��6�=��E.k�OC��6G�(Ti|�朲$:��t+X�����.|d�����;�W!��`>bys[#^�te�V+W�Ɔ�ud�o+�(G)��~IN�!TF �[�G�R�/�W����Z���%�Z�7��(�m�v���9���co�3A�s��qp����D��6�[�@��P��=J{r^��[�V��u��	j%r�P���u����|w7�J8ol�f�N�R�<�-���`�Vж����_N�	�Ol?z��JX���!`�N����� 5e���xb�����@τ���
��Y��i�'9a)��@�� ���HU-%���=��v?��=�6�@��U�\������Z�˿r?�b㧚����_yua-��S���l�Cg7RZ����U�Bؔ�EV�e���ݛ�>co���ߔ��y�.��\�8m,�灣[���UY���UµWJC+):��6�^�s�,��D��xy��꼰0�j�U\�[�J3�jTy'��}��p�yk�0	��Z�ƺ_�h������D"�H��r��@�-����O6ǥC�j
�Q`Uv712S>��6��u����rӄ������[��N�����ɈBԕ���Z¨����v�7d�_V��.`t���+��p]d�A��D�lEy����T���f�����a�G�w{z���J�r}wF�(Y�æ6Cl�S�m����G�����:��ʬ�n�Z��2i�Y56Y�/,�6~sv2�>+ݻB���ƭ�+V�U5�Xy�!���t���<�m���f�ۋ77X����@D�u�۔�G����<zE%q/㗇}�n�L�:{���i�).�)o-	����Hڅ�����QP�:p����(������ ����^߅��zC��1��@����,ΑBA�����t&��C&Q�_���	�-�`*�����/����]�����l�����W8�2X������^fձ�o/��ϷA�2p�ܣ��$�c��~�E�k.,����_�z%ո^D�W�o�	����`��)}�6~�g�d|ʖ�tHd�L?�������d����se��f����=���XZulf�y���׷<��sy����y��;�9Î�ս���~��}�;���=�U��Z��9�U��3u�c�`э-0�W�)�gCL�����=euP���<� ⎸E��U�q+��i�s���LʠM�l~`{ٰ��kQ`,�=�j�I��X8�����#��]�Zt?P�Nk������b��
Z��Oh-� W ���s5��kb��wC���|c��򹎼Z���������n��~�D���;��W���޶Mˋ�����P%;s�^�y�u��(�2Y�U�����dY\Y�ǧ�ǥ���<�z�ބ�Y�<BˢcWP��#ܛ{k-?RA9�u����	_��3ђb��E����E4���.����Lj�'x�$� ��E��3O���}y�����'���j]�7PK   t~�X�IM��  � /   images/86917e2b-5e70-481a-b4c7-aed39e2d087b.pngt�P�M�ED�~�t>��J��"(�= �	�C("�T���B%� ]�=U:�C�Pn�����Ν;���{��s����Gm͗tԬ�  �N�� �
	 ��s�*��!k��u�Wƞ ������r�}  n�ʋgz~ikxH,;1}�p�'���tn)E�EG;��ſm�3��ͦ�+m���0�΢��d�T�O�B���Țq�8n5���t����!1w��?�#��M��έ=��ݟm����gv�CLŻ�32֋J�։4���VV֋� ! l��!m��)_��.�[��]α�S >]O`�_~(BiJl#r��lI�.� �`֗�0W�a��?ư���+OϽ{Q�����1\��yQ�鉄Lc��l~�}�(	=>\8�(��z画~'w?pt&eHCwQ��xJ���'��XHP�F	sI[�ܛTN��n�e_>̎�8iHLv;��+f3�W���i�tU����\� ��L�o�"pUMI��Ol���@Y���;#o�s��Ōحj8���.aS����G�Yײ���6���)�*f�r��`��������_Z��#�a\x�;���������n<��㛪�k��k@a�����v��@��Dy�]d��PUrֻ�����bJ�/���>����k��c=��BV�V���?�N�=g���#�:�|.ƍR���P�t����B$��9EҾv<�4$�On����â�gP�ֈ��U��o줼�ْ֙���W��� Yr�
��U��2�߂DUͿyv��L "�H��+��P�J��.>Bm&���N���&��ff��c�a\V\}w��<��A�����|}",0��K*2�����k滠4��M��7V�E�A�b���W��CH)amR&R����B	���M���3[<(Y�z1]Ǜ���F�,����\R[���J6���2�&T��,��n�]��%`n�w�4fB\�}4G��7۔�+.g�����k��;�˳��!�W���mQ`5���ϟv�f��kTB!�̄�	��Z�QS�e�~�s��8�����e,�3���"�=�G�;����C���1�\��3���7�i@@M�M�	>w��k�or�X�K�0a��-/iB�Kt�	�%ai�J��W� 俗��W��;kTY�<����H�T�g�[��VS<Zeֈ֓*]|q�F
�����������obE�|W�"�wD�Ԙǒ�+�=5{�n$��Y��{7hl���ͺ�-z�N?��3��?�ܰN+H��`i<y(�y��^�R���"�±_?�w9�M+���g�2���Åg x�����ٙ΋v��������k����l�eD]r0�i����z�2���}�&���]�k��zw8[�~�DRa�K022*���M.��:����S|R|�]%��x��8۔UJ�&���(�W�����]���A������
�	���"ͧ_{���m��{�	b��\��999c�$K���vsf��@śN�nX��c	q����U� <�m��S���������FG��ة��iҌ#օ�q>������q���xT�0��SQ����Sc��YԔ����'��ƭ^�8>N��-�rF�_;�F�)?o@|�ڴ�h{S����w�(�.͠�T��񒕀ُ����_߈_�`��?#�#��z}�V/�/b��Z4�A�%�`��OĉU�Z#A]=���Qe(��A{�� {�nu@<����莮v"��2�Kr�x䱶������Ӝ8yoε��V9(L&W�k�M�r&�D�t�����TW�&�"M{w�\v� ������*��Qm<����2�g�i���wS�G N�[{:Ϻ>�yu%N��k���N��V����F]nI��^Ҹ���3ׯ��~R98�l2)���"�u������_%�����˞8�2@hkԒb%ĳ���_$_�yD�\���/(��K����]N��`��M��o_������X�#���k���G�.E�;�Vʠ 3+G���<;m/H�!{�P��I-+�Wפ%k*e�wih��-���	B��;خc�jD���}����?ybbշ��깠"K�u�J54����-��7hpѫ'�Z�ʘ1�ԑp˦�)�T�&+u�/�F�y��
������7����%H���ތ#sD���rC��\�\u&��'�|�����m�?����[����t��kN�f�9%&&z˝&�V�x4i��bT�^����^����>���:w����?��!/K��j8P���㿹?�&b��=u��	[�<=]��T�᳻(�.��n�YA�x9�{��a���,��Rā��/��|ҏ�˻�+�k;O/��|'U���</��h�J��o��Q�Z���B�f��b΍�A�NfF*�4�f����Ir"ݹF��F�.tX�R�>�1(M�J6�QE?^܏����<b>�]-��)���պ4�%9Y�ʤ��?�߾\�4��a[w%�UD��q�)+S�z�~k_9?�I<��a����G��Jᖻ&��q$���L݂�_ªx_f�BW��"��7���i���*��OX�K�,��M����f�3%�#-�:��3�������B�a��Z0�P%&e��8���Q���h�d(ۗ3��2���#�F��#�[:�El~���e�o���L�G����2���+Cp�zP,�>�^u��e����,�Ӽsݭ�X��.3?���Mx\�~������թy���5��]���F܈��U}-Is9;d���I���q��B n>���7:c)�P=�e��_�
�?v�B��K�<�w�����L�M{EN�� +FF%��=h��Ν�]�tN����<r�y���gha<�We������/�ؙ�^n�~&��t��m|,��pך0�[*�zeZ,Јj����ږ�0������`���G��Wx5x
�9�DO�}/�ǥ�S�2~��Sm�����F^��`dpc6���7�m���F��ݘ�j";�£�#��3�֩�oa{�.�|)fe?�I���7�m,�}��,z1�U�i�ľ�����!Kjo-'�j���)�{0�/W1Ex�ğ��}Z璱�^�F�|�����U�,`0�7:33#���E���f��x�T����nKU��т.��!X2ܻ����%�ť����?-� m<x���k��6dJ��!T(�.������u.##=�cXG��A"(W+�F[[ M�����;�����U��/��P�ØWI@"
��#�ݝ\5]���1���#�^65�XZr?u"�OOO	y�^3�W���yZ֚��6+���T��ZT.�Y��X����Xsã��o0�yD7�Ƶ�,��bXȠ�kx�tT̖�<�Qe����]�5��/�U��ܾIr`6JJV��P��s��Hu����k�$���[�
�s��$n�_��r��!^�$	�F"�#r]�V��Jl;���|�2j��zy���]ש��#1�b�!w�3�B��j����븫.%��d�S[��;�����u_��٩�t�'ߚ�4������;���2��^4߇��=Wk�A�Z��4��K�$�<;�&%W�eR��3���>+�@J���SL8 0�0Q�%������Z��L���V��o�9���>Cw[���OOT}E� �I|��p�u1���Z��}5�\�7��y��_0�3��l���Kf�TK�)�����3�����g��ݱ+�'OV�S�����.��QS4!,\����
\�������,��9gʡ�G�͋�?|~��ZT1?�x��=�`xnLKni�<>dbpz����B����{a�[����d�Cv��(��f�O�'�1�؛Ҿ���-ҿ��F�E�/��/��?hU;���QvBP���'=��|���X;���v��I49��J>��d��c<�ݖ0gRgv Cs9���m�E"�������R��Y��-�[�~�/AԒ;��A���~Z|��� 5�[��<HWT�����Dv!�Q]l�_2�?z�=�W�Mu>���4z2��b��元U����g�T�/�X��_��G�˚L���_�ƪf��=˖d]�o�\��?%\B6ʅ�E�@ �$vp0q�g'���?�N�L  ɸ�-��?,j�����P�o��k��QTj�\���'���\]XX��L5@�+�R���u8��/B긋����$G��͚�a�������ԟM=�:�G��Y6�{��.�~N�nd� h��?���҆3r�Ռ���y�LJ�b&}R'«S,����yH��duõD�ń`�l�����!���A��I��)���ߚ���q��@����	IdR����\�-o������y�]Ҟ�zE��Yb��*l���|G��*!=�A�8G��7}�y")`��<���Ɉ�,$�IB.@�
�z�>�:��u��a������w��ﻲMS`ك�l�\M��Kt>G�hŹӼ�"�x� ��ʵ�qbvd�rJ�����żu�hٺ-2�{����	&c�����_���c�cAT@��Q��|e��?y)���憽+������!������b���U���IaȚڑ�9+��E4-��Z\��z�]�E�(E�-i8�r�7�)�+|f���F��^�
\�Ԕ׏�yJ2{�C[���g��-6 ";���s27�;�Xs7xS��[�[�h��O��j���J>��R�'4���dzs��bAomqV�H���ǆm~�ǌX��ӓ)�ceBT+)uS{��ۤ�{	�}�ʱ[kr��f�i�x�cڂ"C(�`3��Iqx�y�%=
Zrh|�ED�����)��o�)���=}�Qr4�ҚSh�T��5�qu�^kF]�H�������6݃+�w͹&W[ME[-�q��s��`��X���܏3Ԋ �}Rn75�7�W#$�8�	;�z�%U�����JO��v��[A�g��]��	���4��l&|(-yɎΐ���'�ޟ�e��*�K�B}d���K(������������q��z6�X�Xv�!����b������İa@O�_`7,`|WϐT���t։�!
)�4V�d���£�>��ߜ��u؃u�	���
��*��X%_uz����KWT2�.�G���f�"��9��.1�COR��z"n���#�����ɕ&����f �Fۀ폠X~8������K��2Tp�y������c]h���n�ʬK5���5=�7����x����1E3�(
�b��]�3�B����B|�N�e�����VRώ{$��h6��!3�:��f���3d�C3�*V9�)���e�Хp���Q�g�>gux	��e'�Dc�An.�����o��~5���.G�a�����/�:�S3
\��	) 3l��]2j?j�H�ُ��XZ]�2xV}�:�=3�b@���	^!�W4�
�˞5#�5��u�����N�!��%^R�ׇ�¹P;@қ�����ۨ���1ͩ���ƾ���JSZJf*	VLI���a�Ѱ��q�J�)_��������C`�\���otú��ho(��#"��n�Jt��T^&��+7ƾ�n���$t����&ER/�>�HO�\�Eh0��淟UI(�I�=��c^[Ð��Dw�{[T!��bk�d�F'��Y`���_5�ҡ����H�"q&a��4�,[�0�a*0��2�htϓ8 �l��������z)¿���K�#辢6��ݚ���.ݜ�+����ևup?��*!�E�R�ˇ�W]��ee���M��{��5�,���3�s���3�[$��8��%�߱�g�5${\��'<��0'Bhel���1���W����L��Cږ�s�����~t�~"_28="W^�k�j×�o���ع$��s��%}�P��/+,�h4�Y�Y$&���� Fn����I]�n:���,-�x4]R�W�5����_�^R����fי}'o6	@D����R�m���y�<�dI?����Ax^Ĕ���i�D�N���|���Jޝ�~�?�/绉U�Vf3I�ݡ^���N!,�yWVo��͖u�N�/v#EA12O�Py-��Z�<�Wb�?ڷ�T�N~������kgD�a��{w�).�������9��E���f��7H��o�R�ݲzt�U��)�ƽ�J�"�������&h1�����O��l���i��Fo����
�{>���ť����X1Z�O��Y�цE����\yΓ�w̰��&.� ��G&�K��ث�@M���bB)]��E0����3f=좓x�,6!ˮu=_��dZgU�s��}���~D�`/ �O�u7J�&pV̊9
�zS�i1cnkf��WU�Y�wt��f=(!999���X먨(�)����i	�zj5�ͩ2�m�t�F�Q�Q�AS�;�斿�A���~���z/ַ�ʻ�1��)J�=vb������Qtp���gq���߾i]m��|��Le��)�TO��ݽ2V�'��~���퍛`��Ŏ�p
��6��3%�yZm��&��u5a^�3H�pZ�L1;*ڻ�Z�������gt�k����n����y˜3��W=���Q�d�^h�!x�����9XA8�$g��S
�adw��m�p�dw�Cy9t�dȥv�T|(i?�3zf�4��KtAW�_���F��B뽏p�G��X_��Ί�F���]������]-�&����\���ҋ��ME>U��Q�`bx.�#��._�$�Q?�ԨC�H�`��zi���za/�7?�ߨ���<2��)��>󊐡A�{��	./��Գ;"����s?A�܌��͌% �ïfntgʷ q��ϟyZz���N����L=��́A��R�e�!6x��ax	C�H������n���K��j
ds&��'�nb����NSa���[�B��䝶���B,�з߯���h���A�Q���d�Q���Z� �̊o�E�|��?��GD��e��Ų�scY���*e�i��ʑ�5�~=���)������Ň��^d��%L���S�^X�]�"�>������0�i*�R��X�h<mG�+5�����uՊA�B'���+̈��Z��$rt˒9Mf��i�ɕ$����]�i��4�H]&L �]R�c��w���d�&qI���2�@U0^�
�yA5�0aF�,��Cn-�w�#g�l
��Z��L�R8����;��T�>�"3�M޶2�����Y7���wwqI��Af���
���f�Enʹ�3`�J�͵�]G�8�HBs��a:��_��_����I*��uO�<��!a�-َ�A�FB����W�q���3:ۯΐ���v3����
�J<��� ��u4�c��	�Q?�,5d�PEHt<|�����*)��Mq���3��ҵa+%+��w��3�=�r�Q���N&!Y9��o�ƾ����5�e|��.��rf�]Yl̻�	k��o��gV�M�սg�Ş�&�(p�fXI��3��  �6!���[��,A�O���G���	��l-���Q��8�v�*iD��ҷ��]:�~��0h�$f���FqCPЬ���.�E�}��YH=D��7����+����|��'��UN��0��˘>B��g�!jyz�jk�{A���QkqĜ�����
�����T������88��ZpHE����1?�����@zU��-r쟛eu4&�\�jF$8�������b�ī��x�k.�Q�E9�y�-ε��<�	l�ϙ�Q�Y��KCƋ!A��7?��� �j�p��,,"޻Sgt�5u�w�LIT,P�P�u�T(��/��c:
�gqEj��֊�����Rr�9�D��|�r��FF{Fp��!MUE���
&)B���W�YG<��cx���q�wYX��2�;3��m\�QmY���b����+�y4dq��3�"�f�e^.�aAX`>
.���g�L�6p�Dh���m�q������^\o��� �s,�EW�=#��K�`(S�b$��2�Bv��VW��n,�����p��Q~����xg��ƴ�T��+��zۃ?Ͽ��(  j�/�r����h�&xC����\y��%��8X�f��+k�H�͇��-�ܘ8��?�R˝��xD�6Km��te>�|�m�T�Dr��?�|1��w3�4�;c���n،"ո���\���	�U��ĕ�>$r��^�&'�<��"֜2��N�G�|֐T������w3F����w����l2s/͇�M���}�'S�79�)�1oi4�i̔o�ۤ@�[�U6�Q�KI�$ܘC+���� w5!\^R�"m�$K�=��:`YY&�����Q�*[���J�8�͉O��T����>Χ,.�ppY6g�ӛͅ�R���B�	l����Br�8>�wR{���(��6���v<�x���H��"_��l � ���"�����֒�|��'p,b�P��D~b_�5��"�=m)��gh�ܪ�1���\^�(�X|f ��t�ʸu�ΊZ�d��a��=�9 }�M:�8��8,���:��8. A�Sg�u�Vuu�Z)�/��u�g�~BekLW��&$����.����kՙ�Ř�̦�H<@�E�S��9���b��l�����A�'�F$��Q�M@��M!X�rt��!}��x&֦���6����+V?�띣/�j{��Ѩ`SQ�g�B�<8(�n_C�d��oe�����Jy��b��3C���Օ�ޅ����mc���45�(p�S�r���κ��4��z��VB�>�����r�r��H�Ԃ.M��������Z$��p�3�H"���%nD�x}��sa�:T��ۻ,��<!��j���&�%��tvvu�z��Ĥa{/���G�-%hRi4�9�s������1�'	��k+J�,�ܩ���*�I�+�:��+i�� ���Ͽ�j�?���k�#�p��R��&s�>�.�l~�=#E��M�vk	��g�X���WL��|VzLE���`�ׄ�ce���#&����i�19od�dUԆG���Uڔ{�L ,��F����^����-��coY���+1�
|��6��A��'q����~��������Ay�֖�Q����҉7�=d��`���h}�wz����Je��>�M3��X_��!'\�c��x�N���E�Ɔ(����wJ�N��)��8�t��vH�Ը��U�}���[ٗ�T��h���	GM��(�	�1�X*Ze!����[[s�i�
�QV.9���?iʂ�� O*��[:|��=DE1���
�	���!��Ϣ>�ۣՂ�+�º��ӛ������v���B�n�u}�%�?`�Xֻq�����i�P	�c���ս<V�܎��ʠ��$x������Od=�S�K���q�Ay�3)89���u��U��?�yO_u	P���;���q�FxeF�N�Ȼ�lb���h����x��I�ܑӇ�KΝ�OW�cU����u6���T��5B/M�V\���e��}��M���i�	}�G;cL�%$0�1��V]X>\�A����o_KP/"�{�ퟎ�%�t�o�mG�9����(v�v/q=t�j[�ˠ�xJlQ��|��ٮ��k�d�9�~�����@��'�/�=�?'S���|gVfo{q���# �d(�H<=��~�V8��u��h�%���Tk��������'����ϑԫ��ň��v�:W�-�}��=~�A�;�aT�"��_��#P#~rdj
;4����FJ���Փ�t)�m�teZ3akl ���'�/�G��;H��}�Ѐ��H���(UF���K>���ŏ.Ԕsu����]1/ž��$[�����A�F�ݳ�����q6F̤����u<�Đ�3`�2_���P��h�3��
 lsõۢۯ���+�f3[1�����x��ČyL���?`�sx�,���$v�erg�l'�$ˈv����[��+D*�6�\�p�KA�c��򯜁�߶�=�S�1�P��w�( �r�K?1Ì�0�o�ū�D�ӟ��}}W�ژG����y������� u�jŻA8���jߙ�NJ���z]�'}����mj�c���颉����s�D&��͎����X/��.=��A]���׶ݳ��w���d�&�c��#�]ȶ�1��<M����o������1�-h&��ۻ�3$���f������2��7��η���pI�9��Zl�E\�����i��KAxp����%��Qw�qE���|*cfZY�k
n``�
^W���@��3�2����&#k����%�Ϩ(����B��KљK���"��B,.n���\娆����c���޹��m1��9ssJ|ͣGZ�������<��N��a���0�.��avz��^#�����ݘ��gdOt'?c��!�H��p��@!@���G��錄ڵb������ۉ��~�l�����Cc��b��
��ӯ쓛��	�v:BqYo�$_���لM���l��'91��u�=[�+���J����{F�(��愂�)�,�Z���/2�(�4�V�	]SX5�f�e����9��EJd�K�S����.���9�*�!�T�:ι}�DX���k�����=��屚!=F]Ї���v|����zv�K ��2D/��� (ة���-���8��yrM��A�r�J7Xʳ���LL*(���ڿ���v9��- �������;�)S?�����/��?�7���q��������"l�@1�� %]�3鷩Xxٙu;�x���>��)��%��l�[.��IQ�E'��������A\	ԗTR쎤 ���ۗ+����\��{����������YZ��5<Sڊ4s�=����^�'���Џ#98f���.|k"VЀ�ZCs��`7zy�"��d2����*��7���ͪR��C����V�I"\�kQ���˩�5L��"�����v^puw��c����&^7�]����.��"\8��o甪u� �������;[�\�cwoeO�{�?�$75aA���q�n4E8���7��u����^�_���Q�$&v�����^.�4�.w������	��B@���ڴf��+�Ϫ0]�9�@�P�
�l�̉�s�ʟ�����n������]���ȕK(�B����>�!�y�w��6!x�8B�{C�,�Z���j��/�W���W-',����"�:��ȼ]쁂*����G�=�{�*�2�?w��b\�3e��^z�#O�o�y���&q�+�%M����gq��W�"]�WW�2P�HF�)��(���1�f�U$X����6��e�Cc#��x��g�������D��*9�����ۼ��ɼlil(qRTrxi�H����<��_7��!�nV�rrT '�Z|#ь<���_�C���V4]���;��Q5�e?A\	��85+ҵ�l�dۊշVp�W���]���ف9����	aX��S�q�	�r���a@@ �#I�;X��ܗ�=Vͣw���r��*��ߑ� ����ܩ����o�ig�*��[�X�5���1�1�I!�Ͻ�*�nt���T��w�u�Kz��T!���G.dͩ�˛�&,T���E��{r.���5��`����1z�l��"wЧ����7g�Iߘ���GC$��̈́�ֵzK�sSG�s3۴�ӧ߯�M��Wn�� �oR2��N�{���&����i�1��L�o=���^i��=@�Z*⎮&P޴���lsK3w���^5uRW@�i�+�hs��|��$]�m���ɂ�>M�"�9�U�U��ֺF�;�p(�*y�!/"B��f���!^0`�m/|9:�W��8i��5�A/��P��l(�rOku)t?���4!�i�HϱiHC
Zc({�sb������F�+čGA�M��y.������}N"�$+��,����:�t����ְ��n��{p��$e@��0eq;���>�j*�F������P� ��A��
��(E�v�+��G���\�?��=n��2�<<4�B��O�N�o%��t�#O)�ޢ^F(������Dd8�=j��s��3����m�c^�6Ͽ�`3��&5]��㫆O��]lqU���M����g��c1@�_�/°�8�5�*�d����M ��0�O\@z�����O$�2�T�V�SΓYKHc䲬����3����=x��6ZN�9�=�ʘ������(�E�R�'�fOE̵�d����\-6Լ���%����6��휀�6�l�ؓ��α�s�GV��7������J}�㯐����Ϛ�=c���S�{:��$���`�|�Y�>v�=� ���ª���ιo�#��n��斫�SBLa��"u�����?N�<��!&C��O��z��dTI�B+��w��W2�jŁ!g-�^}ԫ�
F؛Q
��=���6�K.�0+�*g�;���'�<�f�>�K �7&��!:i�3�K$8G�����(s�I���+��)9h���򯆦��_ ~��&���p'��r��*�g8vn�KR�y6x�j�;�������U�M����.1�nƇ��y�����V뷮�0{x��9撒��rWc2�?m�1B���ۗ��ub�a,� 8���\X �I{\�k#zKU
`���Q�fX�?���o}�^�B���O�@i�sA���MA<���#�W:��=��f���"�mu|r�T䝄���c�{ބn\�*�zE4?����\n�r�5��^m�z������`7�4Dި{g�"���������4����vKy7�FC�N�>s�<ב�*[�H�ɣ�G޻xhXw8�5�naY��ԾŔl��g�fR��{�B*����p]8��vc0�c�I�s�8��%�fG�[⪤6��fi�TJ(?<o�1۷{S���c;S��Z�o��x��2wQd��t��ӏ̯nG�u���E8R3풤�=��ܸ���١�P�n���ц�`i��ԸyfϢà��CxO����ؕT�*�P�D�
NC	|f6ɷ�QR"�
M�`Wg����<����fv���h'}WmMW�Պ����*+�gɐS��B�F��z�}0���v�t����z�o���l��M9��^�����%���������E?����e�g�����6��Z|}�X����3zNQY��vS�a�S������sMGUģ����-������֭������VS똣Mi��A���z	YY6�oPh���Ij@݋���K�����{���{=� 곆	�������fr��;|>�����sm��Q���V����,.	k�ג�%�̩h@��PS?�R���/䀬p_�ؼ%�[�}CԱ�W�N]�)W�"���©��YB�!{��Z �^,:��*㻮W��G��E���LA��<�B��B�ϠUF�WN�NX�z��BUy��]���ƨ\(bբ��T�[�Н�	[��9���[e�cͳ���9=-�FȖ��,C��Iţ�:���qI�g�< ni�L�~�Y�w�y��ʘ�~}��K�R�柁����|�F�y�OU`�aA�fH�A[���	���b���Ծ=���(����m���K��K�g�q~fM���)\�r$
.a������$��ӹyɲ���+M�m=��P.R_U�[�a���v3�է�Fm���T����"x��7����W��&o*���G�zx�o�S�h뽜^8,Ƃ-b�8Y�0�a��H�\;e��lF対��iV�>&��Ÿ��;1���@�?i�+�9���>��#���7h�%-2�[8����SgSk��W���U�Ee��nd�5=B�X䲂Œ�!t�HR�Vab�EI	={X)�-�#<��V�xFC�ڤ=a�E?�X2H��;u��wY���tv����8��!g�˙��Us!���R�OG2U��m�T����u��j�VLƑNX����)/ܧ"��aI���%���^�_ʜRG�1�ʵ�t����=K�"U��h�B�oZ5�6:d���J &-��KF��H�X��ZLY/I%��稱"WA�Ī �G�FQ�I�@z�|�ƔX�üK����>
H!��#��˒�A5�0w� de�?X�:�2v�úueE5��`�R��O���_jFF�Ǐe8��Ԗ�u�b���A���#��z�4ޡZ7"uq��]�l2��#�G�9�W�6d��E�-=�K�TV>��/Ԋn�ܞ��"�#"S���t�����y1��g�k�f�&:��:�H�����h�B��R��w���cg��f|���7?2YQS�\��no7(6z� ��3..R��u�z9g�o�:��Z�<1�|���̱WaGo4�e�P��KN`ro�wC`ɨ��tW�#�J�
T�jC(��
�lH�:݃�uN���L��5GQ/��v���6��{mN�	��EG���;	�ŕ�P���֬TM��U����2Yp	�phiu���Vݩ�GS��Q	�td0"����_����I�xP?d����[��t'�6+E͔�U -��l��2	�ˡ��[�'�'S��了!�}w�/�w�t�����m_��"_����7� 3Y��� !���ʑ�r#P=�~�B�'p��P��/[�	�l��FNM���|)��Y�Uױ�灐�jtr��<@7t+S�Jl2��T�.�z#^}���wsL��O�Z'�8���s�`���<�x�շ羡�UD��V"_~�ʺ:~ӡ��6�I��.�T�'U���\b��b��X�5E��E��ӓ֖xw�jz۵l�0�Á����������,T��TT� m���+@�����E׌2��d��ISW��1>��KKރ*�^��6����h��+V�R�$�p�Q�1d�9�)��)� A)��냁VS���ဇ}��'}��K��^t�g�"t?�w��
�5���#�;��/����Y�@V����{��L�@�NR���u���������W������\�_����y�^��xt��"v�
 �]���/��}��ywl�>*���us��"��f^hi�2�n��5����~%���m��+����;��'.��2 ��^�b�`U�jC{���<��<�<�-�3�ⶵ;I[��u;���C�����Y��e))A2���Li��-<C��ky��b0�9�/Ä)k��vꞱ���'�C� ��YA	�o=��A+h��lK�@"ָaO�j�r�PBg+V�-���? [�w�N�g�� 2c��z�L"��8ӣz<֙B��P����g����#Z=ߩ�]]]�� ��H���K5�&��S�n�g���g���YQ�9ʣն��F��1��tnʰ���.��R��!�\u{��D�KK��-��IЀ5�B�L�������&ʣ2�T���)L2���x�@G��L�?Ϸ�﹐�qXI'tt*-�t��]����wq��*��n��2��d�+��1�%���� �������Â�󼵷@Z`��B���ު����H8�����7t���/eR����T���|�>*��!�W��$�x�@��M��&�4Ҕ痒�[�������g���A'���Ru���2@f�g����^�#dSðS�%W�am�<�
n������ m��b?��|�]�_���{��=���e�����I�V[;��W�8�D��&�e�[-���T�Css���y��G��>6���G�I�B]�]�������/�n��~��Y�¢�h�E�7y� �'Js>���}{U>xٓ-B[*�>�6Z
���D��L��`9�K8�8��&%�Kv���{H�2�l B=3>@.
�M��?ww���. }�I0Y���Ń������Xv~y��l��Ez�j� �9��1-_��ش���K�_��p洯nd�2�#&ί��k��S����ps/�`P��ϩ�E
�\u��3��4�<W����I��gڌ��JU���*!6U�r�K���;t�[T� �]�A%3d(���:���7�w�6{�	Ts�82ݟ�^��7"?�G������X�]p�U�P�<�
؃������2|䘶���k���A�������#Y���ӓ��'�h��ʶGX�g�hHi���d�T��q�(R�W��@W���w�}��?X@��s����bǎ4����vk�է(4	�3����>��/!��O)C�w?���^)�pv9�QT��X�Vg:����H�agqW�UC���)��$�=������R��IE�L��E'���8B��	�D��LjF����1���?-o��>�a�]���"-c� Q��&a7a�,9�H������E=���I� ���͹G�Qc=?���ߙ��O���E�=�Jb�29����h�-,3��<�6�N@!0�Wa�OJuo�5l�d%]��n4��C������|��w�B�8�@�29�mDN\;�������3'�H�*S	�		���d!�2��rk;'�F���!`�/-����^,ϟE@���
�"��[�7+���[%@:/��)L��0s�O�ݧ�,)�b��z�r� ����vi��A�f��Ɨ��ᶉ�\�p����� +Gӵ���9���J� g����X�i%T/��.ɘ���(�?�����f��n��������ao����OJ��B��.��%;yG%�1ٳ�c�k(%$�:$ی}��6D��}7�R��Xg��o�?���|�����������u���:�\#i*WlW�W�ΐ=�Kp��K��:�A+�k�2O�`��Ce�9�_wl�]L
̥^��on��q�f)��J���ԑ)@Od��c��}z�S�F=͑�X���r��s�@m /Ņ�2����ъa�1�F�(�$�V_*�SH������U�987T��A�7�ʋ �5ٽ��K�(*�3%!.��w�d�������ꆝv�����MO�Q�`��Bb�i�M#M����ktfۏke�b�	􄸷�3����=-���i��^u)������_���ǟ�����_��p�ݲ,1ЀM6B���嶱v���gG���^�,��<����`L�3�Y��%��ÎO^>|�K��'�s(�P�������HA,��qZ�-�|m��"�K�b}�\ �M�����	�V�����Ϗ@�A��~���Fn�y<����t���Dk��&bz�$	���!�X��Yi-FZ��R�a���J�
ms���noyt�At��L������,��V�߃������֖_��zv��-9t�g>�<�cr�x�t?R���J�,Ò7l��a �a�c��
�aN�3�0��
��_�j"�V��s�j���D�av�F�J�#;�����n�Rn��k��{���\�� ]��Tζ��W-�w����.}�(�u���6x�,��`�U���w��_�>�$���ΛtD�S����~�t�Y�G�uKԍC��<�uW��d�,]��\��Ϲl�b�������s^$���@�7+�:uMM��f^ߛi�7��1s�_�_�;�Uu�����gb��� /#qyS#ϴj���:����ZS������0���L��L^����Ҩi�YC�n��l�Z���\�nz��އ������,G�^�n�ؒW�0�lC���Ք�c�^��v0��$Ǖ�{6�^��o��F+���xǵ_���A���� ��_΄ e�=O1]�w[��y�QC�O�l�&�_0,)��`Zm�97cW	���o�4�����c�V��L;��_�7��͸{T���f1��?h��<��S���)�WeI!ۢ3+D�R�61�ѷ+����7�/�,����)���'�;�� ����̕P��z�����_s��mY)ȭj={7��Wߣ�N{�����a��'�4��OU�ú�6�L��QQ��3��`�z���`��"�-r����k:�8
F��c�.L�O^*X��u�f�8O�b�[fǓ�r�^Lb2|�ogLx��VIڀ%;��<�rN3�"P���m��O� �x�ZQ��);<OѦ��H�<���S��]�>W���fQ�r�`^�=��N���|Ԁx�ς%V\���cM����'�K�ݢ��f��,����S��t��B�>p�ǻm���~�S]-;&W���DgeЧd&yt^?��������"�g7	�W1��{���z�F$ai��H3����
c351���\�f�������H��þM������kM]�G��Mj�v�Kb�G��8�Zo̻�a���".�U2���yw�MF�Y��^�o�;3�����偛e���bJQAyY���&/M��?�s�؟-�k�S�j�}�r$M�����r�W�p����Q9��}�HM����=�z� LD��*�-��`o?����2����<-MV�{�������z���A�u���I6=yw�z���)�� F3O�(�&||�/)P&�����j���F���,��+�L��}���}�hP�yO� ���d�d�qDo��  ɾ�m�&7ӑI�%.�S�������8m�vN뗨%�./�VT;!��b:�ӻ-fM;c��ȑʜ�ͼ�Ѡ�]�b���pyA��,�����g������ii��L����Δ�p$�?�t8A!���fyw�Lz�����y��Ȼ��H�P��� ��s�J��¿�)�@��ğQ2�MݘZ¶ފ,s`�=g�5��"�� c�*�:��*I���"\A�--,T	����c�L�f>���*9;������Ҹ�y��,N�̷2�� B����)�,N���~S���4�����ʳc�v޶��,t��� N�������U����mjz����ޮ9��[����$�����c���އ�;�4��9���&b��gHf����o���N/�p�Ҿ��i͹�.n�������ԫ<�v������F����&nT�bl�����'G�kQ�϶XW NT
������ެ�'b���\L
�TƄ��X�~�<X�qr���v�����Q�Ą���F<��& *��/S�AMJ���0&٤�k,�T%����cW	�8�&����QU��m�<�85@!�������.�.���D�&<A���~4��I:��˶z�oA�)��>wo�	�r����({SeI͓�>v|U�*�ýa�O��]37w`;���i�������?o� �+@;�îo\��#���*{�}�����f���L�^Gz���-��I7�Q���=p�
#{r�~U��4Ihr��\���^�~�u��Ʌ��w���u~~_�Q�s(���}��M^R��-6?j�\8��8Kƭ@���>:�UeG{:6譙��(.����2Oo�9Ø� �_�`��s�z+g噑�����e��&yQ�c��M����� ��XO%�z��t�ɭ1�E����}S1U��Akd"�������U~7�?��R� _s���n*z�Dא]����si��Z�eZ�y�@�����������e*�/zȉu@;�<��Jh����>u;�ཷ���Ӕ�A��x��rי O��E8�S�z�5��ϱ�K��[��5����p���X�b�}غ���{��5V0�ݎ��sF����u~_��r�eN�h���F��vW�#�d�Ŏ�_>��B��� -���޳.��k�0.&�(q�5��oQα�/����A1�����.Tğ[O��Ĭj|�F?֝����^�?�_��ۖ�<�-���ƫ�%�;k�P%�0�V��9e��"��T�L�8ƴ�4�S�yz�8���!��9oȷS��Ci$�6��{F{��n?�Dy6�A�I�5���"�3��!9m�s$.g����"���-O�1S_��1  �ɼ�+8��|��ѿ��@5�nX̛�NS���p�A�j�7�n��&U��K[�IN��z����[7S��Ÿ��f
wxj���&�W���ɵ����=���~W��B��L`qW�1�u^��̸g*���;���L���N��e����!�~�������e�\%㎼���nv�|�+�_��܁�2KVje~rܮ�-��k���c�O���i0ip�?-~��i  <��97�S�n�����1�tJMƴ0A����؛��6��%�0H��C}�#��f�0M�r�?�n�ؙ�sě}���J�c�����+��b;1� �{?����� g�VF(�<�Xި�&���%�-?�.J�	3 ĸ��vh���z슌X�W�y[�ϪR���U� g�]|����fA��	�.�z6�e[�l=Sa��<���e���3����W�'��$�ׯľRs�D]j�>k#2Zk�T����}�� ���\��3~w��[F��Go��)V��[d1�oo2d��ĈptXr��I�� �$���.�^��{���`z��ڸ*�ePբ_��l�~�x	r�7���h�������� f@&f��i��(>�ĸ�&`�b��ը��lT�cN���yx3��h�A*ǹ�_����I�ݖ����	1�{��01f����t�V%�p���n���\痋���h��[�F<�ty��M7�x-@J/ܼ�{hbUr���o<,����Z2��H2%t
�CeK�7Qw��]��~��&�q­���>C�L��R�|�Y?��{���b�돋���٘�5��>V^/�͑��i�G��M��]���ظ�:�����WoԺ�m@��	�e\^����Kz�܉oɞ��{{K����c�P�9���\���ȉ5�����lb0��GE:j`��?i5+�^��9��wd0)K
��~�&'q>�o��y��F� �_n~�!���M���ה�f���>p&Q狗��P��Mj|T|�?߯n�'�?I;�n��s�f,�ٕິ�Dj�~;?;7�C��*8u>�E��D�����=�B�:O� ��u	Y��H����OuO<NI����҄c�e@;��Ϭdߢ�D�'vrk|nڬo�v��O��^��$!l06FR5�����"#Mȁ�� c?b���	�;�#E��x�=(aa㑤Pqqi�����ȼ,M[^���$҄zU�Q7�Հو38��1�=�4�x��	q:W��ieD�a���εU�/�{����W��N+ߖj-?�ҁ�ؿ6�"�;V����U?��dWvt�
L�1�I�)B�����8r�_�ȬA����mzg]]]/9��O���_���]��Pa��V�ƨ_v�O��ɗE�2�7m��7R�0#�؊���F3 �?*�g�����Z���-��ˬ��l����9�����!9�ӛ�g.����Ο���;a^���G)�'D�@)L"��?��0�=�.1c��G�vԕʾ�� ��Ƈۖ�b|~��6=R5�}��K�;��43:�M�ۏd�����s7Y. @t�Q�y��u��goe+
;5M�X�$әZ�0���B��V�z��-����;fR�<\��3�Y�`ͭHT�����Sr\5�t��+�<�KԸ4�>��I2-��z�9\l�H�tz����Ѿ#�Z�j��[A���1��j}[Jc�LT���į9��w<�/B"6���[������Q��m�6u���X�d
��������4�ٟ�L	��)�l�6S���y�ޑ����zɑi�NR���罏�+�Z~D�.zE�R7j��n��I�~s��g�EcU��a��K Q\{31*�1��&�Ɂe|�{�	��Z���j���^��@4 ��d���1T��0kwD�1�\G�h�v�*�,����O`�t_��9�T�d�8�X�]w e+Nai��p;���wE6iw��O��h�:F��p*lU���"�}?��X^]�s�~`�M��߆c|����:�UMV�`n�.>�y�~3��dB=�'����<���� g�-Q��'J��u��{�ؐ?�Cg=����v';׍�B�j�H���(�i�E��[#8?E���O�Z��9�Fc�t��y�Pa6�1T�_z�׏�/=:t�8�|?Q�57L��P��y�pR�3LN���T�E��B��ş�]FO-g�6#~Tܨ��tF\�t;GuC��h��"$=�5��6��SSO%�"-��t���N/K��Q*Pk�V,E��=xaÖ9"��t�vΒ]�G�n�c�c��]��X+O���P�i��34r�j�}[�M�Vp��2-Zz
�w�*�h`V<݃6rT>�y%���7鈁i�g��r��lM8��������)�r���8j���-��7��V����j��m�V`�G0���W��@���*��=|��ތ�x���j&a�IM��PnW��wQ�CꖊC-�\~���'���~*��1Z�j���&L��1�vS�� �v�~q��)/����nm� ]ǌ��p��4bW���n�m�#�?��d�'WURkdm���TS�
?E3�h�] �D%h���ܽu������
Ʉ'�OϽ5�$-��ob��~�`���Ǉ�aL�J������=��?ˋs��������uwyr(��J��C�l�)h:�k<�Q���P>FbK�^���ƩI���A���-R�Z�n�x-�s̎
���]�	"j��t�2�� q��N/ �|�����#y��mi~���>�	\��UvG6?�˛����9 ��1��v[������C�,�5�L��W��'A����+���hn��}�G/ʮ~�>��'���q�1_�YR��Fk��   V��mD�1�!Ş)�Ũs+\�z�YY(����Oп�a�{'`�Q ��m�7s�#�����T��:�̣]w�$I��>�کv̈I���p��T||Z��h{S���@���R�$�3W26p<�>��[
�x����q�a�t���.æA�T������^Ml�����|b��&����jTOKe�r1��o�
�^�vŎ_��߆&�,��"�n����)�`�~�y�<��"������ڒ���!���ꬹ�4���#��W����Q=���+Mn��$�O0�o�]}e�]2.'� ?ggg�n}C�8��W���X�Y�!����W5�L",����!�� |�٣�KN�T��ѩ��6����؉��N��+��G ��v**G32��f��׮����8Ώ����i���&~�^��;��vE�7��ZI�t�3a۴��HP�!f�σc�ʐ{�У��F�M���������t�u��[1H9�!�O�& �4�`��}���?����I)��Bp7�Yʢ���#�ת��؉V�t�Y���G��w�e�%׈��u��[���
}��k*~�0jķ���Zw��V �b,;�7s@���磿2�-��)@�����⚪֤ޏy�M��$ªg~b����\|8�K^vC�� 3�w
)I% -SԹ\D�Ŕx�O� ���P��Rn(�������h�sg	w��\�V�F:�QT�HB;��NNHo�}�Z&�M��[ �d�p�����N1����%��o���VBe�g��R�C��<\�y���D�(�Y��}|�+ֆ�Yݷ>_.�m�'k��vՌ*�+�.��t�{�nZ�G���?3x'}�U[���L�E��5H�Drr�2�����@���X�zy��6�<��ל4S94�I��9�=����#`sPض����@��K��)�ئQ'��	�§�N��6>��[���`}ѱ����^�V�����6����Q@���o��7��y�rk�
y�r�9`���,�=� �c�{}�3BJmp��;MPvIy"�I���Z%�7���"�L�[��6�]=<ț��R\s3�@m�����$��Ag�}�]��>��Hd�}�6���� ٟ�<}&����.�xYJ�_{k�!��Ӌ��31�׹k�g	���o����E�D 5��[0G�Θ��l�S�h;�\�VeƈL�K�����N��yP���{�,=0�gK����, QE��(��[=�����]��0���7x%�,FTT\=�@>>��\.H�)�Cp}=%' �����h�ľ����"[]��G���Z�}�,M[!J0�&"�5�4-g
�/���z
�˞B��� �I��ɕ"$NŁ�ʃ����\fnz^�v�嫙�oΫv���}�٩(�s�P2^�ٿ2����{��ջ���o��|8{٩#z�ŋ��������I�^���X�d$�+�h�F^+g/4��^pF���j|�����X!
U�?��-	��LZ<yM(��*��e`������Ķ�)`�:+�'-�V���mMLL��=<<neU�4���]$�d:9}^{Sl�DPZy3� o��/�+�~�	p�:��4�Y�]Su��r�ys���I8Y�i�fQ��\�`)r��C-X�=U��;�7|O���M��$ ���>hfO��2��E� ��U�/-3sT���_����V:fw9���ٝ(���x"�"�1�'��n� R����~��I�[~=(������cff���1P^ڻi�8��7FY�^g�(�m�F��dĈ��D���K�߁�qTd:�s�&x����u"ؼ'�U�����ws�x�t�'����A��0RtG���Ɛ%�������J�6�[t��t��>�
��D�~���H���i�g��gg�u��F�������A.�ZT��ӿ���(��
�e�>)k���V�n4L�W�{�hk]a���NA�겆���uh����%F_�0��:,���4ޛ��o�,�r.6	Lqz�y�ީ� �!Y��sUOe�s25=������P��-M�+�\N�����������n��}��?p����iC�d1�����d�t�	����B@�|��m#uuu���?N�窿ƻ�qƋ@��z����&0|E=� �l�������X����ͷ7X3~�U�M~W�\����yn�4׆��LI�!Z=��e�9
*<��E�P�z{�yF�ز�(���/A� 21�	���&���N�c�0���K��eML(����������y�*�%�����dT����1�B(�� �5}�p�-�e�A�`[�c寅����at��C�kjk=�&���UU��L����b8�g���@r�K�o�{��몯�>D�YH�'<(�q�=����^~M������U��E�/�g�<�h���ݙ�ܴ[
�BS�\V���\��s�IO��}�����^��ع����k<�o&JѴ�����U���U������~�qO5��-�`¡�B�(Y�g"�e���x�X�\�iz��Tp�>+@1�`�3���Y��Ƴ��j�h�Q�s[G �oJB��z���n�����yA>u���?ƌ���t/�l|���9`��z�JPI�w�x�󍪢>�K��)����Ѿs5�/L^:�~g���ݞC,t���5o�(�.�h���$$��� �����Ì�"��yT0�ٽjF)ȰK;��D��T�!* 7�q��R@��KG9/^,KII9Iv�r�6�<c��#�f-y�Y�W]% qб1C�\c�:}zls�����gf�;t|��z���^^^�,�tȌ�����h��@}ȃ��>�wۉq�����7��)����=�Y_��h����F��׶����yz���ـ���ɀ��B�dOUT�[yRH���v�Q�Ea���N{9؟���#6��e����6|�2 �S�z��T3j+t���塟m��Pq6S;:@�ΣU�GS�Ffn�
��-<2�LR��'��T��w��詩��Q�Z۫J�	��(�����������*M$n��cjϽ�G_�gh����Q�5;����bO�C�y�#�t�臡�+���^Jy�(����$��������_\{�v�$�����U/hb7�}�|x���2�������'1?���f����uDJͰϗ���fUˤ7�&峣=+��N�R��!c�{���xē1ğ�5���i��ѧ�nC��z�mgŇy�����5�v��tI����Ww$��_����)���t��?��^�0�T�9��kc�ӄ�l��|���g̦�� l�قA�>�����x�}`�s���������AJj��ȳ�v��n)daxz`��4MwW�r����$�n�[&@r��a��7��
���� ���9��&d��B)�M��ɾ�8�ώ	C�ZS)cc\7ve�ןg��q��7�.vv������򷗖��k��e�!E�Ω߹�s�j����g��kHEhP�aX�k�-��&w��?
>:�	�<�m컷�wJ�Q�ݨ��ny��kך�LM����nn�@&$p5?�͛U��(��@
<B����vy���\�nπh��ji��lE Qi0�0Dy�4��V��D��ρ�ٞO��0� V�pQ�~��h�����X��? �����/eo1�w��!�6^+��k
ս+6��N�d)�aMr��M
�X�޹�h�2=C�i;��Z��p z��vI2H�{��uO�\��!S�|���0�옃߯��w��H���8*�h�|�6~�X\���GE��aT}�Cu-Pͅ��JV�a��f�6���kb|F��Hʬ�>�iG,	ڤX�'=��Y5�&8�Pzm[2l�;ܶ�NF���2�a\s��~z�y�B�|.TV־���P�X���P��XAS7��>�n �vNx~�a��ݠ��y�X'<�02�A���A�p0������ey�)Q�|E�W^���ATޡ���has��n�r�TŐD�X�1Ec���k�j6�Vq����SCL�\=Yt���h�y��y5C'��X��g
���-m?2]�������Ct�6�SGyB�	q����O޷H�a����%� �W�A� �/\(��bA�Vh�eʃ���I�z��ax1i.��k�kۍ�nh��'J9�O�]0�?�q�ٴ�+)sy����*��ƹ��w�j"��ȉ�����1Nx	��/�)�
���jVr;jɋ���%KȂk(cB֠]������G w�q�����$�m�ݜ�����Ъ��Y�S_�!��Ň�G�{��P�NŜffA+��@�L�`��8zr���,�3�����O�����w2	�I[d��3E��)�D� |A��|�٨T�א��kp�>P)�3
U3���dg�m12�d�o�z�dG��k���ő��㟉W�C=>�IX �����M`�ǆE�R�
������,T��f,�ؙ
&׬�cFH���̶&��G5

�j���/� ������z��ޝ�ü�)��vv�P���Ȏn��`�����ߐ��+t黱B���eI�e�D���<��=[5z..9�L�A,��G�[���$x�:;�a���M�`R�:b-[��Lt��W�u4b��L�:�\vz���o�=9A����N���F������="az2hr��k|'��)�?����+�N��*����<r�pM'���;�`�$ҩ̤��a�^T�����bD��|�og���#�����ȡ���N>3|��3Qƽ��'?�l^�*�8�4�� ����9�\�c�8��*ٖ7x���d�����#Jv�M�ȿ�6PD�@%��v�?R~�C���^"d��|����]"���iK�ML<��E����c��A5�����G��vݟ�/2��B���^6��� �,������r��x\1b�M���cVυ�ռ�WM�P<��Q+�m�n=��v�t�� ���~�����|ƍ�����eL���cq7�#UH���~U�m,�㫍��!���M��Y�0	�r�X��7��,�ch��~�;�Hy��A���M��a�B�xWb���ұ�/Q��u^�޳&�I��h��`zG�o�m�7Kx����N3�F�W�����
�$~.)�~�+k�9����c-
��o����ڳ��� �`���2��l��Ğ��=��w]ZYҕ� �$R�{ Tō��;d�����i�]QN���^�L �1���
guqt� ��vm>,}�>�5C���w���9<�]3ܹ��6	��^��z#����kb}4����5\"�\>)���_��04�Y��]ܜZ����
��������-�T�h{���&�c���� 	��)��r.��,Ɍ_`X���p�6}��g1!�p8+�h~q~�Pn��G�e�R$������o�]�؀�U���G�\�z(��� ����L�S��%�s.3����~|�?:Ϭ����/6F�����57�	^q<~���yk�ZM%L��UǉB�v�@y����~c*&��a%�r)l���n�*�UbS&r���;bXc��c''�ba��P�}�W|�߂��a�̀�]���Z�kw�i=�,Pf����?�����=s�\��/���NK�@,yPa��^�I�3��5���r;C�Uכ����bX�Se���R�mv�j�ߛ�[��řSk������Ģ�R{�z��b�dO�]E����5�v>��:M�}.�qP{����0��Ă��Ǥ�% J����� <"
��}U?Y�\�b58��q���Q�C(U��3o�~wW�����慑=���~
��n��_-U�O�H�7sC�E��~șM�qD���	
eF2.��y�p�Jr��/�)���/�+�>�d�A�?QI�
%w��Xy)�:�o$���A��8�s�����6���v�ޞ�u9�:[:�n��̸��c��%
҇��3�M�F�~��8�����	�/R������k��H�bVxr�[[?�@7ϰ�zn,%��{��j�ڈ��j�"/�Tv�o�%����e~BSAu�n<|0V,&�RPd�d�K�=q�����l�l�ئ�|��
�LLh�>~N͞�2��cv�o`̶֙�JCo]��~������Gp����
� �+~�q�Ο�^��V��n�x<~��I��b�<�#;���5�6))�h㞼�aV�C̾X����f����C�ׯ_M!�/�K����y��pԐ�S0�?�Q	���/A@��J�	BN���{:�<5����*����+�K򍿹x�pag����o[5�
r|���rS��>/�q�������@�H���c�q<Z����'���ǯ���yo���R]E��>�<�\�p�6?z[���T��!%Ssk����5m������	�5I�zhn���Urr���9����J)u��a�z���iG��D>i��,����s�ߺI��`�x��/K�))��;��ID����D����m��|�4Y��={?��?r=洸�(�Z�!�V�аp���Z���i���nw�`�p�����O��(d�g�"jd5�;�_�84�08�a{ol�
%e�8��Uw�Ƥ�Y��;���7�6�m���O���͍LG-l%;Kuk}T�+��
��Ɨ:�.��N9����]�ƀJ���������D��-�:S�=��FF��K�w��`(b�^��Z�;��;2��fB�#��:D�i��p��nU]Zz��S 
���bbb�MU� �S�\ۛ��B�J��lXnk��^ y��,9&j���9 ���@U4H���u�|�p�<Wʣ���AW��=h+_-�bov�P���c!���7��������z�ˎ�L�ۘ5�^	j	�/�����k��c�f.��N�O8R��kΥt�I�֨ۑ�g�A��M?Ɲ.i�I�?�ň�A�a�.���t^�����%��t�az���B-h	�C����_U�Tu*)cv�v�Zḋ'�~wNu�ݖ���*�dk�-�7g��Ԡ� ��h�ۀ[⇗�R�r�5�(y�c�lk�������K�]vo$����n(�S�&qRSe꩝��:�ȡm�<G�2Lk�w�_���WUTTƟd�*�FM/���6���'7 ��G�\`7*���Qg��҂b��V�a�4�p� �=۱�J��QW��-�-�s�9����T=�Z�ݵ읝���M��*-��p����A��Uz[���Aנ��4$n���:�,呋Yٍ�Թf�oO��QČN��Ի��(|#8g�ylUVh����ƚV�T�!}t����n��]��Op�����gee��%������!����~��>���n-����%��0�������	�<�X1�z|	9��}���Cq	����lq�k�M��9���#ʮ�įCH"���.�>u�����`��EV���SH���p����m���2���&�ƫ��L�e�c)��]��+Q��2k�}����������.I�L������^�~FXXG7�,����k͈��p��h��i����l;��s���\���B^�&~�?�"����?|�"���+W�"b�¨���s
�j72d� .���g�F�/x�W�+�#d�٣����Q���ю�9���iJ��\8�o��	}�fjH�>��A6���J}p#p�>�y<z�5Z �if����a��DI���x��ʘ\�f�t��3ߥ������B���3�O�3����W|(���^ipG�t�T�|y,eK��=�PE�^h�]/$�&F2��@����s$�Ӄ-�\�/�W�-*�=$g,�f��
-Ɗ��P����D��T�sDZ�ax�C�L'�7����ʞ^y'�}`�돑�.�}�j��i?��
�8'����D��a��'k�|��tGVvy�E ם�ƶY �`L����I(�ь�P���Q �v�_�&�-�j&��רapb[���~��D~���}V��N�@w�0�z�8��Uhm�o@QW�l�Hm��q���?�F��#��'Qp��Z<(�p���z��^	We�w�.B�~��9�V�8�T�w_v�Xﻹ􌈕5�.���6g���~�P
��sK��F�-�>��ρ��~��t��֏/H��� o�Cw䴦�T{f}�@.3�m������h��Ғ^E��DV�o-cbJ�k<ږg@�x���`ƍ�}i���˪խ�6jЁ}�(��\a/,��p��鷛�����z�\g�z�y�o�Ӈ��~ !B��g���r$�qyˠ��M�@���xf I�����39���͍�/����	�R�@�� ������s�Bb%
�T��An�OV��u��J �Mx�|j,����AE�aU�,wuv��M0����5��6��A�]�8�h����Q�W��ey�f`�m1��GA(�o�=���N�(ڪ����i�< ����s�z�ss��1��x	���������5� �_���vc	�'cd"�E䋿�1���>$9k�H��U�����R|�*5hi��Z,���p���ަq"(�f����p)���i�����X3���a}�j�D��R�ӆ�Ө�\��Ɨn2�!6�2Z�/2�rh+����<֍�bs�
��5�}8���ӍB���9�����ڱ&�B;D��}
K~2{����i�y������hZW��1cT:t ���2�*�s]���g������O���'PJ��"*�k�v++������0�P#MMM}2�����x�L$�{�s�����5$J�q�%&LZ�08��yb��8-qw(����16��/�W��(���a_2y�'�RҌ����0���Ws6�r���5���ncz�O#+�KH1g�+z��H(���W"�7{ngJ���?(y�- 6�t0u7@��F^��{���P���o�Alw3Z�T�~��n���C�*	�4��4 ���[��u���j��=E�m�9e�T�aT>k��z��7�}�(9T(���&^v���z	��׭�~oz5!9�����*CG����>rV��1>0/�ի�E���D�P8"g����_��1�:}���ݻYOD9nף�!%В�-|�(h&�ٯ}�E�3퉭����������˷�����չa �{a�B�+L ���V����H<�o1@N�&6;%J��U�̃�����t�?�/���'ZKJ����7��M�8��s)���
3�Eu��f���Ń�2�	����8��@��)I"\����ڝ�s՘+k�ZC��Uƣx-���{7��D�-�H6F� ��]9�n/���ވP��ZbFI�����$�~�I�=Jx%8��S�>-�CLn�D�nd�^���Q;�L�X�v�W�5�3��w�oy���)��H4 �i�~�6�a>�
:Iz�AXv�.�qw`W�G/�)QW-X} Q6���oEC�����n�iff���J�~���|k��\8y���Y��L2�z���wD��V��D��/�> 2���y��tXW�q[g��i��E�bJ������P,��[Rmʴ��A�a#�i�CQQ��rI/x���p����ST��}1 𧨧��Cܗ��.����{���ԏ�}}��>��a�?!P���{;4����p�F]L���w%w-h���{��`?"##p��ǟ�$�6�d�d-�$�ppH�\���yH����X�~-L�|�94��DsOO�:T޲	$@Rԋ��믨K��=�#� �L��S7I�_E�5����#)�������1���%6����
iy�B��Aȹ!)+{i�QSi�{-� �[)g���x~5y����H2�M�=�%F�F�.�ǜH����P3+�_���EH�$�-�鲩�B���f�P��HG�xwk?>74v(�RgA�q��C�@s��\��%_�ӿ��\o8b����������#��HEi�c.��;W��R�;wg�w���<��(���-.a����+Z�X'�ď�w������Q�e`>o��VG���@�d�o�7�2��к�?)ciFQM~J��yQ�� _�=ӌ�H�4�%��N�u����V�J(�3洷yth��p�;�s�-��FY��{��}��)�W�E:���\�]���jx*[�� N�����u��ԟ�@�n&��}ȝ޹������&yH��z�Z�����)�M���e}��|���q�e	1�X�+��Mb��^�<�8_%
��K�����
�uL�7l�p$�� <RrG�䫆�nUS�Mm���6�!c�c�mk�o% ;�y���O��-	�o�:e)�������7�����(�Lh�/����'}�0�h#�̇��*.%�-_b��-1,>���[L|ì��>e����Iס�E�F�[�3z�+㮹څ�v���p5RR7M yN�c+��H逅X\%��c/	��h7�a��wU]�#��F0��^LެA�����t�|�/�տ����ᄌ2�šf��Sм[K�h��r�dA����^1@�J�F �4tˈ8�ძ)�n����v�"��tr�4\�6i����B��K���œj`��g����v�!�ߴu�E��j8���l���C��K�=�PU�����c@	��3���+C^+!�<�}��ٜ�D���%�7�ON�hLكg�T*�;�MOMI�%!+���?.��Q��J ���R�Bw�(Y�Ĺ?�-�r�<��k�#��o��f�ع0cȾ �S�K��³�y����6�̑P��5���z���KX�	�zH����;�+&��,�_\z��.�R~�l���,�_yH�|�����4Ld�	�X�J� �jM�����X2�dx���`7=r�<p{k��;b�&�H�G�G.�/�\���k����ƛ�$IӴ<s��Tyc-=��/\��~��g�ʌl��K�Ӧ����(�5oB�^cL5�r���ǀ����+����Yz&�����#��|��a��@��?fuYE[���J��ؑ�ګ�L�5K[{ob��EK�BlboB"�����|�����"ו����\�q��.�Z-�W���LQ�[�,��>~r^̣����Xw�Dj�g�\�6B�����
9`֚D���K���ۡh?{���gx���r��,͋[��|q�z���"��s�2L�?�}�n],>��)�>�&鱐��7�z�a��r����"�uRꗠ6�����
�4G!p�5{�CD�m���,��ӵ�:��(>�X������GZ?	�iP�C-Q���犆^5�O�i�'�ɽ�PmS`�?�&�h�ٷ�ӱ�cx���F5!9-Ox�[#�ޓ�2�k��i��9 ���\���f�^i�F��0=.�~�l? ab�k$ �'3`��S텼�2����.�c���g��W8�}N�.�"1&I��h0LU%?�VK�^Ɯv�h��<�Y�2��]ﰣ&(��E	6��i�4<�G6���z|���0�b��B�f�6n3��`��|��KU8ը�	c���H�gF�^��1.���5|�%a�����E�N��=K}�a��VD}���Z�)D^ P51X]n�P4i������AȄx@�=�eqi��k4®f�"�P�C)��ΏE��$�%
L�U�}�z�Af����{��:��amQ"�=�VS�Ov��{\ױH2
��R�0�K$hM�	L���.P���{��p���C�ɘ��f%޻�c�{cC����C7�)7���C��<������;_�X���b&Kۏ���MSҠ��F&
�捥B����rk�|mt��^��>��x�?O�0x~�=��!�_j8�*X�f(#mA�����c��=.q��Yv+_f�e�����=��Z˾�u6_�&���3 ��M]'��N@�K��.E�[	�&�$Eu�2�2���R�J-7l�7��a��r̅3��\���N�y��w�y��o5�hn�S\�<�$����Ѽ�s�/�I�]T4�����|HM�ݤ��R._�2\\-�<䛐_�/䗃�{#��v��E}�j��ߐ�|��.�C��f9Jq}&LF��C�; #@���<۟������uO�}Yc�µ��rH��w�����To�o�@�(�`�#�lΕx��a����d{w�M?k�4�>Z벪�����0��rXn�?��Ee<*�k�u&臅䓫�T����7�Z������k���O�����Qɱ�n#*9[)V���3A$�]g�/���Yc�����G�3QA�G�#@F#���=�N8%_��1�k�/٪6���#��IH�y��'B�X&`h��K���m�m6!����5�O��|�w� it$��|��o�����A���:ﳗ��.�s`]��̷���hE�\;b��P=��1(z˞���-FO6�?�"�{c��������D*���.]646fL�-�x�M�ˇ;v��~��uz�ZA���8
��6��cE�kD�p
vV�q��H�$�!�'z�R�?6jRω)�,��1K�z�1�z��}�7��lֆ8�A��N&|*�m(w��X"ͣ�/Tlؕ5)��u����I�ƨ`ǵ!lȤk�Ž`�c�vU���o'�q���j�8V[��4�|�5)�zۣR E�ċe�~]�7�8NcB�iw_^��l��p�֧��Y�żv�pB�vuN('4�����90�H��]8l�;�
A#�o�{��A��4�js~��nq���K�"������Q�J2��}�!.GTF~7 �L�P槻Y��go?",q�`k3L�g7b��� �D�q_�x�V%:�oD�6��:�B3 kI����Q �K��B_Rڦl�;V�O�ةB����=�h_.�3�=$������n���Y/�ދ�,sW��E�3�6(��RP�ʟ��Q;�@��$���K|���X(C�����7v�|����C o�m��S���[�zWl�����CUEn�l�i�F�_�'wk��;�)~jjE���]��}UpU��vN�>�w�����H����(Xn5f^�[ԩC�-�z���h�:ܡnU��8/��{b�vs��T�ҭ�9(HJ����$xGѡ`�@1��<��-�&O�B�F��������q�����y�(+�vK��+D��J��U<Y��DBN?�&v��55���/F���!c���� ��Ec�M�iDS����<Qrh�Z��a������GO]W�~]�S��m|���,�^P�o�U�G�g�Ʌ���<?�������5��n� f)�7Q��1C<Q�f�0��t��-�^�6�ނ'k6GSfk��gz-o�5[D��U̲b|Ф4r)�3���{�R	�/��ܸ��w��r�B`��;=�p(�6�	�ޣcTLY�ku�2Z�_�<��=��h�׵~���ha��de�5d�B\\1��GI`vεeQ�󏩨o��x��!poI��1@��]b��^3��8a��4x��Z�����L-�ue����EU�������6i*rtndq���q�`w{?���̇l#�>��bAQ�7r|�vԟ�����8t�����i *���up�W�^�w/~�hp;�s�����E��D�<�Wl�w�����;\>��i�.qE�Ĝz�K���)����O&�Ӥ�:�|-2���e[�ޠ9�2�1�g�����"a�ޠ�2u%�Ύ�!�r���sj��0��^^��@<�R���|Z�y
��������\��s��R:�|��Ռj�Cd��l��d\,%j�u�x
_�$=�s[�Y�g�2W%���M�"���]zl��Ps35«*s/Y-��j'bTYF;�����:��7����j��@��K�:��A#y�;��B[B�W�;7'�5L>`��Am[�q�7�'�w���f�7��gAF��jw0�0S���E����P���4Za5|�g��2��Xw��o��� V�����-w.M����8?���g�b���}b��O1�Ǐ�N��K���K���}��~�s5ϫ)��UI�Q]���u ��1����n��[�6�.ܚ\~�j�Z�8�*r�<��g� B�>��A�.7�!>KÏN�$
��G������}��H-DV�G�J�4=�S�nY{�>���ﳧ����'M�a􆰷�^C�d_��%�W ��\�b�O���Xl�d�ޘ{���. ���d�c�Q#)^a�ibd�������7ɽi?Ԧ�C�@����9�@�h�x�O�s��J\��K_�ƍa�C���/zi���z����c�ө����WVW+>|���ie����mG����-
)ge�vH��H�2&&d��5�S���*#�ER���1T�e���h���+�Q�� #	甝WE�=���G&<����_u�I�{�t0Oo����!#�6ZcD����վ�����Q�^1��E}�W�1����:U�e
h�c�º�Ӎ��ueu���wZ᭦�S����$���3O��Y-��T9S?�[îak� ێV��Dv��e6Wʭ��;����k�˒B�3��6����$.wݽ#Qu��S4���$75��r�{����U�:_+&E��(����f~̸ۀ�ww���Z�΢�VW�����n��;����yyN�ڷ������`5%Y��W&���%�fj{�eA�O�ʇؚXtZ�-�Y4�d�WkV��8x���Z�Jm�mS����y���@U�٠�Kw�O���/qEJ�a4Z@�hs�l��h �<�yJ����K"��Bw�)��I�֖�f�ۊ��z���Q��$&��-��L�r�S{j���ZR��X9q��n"&�qGKP�������#���r<�H���,�j$��ׅ(j��.�U�8k�E MN$H���߅`n��ma�-ʼ熔F�3k.��wx���\de�)ڝ�ȎXf���/�L��$sz��S�pV�k�¬�qc���N�:b�l�����<���ݘ?�(h�u��s�`��������{FWI� ����+c��zHL���XG��F��<C�R�ȵ3h[Iϋ�_,l<e�4�_�9������-Q:���a||��K$5	��ۂ8u�z�B��xX����鷽�Mt�6���]�=�P�ﳞ��V���`���\��5�}QD��P�����IĞ��f�/���jM���q�i�k�F�����F����G�~�	F`wR�Uy��`�ȔLNZ���'�(�mi���7���y��G�p�����܋Q5¹�!����7�����*�pܿG���8�|8�(#pS*�[�l&��*^"�_� uBh>�R��o�\�w�7�j��+ĝ�Z� �t�g6z&��$�n�q�S�/B�������/�����!=��H��n'+~[g��"LY=���x�D�7��d#܈3l ]j1��R�4jM@0�k��ʍ���d+c(��ﭼ?="����O�:E?T�:���[9�Uv3�;AbE5�����_=R��C��]ЁUש��?K��^T* �WI*�S������__M���5<Yf�N�ŗ	잗4E3՚j���?�{��G�N�q�Τ%��Ɲ��:[	��wo]E�~tQ�������U�/������7�`#1'譜��t����X�՝��8$\d�G[�RK��y��~A��Ҩ�	�M,�4~ �ڰ1��tm,+8d���M�>#.��J��}<���b8���϶��cZ���d�J��jj�c��{�}�1U��A�*�ΝrI������`�n�����i�]Q���p�7���(�Rr���<� O��z<kj���og�?s��`�]_q�V�qqIH̎�5�����J�Nw�h�y�����t
���e�Ct�K���m�����cq)Ѭ��:Y��4���:>��@Vs�#�$�� ��@��obn�ܰ�7<Z�-�b	�au.y��9�`~��NȨ7��I��(��4�k+���r�wP?�����Mz�>����9T�yW����͌��3|�ڨ�b���������C�f�j���s�O�An��(na�P31���6?�M>8�ǵ��������hC��N�`&��t�d�`����|���&A�C*���5�7�k1�<�g<���65�������7�k��[�M����K���ui�ƻ�o��:'xh ҉����H\��絺���2�Q�*�8�U3E��A'�v��ߡ�6��6B�-I���)��9��8�X��q8�������t�;k����l|��7�ohn|y��������R�
�5!OTnm�<E7�c��:�E	�㯜µ��5^�b�U"��7 T�Z(F&�x�Ȋi��ebI>8
�/y���vA��*�	�O��¶�K��0��,�
Ė��M738�6  �`�=�b�[�����9/N� a��Rg^lA?Xt3/sʪ�c��ݿ�e"q5FF?����6:�'3'����:��z-�vf��t�q3��g\ e�w$5�k�8ڮ'��q뱇����Z+��i&l�8���O�$f���|���zl++ѽh~p8��� ���>YΔ����VW���9l�O��4/��
�}NLӤ�Ηn��#s��|d��ƍT��3/�� ���G�X%{�C&��lc�~��y����C]�py|�۴G�6�.ɒ�V+{n���NA�E�
� �`���|�^~8{Z�R��������0��3��R
�A�6���pW-E�'��\�b�~0Ԇ�8�n���Z>Z}4^��p5t����$�q��
�M����U0��J-�aJU�i�9�U��`����p�
�I�������}�v#p[�=z,��iק8����oB�����z߀?�B���ʟ&l���A<.�!�0��w*2t�(=��fj08��y�n4�EAe������$�O��捼�򝨉vb�4���*f�8��!J^��p#��)��'����" x���pe�Ğ��6��O���7�<(��rRTB{��;�a�Ǎw��$�~�X��oa��O냠��O�y���&���ĺ+���ib�E����,y뒧P�����f�e�j;�K5�Z鬴�d���deօg���{�^�Y�T�%�ѻ&����x�*���u�}��n��oSG�
�^'��=&Zs;�Oc8Ӹ�C��F� ��G(�{��f8�7��kxs@h1��wk�i@�5��d{��d�.;���GPص�W��6�� ��4�����R���G�[����ݕk�q�YT-ѥT��F�Y�$���5��ëF��r�i^�s9nsm�T?J�5�1��g�2I3�O�9⪾-A�H\��?��?�	�ؑ&BVO ������L����%�6QSRU����t��zR�:�K}�l�����=0�lnhӠ⋖�:�=/�ȶ�������ˆ[�t��Z/��d��/B?�o�	�̐�@�`�q��*U�BȄ�a���>au�3��d|�-��,�h��(P2�P��(�E��$�KUР��X˪lS��B���װ�H�]['дZ�Y���\0^+�bF��(H�A�7�&Z�Gc�}�t�yɐ�6مi�I�����+�������-?�N�괈�
�Jt�c|-��/p�z��Q.0k�B� ��~i�o8z�6��K�f�#���ۑ�R3-?��5��'/�u��y�V�Ք�<riYu'�ܼ�z%n�o�]�%��Q��%h��~��M��,ۻ�l�v�,z�
�Ū�_x�f�7P*�t��\�#��HA �k�K�����&���		ǳ���f�+I�n�ߟ ��%���dm-���v�����ï*1V�i���`�f��������h��@�޺0 �ٴ�W"�B��,��F���Ij�m���*UH�,6���>n���cAe�魼��B������9_֤T��lI�8� �H����ST�=�n�}��X`*xgQG���̷7i j��O�#]�}-�h�B�HEn��+�?7&����0�3���$�"�;d�O:H�&�|���3J��5K<����qԟ�:� g�/�2Wc�S�sX��NC�=��"�vG!�'��d�"�Gk�}�����XÔN�qe�}NiQ�Q�!+�ѳfH`'_^g$7vh@L0:,cd��^o��_:&���d}�&�S��� =��M�K&�ڠ|�Î��iq�,Ү'G�6�ؼ���7��E�X���H�m��fS���z$}}x�����jZK>z�F\\<Z���:yL������Ja ��i<1<8ɣ��h���-�u5Ё�Dn�	�6�IIr��^!�\!�˟�}���&�5��h��W��\�x��ˤ��A��=i��-��������oed�%�@gZ���*��_���+h����k�+]�y�=��`�ˡ�v�-���P/(֫=�)���o��.�'h��o��<��,a���-�o������#�_��\�ypO�	d
��/N�3P�0Ɣ�]������l>cx�q��2�����r���a��>9�R� �RHh���f�` .<�p����Ǹz��Q(�I�h����QAM��,�\>zN�b�@�v�-wY8 pܒ/XR,;��lx��3,��
~�>���ĥ�f�k��\9\��^���7�n�12ɇܸ����?�vY*��yMy�M=:9�\tc ?�1�d�����>�푝X�fsZiJ�
����ԝ�U���:;�a�嫡�.�09�)�m%�(�tx��?�d���C�CQ�RX\���x[�������\;�f��$��{�Z{�SP�ݸʆ ��|x�\�'�3m7vsT�FTxhJ�-n�%~�a/�\9�_i���if�[�_N��˟�� �W˛���@�}Χ���;����=�pcֆqy�C�1�}�$�aZ��<GC���7Y�ymF:��,x&�$��fj k���%��;�����n�1�b,�`�3*�QE�F^� S��z�H$"�����2>����g���b-����l�"p,z���>֦���:��;:u�Y��r�:��Gvz��#��П�]^Eo��Y��A�O���h��1%�����O�2�)Y�F"���,/@ bm�`����؄�;()�GM<�k۾�Y^6���h�eE6��qV������Ҍ/x��q�@�WGf$���U�h���~�s�4�	`w�����G�`�����p6�&��b�c1`V�h���ϱ[ҙO�^&�9��V�	��ܹ�:p�߬�IÅI��3�hDa�k��BQ"��Z�-o�`W���ԨW���:�?&mTr@Q�okF���w��
l4@fC�g�l�����6��e�i_��0O͸#�d��R�>A12f�q��Ք��R�D�8����䩣�D�J����V���
�CclT@]q!���F{�lđ	��n���֌ri �<�9t�V�B��j_P�nX�� ��ѵY��r��$l\�:�7�=��������+I0��+wl���ۦ��{��j��ҭ�!�0��)r�KvY� _�
�ѽp�ts`� <�]i�v׵������ҫdd�Yn�k��Am��S�2�/���ٯ��߅FysW4��}G�~��3��HŜ�pZ�����vu�/QP�
��@�����:Fi�h>��� ���=�5P�`>u����Y���ft��<zR#�O�2�8tL��y(J��y`����|hO t�6ٜ�V�ٱ�=a��"K@)Q�x���v>S)�^��3Sek"�8��5���R����\�B��{Ò��Pd����7�'���yyۓ�z�[;�Y|~�]�|��8���1��!�
�Ҩ3��MV��lw�^�3��sh[�y����`�'�l�5���؆��#X��-��2;恱��n��RyS�G��ּ�iȸ��u�l��R8���53��v^�Ϟ]y�(��(F����S����]39�Q��t��:Ąmm��� '�<�[�������<���U��v��H�ʼ�����Ν(���|ԭG3��zq55�q$޺Τ�Vg�w���2%�[�@[��Y�h%��uL���^�5k��Z�M��E�懽5K���C����$�b�g��ؾ��M������۱��zM��m���=�/��i|�v��DaJ:%�w�ꨉ�ZM˗�k0���}nޘ�"9���q��h7�1�U;#���|�&.�̘��k��.F�pV/��y�lȽQ���K�Wx�Y��x�櫉o���TY��x�{8M$�ϑ/[%G�u ����n6�d�5�����H�˟�9G�bv)v��]��:֒j��u�2��(�g�{����σ�Y���&�x�1���a��Т4��J�]Mh]>�zgW���hi~�CTh;3L��, '��p�qղ"��*90�SW�jd�Rb��;�#�/322x외]��Q�����Q�ҷq������Խ��ĉ�[<�=��L��U�T�R)�V
L��2~�)���B�و�\�44�(le�@6n��o;�Ub��ew�$��"b�Qjl1�C� �^2CS���L�p��	������X��&� ���r��?Ҽ{�c�`D�]�q�>=�r`����>9�)$������!��*�1BH]1|Ȕi�t��E[�>�.�	"�����-R�9'�	�)���0�]>� uI�9E��՘G;�:��LsFO��2J��Z>\мs� 4��,#""&d�0x������7����@vR!��@�7� g�y��bͩ�Y`�&�yxmNYU\�x.ǩ�U�������~;��Vԭ��T����>;ł�\Cc�8�PF�u�x�M���*AW�9��B|S}���z�+Z���.���r�f�wu��]�~��f�)�b��T�b=��F^d���=�{���U�`ү���	A�1D|@�*p���E��S�{�ָ���o�5������'�^�5Q���n��wXf޹�xa����Ӝ(P㻒+��xp�d@#�V�x��{;�-'oȓ�O~�sY�тء=�s�ۻ����+X:�HqZ��e�:��}_���F��k�dB��8�B�����6�9�#�A���Et�8A��0r��ʨǦ�dOHe��l��� ~j���s��K4j��G=	�\���;����SmkϏ,������n��\v�,b�����I'��J�>;��>�����՝�D¬m��۝��#�ή����qq� ��3Oy�����v;][d͹�ڢ?����wü��r���' h�վ���88�q���H/�f{��z�Q�0��ލ�*g�����/�b	�����r�\���}��^�ԧ�Z�W����ϊ~ҥ?���v��q���誔��G�.KL�@�b��>��n�x����gHct��L��a��1q�kV��J�j��޾~Z���_&fx9� �X;�\7X��z�V{�����tGN�$hY�>Ց^�����(}x��cM��N���rn�ݬ�,��=/zV4 (�<y��?����k�e��b�[�k�3�c�AW){�<�dZ�z=�n^��9�ɺ�%��4oo�l������k����3
4������'��*�C��\�?Ӗ�j��r�_����zw��3;�Al��r�=<$-��Po1�ėӒ5�g�w�� e����:��E)��&���
H����u�D�#�`��W�U�НS9SK�k�����P�C!��"w2�ފK�Zv���R
��z��_fv̾F�o(#i���]�1��xh�m��`����A^18]��W��`ژk�{���7�4��(��t��̴{��璟������%��gUA�_E�����?��8/i�sP����~��!5�"�L>�������REZd"�&����PEin��ߤ|�0Wld �>Fɪ�:��p�U1�kͧ��<�潏P}���&��~�$qе�~�U�� ��/t�_����޳�#n��k�5�N����F�\��\�#l�l�_���F����(/s��$��>|��$n��ݝ6���+.�_[�L��&��`5>shT�
(T�}b�\>����q"[� ��2�_$!&ƈu��WS��H��_NF���/�+QmlC�]3��U��h���7�R��w��ws���
T�SW�tJ��!6���Z�9G����1&��r��ŋ�i$���+��3A���ެ;1���]�Cm�<�3*�(pX���b�yq^D�:/�����-U��l�Z����ej�Kc��n�|��F˧ȇ��ؓ�B_�lNk�3�Dūb��u����C�@�1W���;��o�3�Ѯ�4�V7"_SDY���!�J��Cm�����b������S�V�������q'��g�nU�I�2A�d _�a���뎽�.��M���%Q�g��p����?#&������¿�����]���X�^a����b'I�$'s'�oSP��(���B�"2��*:�|ݶ*Ǟw��ܼ�Y�3���Ԇ?�0ӌu���i�	)k�I�}r���z�h��Z�ZsZ��F�s�r_x���v�%���S����1w| w�޹>�Z�r��}� Co$�j6@��;h)�����r�`�Z��$$h: BسO�.�R��R�!(�=GK��Vq�'����q�\�b�꛼���7�T����_���V44z�Ѩ���V����(�{V�O�mcQ�LѶ����	]����~�'�8���_{>_��J[��6���Mjy���GGs��o�&+��?���-}I����;�
ʟaǰ9�ձ�����KT'�#�=d�ڏ�TD��ƤVx!�?���&��9Tu����;B��ɸA��䢟$^���O����dr���/P�q��UI�2Ϲڛ���h�%F�}4��MU�X"8b`v� >j����d����|�B����xM�2:��n�Ql �>eӎ|P4�����Ǧ�/wY_*g�c�]4)����؛w%Ը4@�߻�iߍ'P"	�o��R�/�2�Dc�r{_q�1^��g�M=�^+���P,{�ra�V���	g��b��`�C�K6NA�0P�nk���J�~�$���u_jL��o�Öp���zk�;N��}��.�e�������ܸ`hd@ؙ�üjs��ro|53����xGHl�0�*���5Q�<���+4���F������ep^��x4�ݽ�MM�Ɍ����+��p)���8��if��*d�[_Y�P\1��d��D=��$W�Z�[G���[�Ř���U
ͫW�j�V.����2���C2v{�z;6��s7�-&P2�贿xS6�TbV<oӲ8}5���&���Χ[&ϛ7K����,�y��J���o�R�z\_OF�����sbw�P)�ٔ��N������+�_��/w���5c����5�)�� ��F鞙�ʝ������2}lD��ÐS����P߷[��Äw�?d(~Ƹ��y~X���ce���PKi�`}��
E�>��"D���Q��.��n�)�2e�;�E���)Lj�����2�� �	)���q|�·�W}>�������y�'g,�[q2���v�@�n�`�!?���+ȎOU�w[�����U�#�vqyLP놓����8f�f+���I�ur��J ��5�`���
0&fb��r�`#wE{2�Cy���cń��?�j]HzN˭����������J�.���@��z�z���a���l �XQS	�y�25]o�l}��î�8�L�@����0�'��mT�g���(gv�o�!I�-7��b��CI|���\�s������h���{GOϑ��ǕIPߊ��4�'���8��d�l���:�X ��i׌ǋn��K��h�!��Ρ�r��'��r8��J)�#ȶ���(�6֤����s��Ub��nQ�������ޚ_Š��NJ���8H���/c�ХP�ye�[�Ӏ��J���}�Шֹ�;��˸ⅉǺZ���rOl��� E8IuY���e�zΏ�B���bi��[���y_��]u���}�{��m�=�d,��;�vz��C��o��;O*a*_����f��7��[vdؽ#k3�{�M�S�\:H�Fw�E2(��j�Q�B>��ɓr�^�?z�ܩ=&�]�Iٔ��~������5�r�Dh�F�zĪ�F2��{�!6��F�����	�^��_*��}k��9��Nu��T\O�prl؋�s��~�0������ُT�%��KorS�֜֠���
��D�ӬvUU챷�kC�I�A7��T����k	�,�$��@�4��Ж1=0�P^��3��@����e����(d����-f�śdd�w�Cb�����ߑ�K��v�O�I�I��c��Å<c�\�=�(0�'o��0�8�m>�)Rcv�����K\�������su
����n�@��!�::�f�IT��c�Q�g)K�z�xO��*"<��p�ݹޛ�����l���\�ZF_8�������T
L�[MR�ZJr��;����H�̦�e��"��a�݊�ؐ�!j�2��a/�_ ���K��N������'$�֚'�ڪ��IՕW���L5���/��v�sƁ��~�{T?��|Ϳ�X�Ʊ��#���s���;BמF�w�9V�D�U��N�̕���=�Ew+���B��˨ڥܤ�.��U�4�(4nkk�b�6�+���N��`V�
�$=Q��j�?�!�q3t��������&U W��y��.�+P)�/�F�ҋ����+>��X1�	/����jT�KF�	���#�{���ħ�z�������Wٓ�]�T�������oI~���ȥ2i\�h=�]���f��[�7Ͻ��{o���@�Z���u�m�[CC�=���f����`h�hϳY�Ց+P�+��?I����Ű2�h1pXT,+��Pl9�v�!�c�'���Pֈ��c��Q��מ�qw�S��aj�/ˡ�w��8Wm��<x$�������ÔI'�^�~�Ξ��יq���χ;�:��&��J�zo���|�(�O�V�~�}m�M�����ʅ+~D��L��;<�!�Gu��l�]f�z���z{�L�6�[��O��R�t!"YYY�K���>����h{D��"�R)�\^s7߹��u�9��m2h��M#Ѕm��;C���^�z�����*u����E��m���4��_l�i�8U�6ӵ�Uˉk������D[#$'��莛&�iL��`(��O�ew�n��W �^y�4�sUd�;�o�|z��ʽ�"J�Ƀ|��X8��W�;�5&iW�jkݭ�9����=�:�Bj�_q�����l��1�F�."�B�IMz�s_T�YЛTU�[oD^1����V��4���X&=�i.ϩp�������3��5���m)��ʮ�?�2xf��'� ��[C�R]����՞��"#Dn�=~M�ٞI2n�({-�ó3k?�,�W��a�AC�R:�\�nٸ�}�[D���2x��oEVښ ՝S���r%�< 6�LǾt �-��rM��-1YB����;E�|��;��&�w4դE�/��5�YD�}g��鵐��z&E�r�}���1����K��д}��#��}y/6�����F"lx��(���yMt��׃�[�9�fƦ6��L�t'�tO���J�6�T�� ���-�Z���pڟ�S�'/9��c���9R���0�:2�����w"����#��-[t%݈7��)dP��#�L�<�"}��W^�K��N����wīX0i~ۼ~� �mt ��jGu���Y7��%���f?Rq[]������i�q�=���=�ĹS��KV54br���,�-�W�?�L�Z�~Gw�\��F�����#�i �׭/#��1`���QK�z���4�^y-Kg��q�����3vz8�
7��D	 �|��/|[���g��L�^�cN�#׫���g^��/��V�%�Ⓝ�ά(݂�"�վ
��p
��L��!	*�ǃy2��	c���߾�x+����E�e��;Ť�sNqDȰ"ߔ���0�G�"u��t��k�ӎ�x�j�e�,��R�L�v�~�/�$w�������| �h����t/Tկ2s�F���5|g����g#@��*��p=N�?Gk~��*�Lo��i�����!:Î�x�tIf
v�W3;���G�҃�uݕp�q߲,;�3�����ޭ����()��5K��e����l0�t寛)%�}
��F�Nc�)-������>�<��u�<>������Zդ{Մ7�g&�;q�?�S|��A�r5�	�'[T�EA�/���<�exN��*3�kF>�SL�M5�٪����kye��ɏ�#9���u���߻U;o����?7�G6�v~:��ݰ�n���?Ќ�Wr7���V�C�Ta^
�A�t��Cp�̚��k������jQ��{�ԧ{ޒ�b��kt���Ov��Y�;�6v'�o��Z7Ґ����2���4�k��>���A��t�>!�li�"���"��y��C�\����~4ݑ[U=w�+k�K�7ՙI{��0�/uN1��ŽV�:��9���=���aj,Ӡ���	 �����؀;��{Ey�%�e�U��;	Ǽ=T{�g��ll�Y�ϐv�t�C.KܹЁٮS�Y��d��<r)𶀝� ��*BI����,l�(s4M��]�J��oLn�lG���� ��w�{�ڴ%��F^�]0��������J�~�C�o�fo���~v~�F�ч�z�f��z@`��:9������r�C�s����������t���.�����؅,�����S���̙�s�ԗv��p���.��M��U��o6J�ì�U˜���J3g��4�]���4�[���!�;���E�� *pq�11v�3�����ҥB�/֛��?sd�l�����e�x����6�L^q�$Ȇ���Q��V�ˢ�*Y�H��d (fH���92*}C�w.��W�*����g�X.6{�R3��Ȣb�=��P8C^����C�v�qL�ªh��R)69��U>B�o�����[j ��х~���@����wY��'������_k<�6,��s��V�=� q�"�8����rx����^��|Z�L�4�V^��g�D5���"�x
�0��gI�ρ�(��.����������v������v�?T��䰝yh;\�o+a��9�&Ө�mQ{�˫�OŖ�w^ϻ����2z��+
�=��=�nt5���|E�D�>_Ӳ�,�?�vz^\Kcu"��B=�ɞ�l�v.6�.;��m�H}ŝ�������k;e-���Hs������ő_/�>�%Q��9����R�L-j��*Yt	F�`0|]v�s����i
�eIy�+�[?��\󒞚V�Q�⻱'�)-�0H݊�8o1rn����P�j�v�x�ko�����U"�f;!?.�7��SO	����$ϙ�Q����`sR~'���x�q�/���#�x����ٲ��w����e��윜k�z�d����� G[�n�{�"�5ۙ��7���e��4kҨS~ݠ}�R���c�΋��*������8���?\2�׸���Ιcj�V듥%8���/A������e�af���:�v����o8���]0���[f��^jE�YTo��9��pc��ʾ���b�W32�*�`�6V��NúE��W�[�5�E��3��VB�Bj���F$�$G
�����Jww��KF�����ހ�P߿o<>���׽�u^���sϹ���{b�l`�@����؋��y����k��^f� n�W��-�=p�S5t� \����E���C1R��+�*x�kט�:�}�O ��|^Pz�ܬM�qu��(��;��.Ŭq9�%a��C�m[�;�[q�;����[������M����[���mY��2�<�4!�I̗�o�Ń��r���F�K��=�Lb`L��+�@����j�j�8�0��<�A:���+ڡJ��p|���9��lV����Q u?,���w�̏Ayzf2�����K�9F&T���M�'�wx��Io���G�6h��.	��X3Mz������?�Hñ�~Xc�$�B�m|W;��w�O��xP[^����zW$�9����$K�dX�{2'�s��8�|��>�84���L���Zr�țH�2:t~�ǻxxl2��+ZK^t��P���j�?j���gt��D>me����,SE6w�ЉA��,���uƕ~���X���}+�ߥ�9��o]��+��2+�l��1򶙀�z�O���age"I�"�f�� ?u��B#�G����XWY|p�����P��vH��_g�OFX2����MHS��3?
fȔja��fJƫ�Vm��8gN�4�~a�>����f�i f����KJl淾����?�0�(5��!5F#���']CޭSY��)���ӈb�f�¦̦1�!AQ6�7\�(�=�T�a@���9+	�u�uF�����܇lN4|ڥ���? l7��4YQ�2&8�x��"cQ�'y%<�}\^[Of�i)n�?[��Z�шC���� �R3�i��ڴ�ʏ������eN"P��_�R��R̞l[e��(�PZ1W'Gh��[+��-���s1K<���d��_���I���m<�H5�5T\1L�"�&)TzJ*]H
U�%:��CzM��P��|����z4FƆͨP�x�'���@Dd��JQ�&.�b�h�<��,=��`������T�vE����R-�V:r��ÊL2�_U)��:3�`��,�ZQ�O�~ՑZ����H���*���Bi'q7;1N:�YM�	-%����J���l7���{��X��֙D��Ż#UlA�Lu�F\^���a�UX��ū��5���-�q�9P�������kk��MBY*�3nh���P�ԃ��z�K�Q�FH��JJ/��h!�vn
����R�ψ?�P�p��Ti�M�G�or�_1��-�Ŷ���7����vz��hM+s�����B)k��J��c�q
l��;�f)��R�<n.�W����E���8�E˶�j�	��Iv��:gyPuZ]gMY�pL����,*F��+�A#����j��>fE+�t+0מPζb�~>"h�.cĩfV���|߼�xew0cx��ƪ��E�ז��;�����G=��`�(��^�y~7�{}}S�l.4×ҕ�]�q�����5�Dv���� Z�b?�mt8�T��b�X�����FXw^�.���T����NM*�f4���o�\e���n��(�(8Z��C�~��Tw�J����,|UJ�J��}��g��2�z	"	U���~�CPJ�=7�Íɖ��sC��=� U���\���"�u�Q��FOl���qy��~��Ƶp��{�HG�p��8b��0��Y�oԁ��_�p�&����X�aQc�Ƃ��ǏΧN��W�Z��ȯ���t���>WV>��X���Y��`Ŭ�*s��~އ|��q�8�3٥eTdӖNm�L)��'����m�NX�hr�]7I�����Y���C�}��H�E_���ވ���1�=E2E��	A�0���J��}�-�ePڑq���'�����CM��O���?��&E�LoiD��6a>9[Jw���q�a'�3��.c�y<�<	�����Θ�wa9�����~��yχ��4�藡��g��p٨Q��,LH���*�2FՑ4��]�����5V�l\5�Ͼ
�
�p���	�h=���[c�.J-�����N�|c���x�!�n,�O"o�Ifl�Tm�-�� ^�&!kD�������x�Ȟ{�m}�<�`�5��#G"����b�|ԏ1gW?�$�(������4������&��YHx�S�<<
���Atÿ�2�}��Ⱦ,�S&A�5U������T��-y��ڊq��*��>�> ���!��RϤ�,ݙ�~���N�u,��sD�gt�[|D�۲{�}9�Iu����jֻ�nwµ�BpF"�F��	!YJz��k_��^~ ��6m��Nhr9R�^y�:Oc��b�<�Ps�Bx-<Ur'T���B))B5�V��q�S2���+5�m��-t��C�����ςxn�ܽ�5�b|��Eځ�;)�OB��'� ֊�S��ܸ��I�U<�F@���g�'[[/7Q�Q�3_��w�v"�q�^QЕ�0�'��{^*�T�����c)fV?��*�U���[K��P��띮����;=���^]�7F��� 7�x86hۇ�ǎ�^"�*J���?�F���?�\�eՙ2<[~��x������Ò����� �a �$��2)�0l��E(�/��P���Yfjţ��i ����̻BU�]{�hQ�K�� ��γu��}Ղ�����uƑ�m>y{��ڂ�=iid�v�+ʿ�k�`��Q�j�̚^AQk�N��2m�횕� 1�tQ'~&�U�
j��� ���u|���%V1�$q>5�Z����<N�q۟xZ@B;I��	�
�$���ٜ^}=��5�*Y��@�=Ƕ^`��d�l���C>�-�m��7y	�nR��t=|=�v���۔�7��Ѷ�mL�ɭ��z;�]��N�½����T/7�((4$=��ۭ����d2(O\Hҿ2Ȳ,���=��M�q$+`�/p'�DWk8�D�Y��q�eyU*a���Sp[[[����N�?;o��i*��w��[v����98���v�i��#ބ��}aߒ�7����'ͷ�׸C�^�R�9r�Ql�'�C�zR}�Γ>z�4wm� )b�#�#���RP� ��CwF<͡�Y�W$r�V}R]�T�D���_�b|PH��)h��_�9@0A���ϼ(y�_�,ភ,Y0���{܎9㗝�J(_/�)������x$�7m�z&8�|�� �|/}�酻K��;ٞ���Ӓx�0��u[�5���%�β"���DOx���b��9�H�\�сî�ae�3��3���l���ʔH\B�����}׃r��NsJ��j���O>'$��7�z�G��p璮���nk��/̗��~J�]*���+6���K�B'A�fR��$���������'�8��
��p�<*��S�S�������w��d @xeQP��/���j�M�s�W"�v.���[k�Fμ�R�4h�[�����%`/�pb��b���$0/����(���3c{H0�G/&Y�c����7k���fl{�)��z�vz�1�8��~��<�-��itFKzaj�M���V��hf�A�s���A��\4>�x�|J:qV�
��S��G�$Q�ް�6������s������}>��1�Z���׹�ş!M�������O�k�n��Q0g�*@N��m��y��-}�-�!�vƆz�w�w��&s��ʘ��=�|�+��i�`-��������My��KE� ���$� d�����C�+�ז�Ӎ-�|�l��(��W��:��d]owI.YC��94�D�+OX^kɞy(�S�!�ͷ��G��������U67���Ư:��kխ/ ����Z�T�uG�ۍ�ӫ� r>|h�����P��V>a��+d�+�ҋ�6�fƨ�������v?d��s\��y{_}�E�](�()��4��)����������4������i�ɞ1��n��~*+
�N#义�@T��D"vΊ��@�Y�.�y$����Y�S�����(�Q���*R@�^%�r��s�H^��wb0�"�'����~f#��;k��c�8�,#�]�>���n��E��$7�N�K{��ΐ��r�����˶e�6P�D�Ojon���~x�����?D#�9��[�H:^�`O���%��^K�	npſl�%�0�Gi����&[��`.7�y8��if̙�������>BS�%.7i�gFW-��G�.����-+3�Q�[����@4t�x����o�����Ic��Y5I&o����"vǆ���糿�ܻ�v�6�m������?����v{|��eW�` ����FȬM��g�2�oc:8|\Vy���X��H�T�_L�5�"11l�"���ة��X��t����Qӟ�@��#�ѪbLi�i�g���&.�y�U$�w�:��eP���L�+dј5m�Q�~N���3����2S�O�͏/�M�B��]$GK�.M,g+���m�f��M*�Sb�7+�-wqi�4�U�o�{�G��n��������P���i��h��I��ǎHIheK�.14Q���}>�;_w�2�[�̟�5;c�;�S����m�w`/�'6�:�9H��5sb"�ؓUO%}My�l���35�X�O���i���豈3z�䀅0ywku,j�U��#����ʎ\��懮���7[�^�����������x�/Ǌ�m�B�u��f�Ƅ;���kƱh|�X��]�Z9��+kZ���6��{P��/r)W_אB�3�M]Z!���G�f��� ڒ��h��I�v���"=��NYx|���\i#b*�h��'��2 �n�O[����?5*��֖��*���Z�*��>�^AAӃx���WT.�C���6��2<��m�,4bZ;b���7șϵ\�m-��4Ɋ�ۋ��(�ppY'Jf�ݮm$ߊ�tT����Ѻ'p�1�4�bPa�4��9gK���M�������Ⳕ{ĕZW�J�W�k�"���w���J+c�W������<�"�a�M7�I6TN��z��)~"�����7��X�(&.w'	����"�~j��a��?F��n0�t�|_m��'�23;ݦ*A�~ـ����U�|��Ҋ���+��~)
e���Ee��M~BM��z���5/w���?ol��e�`C���\��6��N_^]��H�:H�;�U�@F��;��%e�=����+Pj��]�D�0��0<�}����d�j*ǅ�^����N�!�F�1�����1��u��A�Ȳ�:�K U��HX\F���5�6�@e�8��4jw��#|�c��d���N���-Tf�,�*�uBT�f���x�\�;[��!�)M�{*|v��j\�:�Km5�ba�jӟ�=}d���;��?|k�O
��I���eY��2i:ZqI��GFF���J���~�ܑKF���9�=���K9�Ǻ_#�os1?�J�x|&j�*���~|�|;��)�H�����V��-	��쪵ǉ.�/�I_"8Dqܿ�0��&ʦC�|;�M�fK�z/�IH4��o�ۓ�?6r&q�^�=ư�������
ֆ��ğ�����9���=hB�H���,��O�����=Ӿ������R��x�cV�����Z��HR�Hy�/�ޑ��+(ڢ�
:�&n���~�oQ�i~�o��j�@O�������n�h�KOu��㕺{d���#�m}��q�Vo9��^��lY�и��{[բ�����K]�#�������������l�+}�t/O<���( ��K_p�o�[��f��)2L4(%BX������8j��S[�a�|/3�Θ42tugm+�߇� N��� �5�=�8�5S�4>±�^�|."�*��=ŞR�2+�[��3�i���A��7�$sK]����N�?�5�n�xc|u��q�g^闕LM����s[��t���s3�W��*�e�wJ)��ha��ʘ������r��S����H�#������z�#<�koI�\�P���h�e���9��L UmS��Yl-~���&�ilq�Б��~}�a"ՙ���� �Ξmi���WǵO՗��Oc�9�q���E��5��*��[R�� ����?����O�#���(�����Y���r�[�%]��r��'��"m��t�ʖ�|�q7��l��u�%�$D^�㛏RTB���$������f��g����tPW����	��yB&æ# �*�L����?S�?������Rl�R��%J���K�}w:&Vm�����<��N����8ߨ�JW���pg�����4S,U�Wn��:�}�����u,��gXWCH�~m<��'�ʹ�Й���Ɣȶް���6Qv7#��i�ǜ^��j5R��`D�^@�5p����2�3m0̈�Y��%�X%�t?�%f��if���1����l��O�ҝ��M1f��=J�S��{�6�n�2
���>�x���7a��ڃC��'�ؗ	�s4�'����,w��f�%�2|�(sT�#7�=+-��E�/&��/*�\��n0i>�%Y�n4֪��]L}��r�\��s�}O{").$�Oڧ��eU}�mʮ6�O�Nߎ$,>(�Cr�6M����[��7	a�ת���\�����25G�Gz��0�>����۱񢺤bL���ӗ��'��^ZW8���:+ZN����lm����	�5R�cɲ�u:Z�~c�w����gZ䰱��cj���:���pҭ�B�_���밓;���Xs܏F#xj�/%q�UZdBǟ�@�J� ��c�@��sV/��'��"��W�Pd����j�n��He�4U���Sꢜ���w�uv��W:kN��>���R�<a�1�nx���#$$�W����S~�zԫ1E�����	*�E��(��v.�#�;Ub�|f�:CZ�y8��i]L���y\eHv(���=�9�x��u�-�B��*:�j(6Dq���̴ۼd�I���,���9�& �)�E�~�0]djj�;RMx1��D��e�'l�Е��;�xF�w��ޣ��m��ڊN��^.�`�ck���#��̻+�Z5��x�l�o<�o-�]Yc3�l��k�m+�p^F��"�T��ɯ��Q:�D�5�^>�M<��M��xn�f�9c���(꧓D�C�V���A�	�5��g5\�/�tb�Ni$���z5gU�~�ܐ��e�m����t�&��y�w(���}n��[d"��}�FH������(����9�mka�ʏ#=�UsPg#xd�R3�ˊk<(���jp��a�<��Ύ%?o&��~D֒�R�ȇ��^���)���>�Y�o�L-�o�{��$���NTf͛v^�Z%Ia��M�ly0+��Ix2A��J�T����i��q-���Q�Ɓ��[O�Ù�`�Y�X��w�f���%՚F���ᡡ� c�Ӥ�:V�￼��X䔎�h�����N5��,�`9AQ<jH�d�>ƛ���5�{�J�R~��.R���S&E�Z%bV�\3�� kW߻s��D͏/�^�}���;u�yd�x����bo2ݠ���V�W���t�/$������5�/{bڝ�Q	̰�O=�c��Yl7�$aV�`P��h;���7f|)�\�y�ta��"�<��P�!�Ea#X]'l*6�2� 7e��b��4��^���Б��b���T�x��CdC�F���%Rvc7I^��k4�I�Hc��L��r*8�=IaѬJt(�<A��&Gl�!ˀ�#]�ᱪiVKGQ.w��F��j	k��}�|Dݣ�r�ݓ���l��~���L�~Y������2eqG��䱿���[�~z��j��j����X�)?r��5�I��\~��1A%�öQ�x쳨����h~Br�Uf�ؼUz��$�i��i0��Ǌ�D� �;7h��i�{��`j��Ng���V_�I~c�RC��/��s%�Y�Şf.������T��=�n�׷��x%��M	Ij=G��3Hb��Z��?��8��=U�
üx����Ӹ���̿�
}�|8��56AY
��K�<�/��V��]l�c(ސ��x������N�^"���.wo-���K��U'%�3���N5������=2�x�\��v�@�a�wT��t��-��`����+W:|���&=������iydy[M�#N��Z+l���%3kVm��? s�E��5�]�[8��p�a$��l�[�7���w��P���.�:�ĵ�"M�Ү#Br_����w�:|��No�"�� )-���U(�/%ѝ�8>M?�vC�>��@���_�Q�t����[��n�㟓�X�m�r*!�ʶ0B��[��H>�y�uvޭX!��!��� S��6ש����B���
�c^�P�Xp��R�}K��w���JW  U�����Gw�P��qg~�q�H�Ȋ�&=���ڝ����nJ���ė��P�����a�4�準��=QUc��T+:�.�3{���d$`3�RX8ۋ�	=�&l��fH��TȢ��y��O��� ���Q`��N��S�Q����i�^�5�w�/�~/7��N`L`Qk���T�����)�����& �ɤ�8�!��Q$a?��R��.��%�g�k}�������V��C�ɭ� ���]�Gf�tb�$`�]~P����]�b��=D���OIK�:�"lش�'K\8�ھ���LѢ�ݎ�g5��Z���`��g
�<�G�bU>�nL��l�fP�ƹ��R�́� ��/�����e��[kw����<�򍫠%��=7ĝ�l���H�b'��[��uڂ@b���7Z��t`Գ+�<K����n�(��Y��k���Ѻa�S�D�v�^���n����Ƣ�H���[49�U�ϊ��L�b�ê2_� +���
�+:��b���uuhKq���rk#h���M)�2$q[�]b�=���徜���4rh�&|a��{lh�]�6"e��M���+3m䅎O:�v��ߧ,��O�e��ȸw5=-�Z���5�u	�d�,�����bO��>2H:B{�&׽���h�xQg���$�~�:��葮���d�����9u��#��dSzŇ�	�-�8>�fe�Mt;�5jJ:�����#�u���Z�R�㧩� �� �f�^A�G�� )Py����4�����x��GH�U@ͭu��;�D�%T�-'�:
%�W�T�<�_��_�hD��;��,���@����Y]��_XN�"�����cf��^O<���&�D�m����ID�V����S�쬐g�P�Ő;RQ�u��5�'�Vb"�S��U�����b�����(O��C�e��<]�|�����.ɼ�V��ռ�F(>�#��X`*ꮱ�	��0���>Mi�g��2�s�(grN(���1��?�"��[��oށ�e^�g`sI�aV�b[)2�zΎm	π5oE����y�w̪�����OU�u N���S1���%�a�뿾.�dM�{֔pel���j�	'h��pN����ޢ��|oYݗw�&.E�Z8I�)į��������[��5{u��,�FR����<�(��H����8e��OT��������d�x�m�{P-Oǈ7�K^���BC���ł�9���)���:d�R9u�ǔ�C���5xIn� h�mD��;r��l�����=�w�ȷP��X&�/����դMx^���T�\��i�E���p.��Ju۫2v	,�ȉnE�mѴ�j�h�[K�g�������[��k������:����K��U�#�w)�c&z��Ǫ$�I���\�Օ*�o��n�ص�(q�"@bͽ�w����_�	���骤M>���ګ�ԟO����:94���Tz��K�>�c���@�P��XCq��h��}Z�=UK�G��S;�,y�3͍&������6;,���}��"����j*|�/�X��Pb�o���\�5Xx�aDc~���X�X�X/���;Z;��.���B���m�;Q�8�\�Ep�����UT�meo4��˫�Oq���A�"�{�~:����k��C�pW��YXq�[�eo0u��.;8ܯ��ϡ[�n��G8�L�e�)��֚?�naee���zK����ȓ�O'm��<�Jg�I{�Z]���{ځ<�u0�G�"M�/�V�Ty���
�ք���9��Sz�R�e�,�-�y�E��r������We~��\�Z�YG��r�D �!�}R��c�s��C�d�rV���Q��:��'E�x�W��!�Ԙ��k�M�'B1G�&>3k�2�#4F��i��=��¥,�aX��������O88�����H�ɐ:E�������N��S�D|g>���+��rیݙ�b�HL#�����:��E��L�/�&�R��>ʼ��M8��2�j�^[�yqF�$�r����#M*��wcL�M?��</RM�@�/c,6snډ�d���x/X��yd�af����S���+:H�(5������ŞR�1��!�u�(�j/yg�����C� ����p�բ�\�.5������(ђI�[�ފ��r��!Y��1�醗l�ɏl���]j~�A����J,�{�W�J�zh��&am�X��ݙ���o���2s)��+4��97Rݧ��9�.�Η��ܢq�ɵ��<��d������TX�I�D��˷��>�D�R�����b��ˍQH���ƩY	r����,0&v�\�
KNH_T��T�2&g�:rj�;��d�G!*s^�uа=�4�2�%��O�g2߰���T�j��q��Frf�CU���D�G�pzS���׻���""��[��,�J��蟅�Ћ}X�z�H�`�(�j�hy��R�<��KIۓ��&�7���ٕ�3r�]��n=F����H�YW
A&$�B��5C�����b]6�����=#��߼���ﲳ��Fk(���:=�L^��x&u��A)�z�hT�J�#�XE�����`?���z������rr�cz��͘���7Ό��y?��u��P��c�Zſ�%/�zg�D�3��.+��0b:�<�������D&P���tZI6�����]p��$?>^H-c�l�[S�M$�`j2��j���%A�4Ӂ��7�})�۪��ϟ_���[�����<���,,�B*��`w*%J�Dx�6V]�I'�X!}�F��9�`�4�H:W�W�I)�'��f���LA�As��I��溻�/�y�?������Xn�N����3������P��/�-u�(�{t��{Պ�C9{
L�.��-X)j���')�� �x ��C�,G7�5��� X��ؒ����!W"W<��P ��r6M�/�ëټ7��h�Q���}�μ�wFᝬ�vt��0�� i��a}�|BM7��O��O�ioo4d���I����WW�	^+��Dk0%����hWp����g���r��Yw�gKo����G5�/�t�~$s/�����<|3�1���0�D K6�����Z����-�R����x`{�:��	CUC-��',�N;9Q�mEq�]�R��[��m(���2���M�\<�&���q��Y����fj{q_�h��{i8�f� p}��[�n>o��o� h>��&?�������O[�+gq�������)�T�����+h��⡿�ͬ��(�uk9��������,|Y��(�h�	�����9�>
������C-t�MЬm*��]1-�%���f;==��p�%f{c������)j���c)��Ei�w6��滔!�d3%R�l7�Ή�-0��v�_�����;w�z�����8kz�Ii^VY �b��G�Ũq�N�d��#O+}���[��n!btܗI��
�&h���4�\�4�Sn��I�1{�VL}#{<��i���䣶{\���
��Q��n��ߚ�:����"b�;E}�	5!}�K|W�Yg3W�Km�I����͐G/�W�d��WE
�O6��&$���V|- ��X�����O����j����;M~4������qHC�o���7����
K_�~�O�X����#��y����N��ȹ�B���O�8�3r���o}	s��N��%��YҼM�72�Լ�'��w0�U�'&���=����?�9"��Hk[�@f��|�_C�T%�÷ǟ��e�Y���
U~�\0B�]�m�����mNL��������38�~���vr��c1��ƃA�ԝ��/�oI�ѐ7�8<*��\#�{of�L$�=���������:���׆����Ί��*H(�#ض��m�!�\a����9J���5
�����Im�DJ�/lQ ��U�R˜��<������	(; �6�t�q.�9�
CZ?8�=tp��+��_�&)������0/��?�4��x��&g.�FY�׶7>O6�U�߼�I���X�������1��_�]�r\ƾ�^��'�\�q9^W�?���7�QI��u�{O�Kw�di���|�S�s���g�o9 M������=���� )��-Q�v齠|������=#
�op���-��F'Չ4��)�r��w��*HS�L����PK   t~�X����H   C   /   images/8e6e9996-4250-48fd-a42c-980e5b13088a.pngC �߉PNG

   IHDR   d   4   |l��   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��|yx����=[2�=dOHB6H���Ȧ�
����R��jk{�t���zi۷������R�*b�V@TY!@����=��d��=�L&$di����I~�[���g��9Ϡ�Y�����b�x�Ǉ���'NwC�R�j.�s��u�B��Z�?q�'-jJj��c��c¡�v9�v�w,��G�O{5:L�	}xߋ�mgI34�o��RB��h-��%C����v��:as�q5��Q89O�2{{Z|؟����,{r��
�:6B�U������B̞1}�������N���*�Z��Mya�������\.}2��Á��V��P+ZL�o5M`�����3�)++3(o۾� ={�ɖ�j,tOrL�_�:��E�]�����������S�qy��Mʰ:7�-Σ	��my.�cA�	Ĭ��Q�Oar�e^�3<C��Y�e��w���k�5|���Pw-��X�'V翐�����mGOgZ�.��e����@�� B�@t�Q�֪eR6��f�賸au)}~\���e��^\���RM�����FNz2�:��i'���G���E+�AH �F�9D��59�X��5;e��DJ�V*����8~z�ɷ&'�{%8P�����V6w@�V*���j4t<5!6�ʖ^�4t�	Wx\HU� c�MN����H��BhH04�h��h�Z��׏��v�jơ�N�t�`�0|=0,�H�����c0(*�I�t@���p{!���1==�s�0-k<�b���@Q@���fC���ӭ�8^݂/��Q�a�٥5�"96�/k���7O�}s[��*��,�AV豿��������7�"�X[�������i!��T�wAI㓑7m*V,�A�ށ�GK�i%���p��Ac������D�.h�k�W�I����~�(��f�c�iț<������zss�`�utuu�HI����k���U���� �m���Q�D������*�
n��Wb�j�3�
��	hii��`�
!�������T���a���������CxsW��c��'�e�A�ų"`�*Fŧ�jZpOON�����W"V>/y�%!xx��#8�h)���D{{;��܌��^!:�����0aRRRI�187%%a��|��{��8��.�O��9��zΚ��-�I6���+������������ݻ�u�V�<yR�Ɏ�d�J�PZHFF�.]�U�V!++	I����k�?�8�����e�U�5Rg�w7Y�ƣ��	�"'#���?�>���
M&�yY�F�҅�����~I��r~pЌ#G�࣏>�W_}%��K��S	�������E��zsss1.:wݴy�����wa{�����I�ya0R¼x��B,_�� X�"�oߎW_}� 5�e��F=:G��Y,�8q���X�~=��<��Cb=�����"�����r�Pغ�f^��һ1))ڀK�C����}&|Yg@u�Opc#X��S7��{�,CHX�X;�?�	��n���3�*��+��y}�x���
Q�w�yG@�я~���Lg*��X$��ފGڅ���9���T<YƳ�Q��Y"q�������q�F�8�d�PrK� MVE���dF?i�iP����_��_�w���ϟ�I�&�?P��ڇ�]k�83g-2���Rf���$���g)�C.L�g�ñ�%y�B4�9ߣvS�䖟X���X)q�l6�7���/��Ʉ Zg�&�ؙ��
^/���t�J�`��[��o�>��7��ʕ+����_~�k�-��q6&�&�f���ibFSS~������iub��� L�LG�����F&Ǉ�h���@{[�O���|�V�Eyy9x����X�b2H{��ף�孨��H�c0��`4ۄy�"#)
��:8u�A+ٍ͋9�0c�x�t�CK|>6"�m��n��¼t4wP\݊�-2�G�����߂x�n�Y8��r��100�g�y���D��`�൦f�#�,��(��C`��Bz��q���vY�^�Ǐ�cqs=� b���Խˡ7��%6ӛ
�(f\+��������i30uz��G1�?%��9-@�]\,�f��T)�ع��� �F#�q����Ǵi����v<��ð�Ւf���z�"��ff�AO���!� ���us�VbޔT��eAv2��}�
'cJZJj�x`�l�,vܺx�\s��E��?�Q���o]���q��>��h7��C��&�!o�L�Q�~v��1�x ���D\�R���܂S�J`"p���{N�����GJ�<~�BԾ����HLF��G*��U� <"2;v/~0xL��M$���?�ȄU�O9����Y�/Qdm�������(!�_�BX���������n�K�Y�y�t2o/lD���l�l[��SR����퇫�EI
rRĪq�dQZa0�SSq����Z�;<XK�ha�9d^��5��ƙ4�	���� Afdgaz�,YӅT�����dM�QQ(:p]�bM,K&9�/F��<ܽ��o�aG|�y�z�Ǎ��fbJN���mۆM�6[��=u
M�-�����u ��i���iBPp%N��I#<����7^}�>�P��^HB(������=�P0W�jw���G���0g��N
�UL{�	�����ാs&���6��d塺@Y���:|t����Š�!�E����)QX4o�ģS�Nᥗ^b�H����s|5�`��
�u�'H�3���%2��x!����=��)S� �<����`��F�u��s�a@8�'�����>�'6,(�C�I���IS'K��+X�J�H۬V�\32�
$���<AC~ۋd���q;�|��K��c�	|7�p�fcav�QL�B};�,Y�6�-���pk5h�6�bs�����(�m��RJ�0�,�&�<��M[(����u�`�,C���f�x1��^{}}}$�-��ř��ȝn�:���!�ޡШ��{Y�V���B��OwJLe��Ĉ�����3SQ�I�0À���ɈFf��{׮]�Y[8�O�1]bSvO+�&8�%��vv��7�L>�4-��$��T,�����g���Ѽ6��P޲���֓� ���LEc��fsbDPf+9R�$����Ҙ���51|o߀e�^!I:̜�-��4~�Ν�r)S��|!*~ː�@8]kHl!�TС$r��x�?b\$&Q��x�����vYI�����{��c�Q}���B�<2����l��ux|�NԖՊ���\��`�X�� �W�J@#Ka��Қ3o.N/����~]]�$Ry�iH
/BC����$^�)J���tW94'���G�+Z׬�����?���az�������n��p�.X��;�e����jQ���Z	�LKANB�֛I�J l�Q:%rғ��B�؟2�<A~�
[�m�B�g���_�j����3y���db$��u��=zT ���AV\��p�5��C�ʃ܌DZ_ �/��R\1��#צ䎥�u1��3� �:>�aוH�My�S�$�˗/��w���}>�bB4�����\��:O��:�؂�'Iʔ��-�27���ޞ^�EF�ű��H21���Zy?+ ��MYc�WjpHP"5!F��K�O�<)w`e.���\�^��5)\^���K�Gme����Sl���'FQ���k��R�@}ȣ��U\	�I����Sc�p�e�����5(�
����v��V�K<A.Nr�NK~;n\���Tx�еJD���ߜk��b�j��Q��� W
�m���?}����}��a �{�A�/TK=����%�`���ݗ��QA���6��5�`.E(����X	t�@J��[׉����!-�r�w�}�af5�!����u��Ā��:8V���rrhw�`YBۆ�����-�@��O�Juق��:���pY��D����|_�0z� p9}�Kz��{����0 V
B,,h�����5ea-%��;i�<h|��XK�W�9�:����؛�{����8씧8�\���������/!��'��i�)��}���X9q1��N�P_�jw�)��Ff�qXOLL���o0צ���M�R��C��;)	�Sk~'�D�tW��p|%��D����c6L}�UV�v��a�U�*�4�r��^�N�db�M.ޚ-�=Oo�	z>��D��ϻMNt�(�NEzz:"�]q,��%ם8��=�)����b�F��Q¦PKi�=�շ����p�qM�,\��O6�=h�����ڒ(q�0V�F~���+>�
	̸��� ��2q����;?��w�."8��}p�)��B��Yݨi�cf�4����P6�EEF���q��#�&�G�'�����)��mX`���K��]�b���={�\�Mϭ�0�J��݃�is)P~�+Ic�����L���66 ��U��O%�����
�`W�J����A��FC*�{x����%��l�����cٲeؿ��.q.\ ~����,#-3�Cp�|��٘��.�x�:�a�:�;l�-s� ;;��@Em#�\���"�c�� &6Nji����F�]u8y	�q|��[Ɍ�uaP���rD��$���5��g���Ȁ�hjmC��$uAëf����Pd�p����E*��z=v~�V�^��d)D�R3ӥc&�+Ŷ��S���N>��gS���r
g����K��j1c��Z��\Y<�&V�6���:,��EAA�Ν+JȊT^r
�/
���J�Z��ű�<W9X�آ��J��bs��Sb�L�V�^����1v��
mnz�Y�E��6�����Id��3�>� ~��_I�ݻ{�⑛7��Cu����}Z#�`4�IBg�Х�D����<!+e��Ipsб`��N���{�;G5�.u\l�$nڦ�����;3O�G��?���Ue����c�C�x).(�P�������ix,�_�B+[���>�2��6l/��-QC���C��6��wO#3+w�y����U�-��$�͞�#����W��9Fh�>6�4�Y��Ox���C�슷�<���B���Al�u�F�9E�1�s=�� V�E�z��'۱�D��?Gv��{��K�PY�I!.ܐ��s"t.~��G^/ˢ��hnh����~&ۣ�7>���hTg��(��M��N6l;���(�췿���5������o���� �����~�Q�P=�'�A���ȧ)~�q�z֬Y"ރG����U4g��gh���k��i�F������T7wK�W��C���h7+�����JCTL,�|�I���ٳG@9q�X����dS��!~|p:QT���&���>�(n��f�7����]�{U���O� ��=Ԅ�̃X{�R��*6皚i��۵ՕU�6#_�V���=C�Tu�:�(^�46����@��׿���.�����K���::v�ă�CT��6�GZ�	Q����'���'�s��[��C� k�	ύ[�g��rf|�?�{�R���?����,�RGk�loGVN��Wt�[T@�(���O���N6=�e0�������\<����l�C��<��[������,B\T8
��A^^�~�mq/���İ�(���>��01��p�0P�����8@ԸG,�����yO[�ڵk��v=^ܰ���"�Q�F��I��w
{,r���zS'QgàPU7�E�E�D�t��}=s/2T�%��9<\�4�����<��|V��ؽX�l)�������f�͛7����?�*O�b%u�Q�E����k��$����o�y��`��!�¥eЄ�l܁��]R�:{��e�u��y����4�ysfc�ĉX�n� ��[o�����4�Y1BQFm��I�֬Y�'�xBr�yԞ_�16��WFvC\�	"vc���[G��99�������ơ��$J %%�|�ь� -��c��/�)��{_ɽ7^����b)LO�Cp��˙<����ԐG�[��pn�.�c�op��u?�+;��R��A�%��_�T�O��9�6�K
%���?�Nז-[�^__/%��2È�[/��-K���1�PQQ����������B�������;��/��~�_����za�!.2f��p�NO�����X	yK��y�K���ݶ�Z��p�s�=���k����QUU%���lο^�e����[n�E�8qŃ�b�{}�gX��	6������l�A�����QZ���+"%5E��2[`Z����R<�dq��� צ�<����38�I�~v(�+[�q���ۊ:ƻ���Ĩ0vj�x^;opX<=Av��� ��w�fwbRJ�����A��]a,���a��M�J�U�g6�@9=��51ib��0�w�}����K����if%c�c�p	�����j���'��������_���a@������_5�l��48�x���+����9�v�t$%&H �5�_$���|�� ��t�xi%���>/�ɥ�(z[�ԉ)�@	[��9��e��_Cy��ٽ���k �}/r)��˚?Nb̠��[�җ������݂�da�5��?$#<<LX!���-eT]�<��4�ʚz|��m�~з�y�9��^8�zd�λ��b�hQ!8�a��`��|/=�X�D�{%��]�ES1wj2SE����el#�V}'J���T3�6a�+d��X��c�E�/˛�*\�m%Ƽ�dG��J�|qEjE�r�d���dF�]�p��ε���PX9�����wV���X89��i������Hى��N�fqb�lFGW�j�e7塚��<�Ϯ<��c�u�J�@g���>���|7?����#!2hgC����R<�X]�(Px��0<���r���F\�I�:y8o�d����g���`���@�����[�NKV#9�E��`�-=�PJ��`j��A%v�:�r<�	� .�W<�8�M\���fŹ1>�Lא�����o�i��&��A��V��e��w�8�#tDE��0�[o���n�[j��x��Mf�iSR���-�NLJ���k��yǩ�>:� uTh �Z4���`Ɗ���<K�y��w�ԩ��D����~��a㲒��v��>3M|P�r�eu e�
�����H*q��Eh������]]������J5���Պ�+gG��Iy#=6 �fD�q?]�U	8F�ێ���]|%YV*&�����h����[���/?����K�&N�uw,�ؿ|IMs�|�����������j��AZM�[[v{fg���{7��o �H�_��,�T(��v����C�!\��\�s�s,a0�w��3x�3�Yj�(R~�C��/������"|H;[��7����gz�� 3;X�_��܇c#?i��~�����m�o����H+I�3�B�:m"�v����T+�7�"W��T�Y�(��}��A2��6#5bQ���+�g�صٝ�-mM��]��ܜ�����`���5��&���ge��>����-eM=A��4{�+�D���9{&��Ӷ�4J��:<^���N;~��YAnS�pzݬ��%>�ʀ�NE�t���*��m�C�V���xlN�W��f����֣�)�u=1##�a
A[�N�?q�&�+f�5��A�/��z=Qĸ�o~c���m�OuSN��F�w˺"˟c�U����������[�m�[�Z��
u��m}�0�@�b�k_Y��)5d8y�Փ�w�=/�s��~l�R��dl$��q7�G�����M��/�&D�vI�T���Q��؊�E��	
E��A�۫�X���w2�f��3m����h$P��� H�4��e�+K�.yF�sq�6�i���kv��q5���qa�e�;m�>zW����/3tJ����UM�Uc��s����+�A�fqZ ���tKcZ� 5 |���MF���P���__�%��q��ߎK�r��o��Ʒ�\e�[@�����lS��?�    IEND�B`�PK   ���X�O����  � /   images/90427f57-b7b1-4ef6-8fbd-3930b2051391.jpg��TSA�/z Qz�
�J�.5 �EzWPZ��D�E@@iAzG�Ћ҂�� t�$/~�{�����{�����={���̐����jj ���H3�{����ߟ�.��ԗ��/\��BCs��::�+��W�ݸ~��5Z����n2211�ѳ�23��`db��"��@}���2�Uګ�����p���6���������A� ��I�K���]��t�
�u������տْkB�u���E�/��IsǃQ�m��K<�+3=�����|������.���$$���Ȫ<QUS��i`hdlbjfn�굽���������@��""?~�JH������[jvNn^~AaQ�ϪjDMm]}C[{Gg��O�������ߩ�e���z}cspx�=>���Q T�=���a �Cy����PP���d�@}[��e}��7���8�{���<����l=��0�J,���c�?��c(��G�����i��� / ϲ!�s����~�g)�?1��_׳����^�"lt���I%^�{T�����F�y�;t�/��qsI�p5���)���ַ~�P��f�lBC�w�&T�0䃗������V\�D��� qC���9D���[�u����=�z�5�\�ۏ$F�����Պ�z��$ ����wP��U�c����DB�۹��a����w��͙u��M<��S�&�A��뒀�q�
	Pц�l��Q�o}Sz�~?����Lͩ�v��ad7n����D	�V���i��TEޘ���.���R@�:���ϴ��x'�E����l�����K�u�7���6(��O.���ڮ2��EZ$���T�̥����	\H���oku��zq� uE��V ԜL���g���D� ×���Fl{ې��KV}���&�Z�Р(u��p!�L���[#��J
�޲m ���N(0[�����(x%-:�׺��`��w�����=íC�ї��H9B��e7���7G�v��7��C-761�P���t���K�у�gHuB��_�,���Ƚ�F�Ý.����G��k�BL�����	p;�%5�'S�9��<]��G4�8���~���ٺb�����Z@ں?ӊ�N��J�b��YS�X����Q��/x,��=��ϳ��QRK�[���̧�d����V��ݜ�˭��6̺!4*o��V-�7CV$`� �_{�E��zw��^ z����C5��M����W2
Z��A7��+�z]�qQ5)���W//zu�>�*M��)�ǩ�画sYI���v�R;B�)y�A(�?[�tbס�*�
[�-X�"kb�	�]�'����P
�Z��>�l�W��ߎ�{�@/6��F�������䕽�X�,���������8N��2~����'ne����w�|K���q� w�<�B��ыwm:���hC�EfQ����N8�?6|��w�q��7�ek&�>�C��\�}��pUz�$�B��c���5��-�铛�H �u�d����iS�d����;JP zt����;�BgI�o3o�C$	�$U|l���,�g��[a�Os�(���R���'��34���A(N̬>YGM��0�Rj6��F��ٌ��aC�iD�p�:d�/��l���(^|��l /��FS���9
�%�*�Ob�j�3fr��B~�In�pl y�h�~Ï$���%ۇ��z>\�b��r?��Pّ v�et�EA���<T��>�P+�<�Q.t���Պˊ���S�Fz���s��o�s��G��R`Lv�p\f�*�܄�)�Lj���.������A.;�g�
��Ʌ��
�z�p|0��I�c�R:�cڄxQ�(a�axT߲�\o?������.p�|��~�7F*aA�� ���|�2�v�])_�����q$b����$*����Vvv��t��|O�ku�'�9��~'���'$`r�X�bzK枦׍aNVG�8��B�l�M1$�2w
	x����-aL��߆">�kub�H���v��C'���E��D�!~��
I�(A�^�Ձj��O���S���RU:��%YJu���.�G�6���d�#��?ؾ3j5�Gh&�"+/_7P_ ]4��4�R�g���Fa#��\�LP����f����kT���Z�Vj {G����sϚ��tf�B���N��-��k�|:t�L:�[x(Σ�	M��!�A5SB����m���}� 4�R�� e���&���fT?7�G~�+���+�xC����]��T��b�2�]�����7ϝ�KwFZ��H t����P6��,�������o2a09[5@���m��۩����\�炕{�"\*�dG�?>T�`Gmh[<�;�-���!!�k'�!4��$����6Qj�L95Y*�qI�t�#B@�y���_���܎����
<�0���e@�l4�ݏ�d/'��qi%�%��˛���-aw�Bw���s]��C8�)mdU�Mr�D[���t�A�J�lIӊ9��ҁǘ�g�� ��W����_�X�ó�΀�W�K� �7�Z|���Ɔt.�i���y^ꂏu}?`�	)���!�a�u�Of�7>���r��|
]R������Mf9o�V�k�$J�Άh�6i�N�M�%���2�@p[�ˈ�:����`x�L���]��;����n'��J興��:E�=�}@S�T��$�/��<�;��ebT����#~� ĭĤņ�.����Xl�L���]��S�Ot���G)��6a\S ��M���``��
�N��O<�٨�4���28-��[��-t��p��Y�&�(��*�h͌��}�O�3�&�B��锡(������;�O�=ddv6FZ��LU�)͞�T��G���[�°R(;.�FLe~v��30��ꍷ��bc�h~��������/ΰ��2�LAM��rΞ} �q����i���:+�#�z���?(�Ks���U�CuN.�>DK�Q�n��&jN��S�͝.��4p�,�;3�l}W�hN� }�I�X=�څ��.q=�
�����@JT:Nk3�k�F�ߢAt"z�l�)���2��8��:ZqK�Á�Y0�5�5�ɱ���U?�R��ٙG�_�&97��X(�����l5�4�ê��Q��Ͽ��Wf���'�k�Z`:���N�1	8*)�=XB4��3�	mE3�lq_�o��i$�滾�"K�&{���<X4�P%�/:-Z&:���R�O6jE��e�=�R�?�C9����܌q ���ޮ81�X��b�Bf��m3��5M[\}`ꡍ[�Hs9=״��
���OFĸ�W���:�߿�1��s�n��a���B38������ �k�ZV��OI��]{���-Q��,Y��v�#���'o=&O'S�ዄ����+�O�n����R}aʜ6�����$@�l{��{�N�l�C��r?�9��X��%�n����H@�`$�b���~�2��	ȏ<wN��98ң`�5��	��x�?MP�l%ײ3�3�B�$�e7n�R�F(�<7��M�Dm�ϝ��D�h�#/�dz������Yt*В2ɀ��g�f��sy�b�X��P�D�F>�L>!��a�hK��wjŮ΅z%>y��u}���v�δFb��C��c�)�q�W/	�V�w��?p����q5��(��ޝ�!j��e虽��֘��p�˷g��0�;��c\u�GIPx �Ɓ�����|:%��M�`��ˈ��.�YY��}��z���5W�-�Z>��ZEt7�s��8��r��ftVĩ���!ޭ�m߸���Ƈ���*�{�����K٤�$@�Ѫu.�Xu|o��n뢁h�s��#��=��x�����fC�Y8˳&�-�q��3�qĥ�1������nǙYE�"{�%�J,�c��bA����^!��M�c+�
ܫ���wa�߀ӹ�w�f�ZCM~Y|�3�t�"����H2�@���ܨ�90<�������VW|�l,g�^��p���(5I��G�|��bEEַ��G*>Iz���е�_�RI�S��@��ص{K�p<���i�J����'ׯ��FKlA����jz�@#ٟ��(�����wQt#U[�19�;�B$�����&0�=�����*�`9L
��7�>7ᆬ8S!�{YA���*�u/�ԔXˍ��L{E�;RYk�Jy�n��Ϳ���ǩΔ:�@�� �PWЄ����A7�j��};F=?���������qL�ӻ�7<(��a���@�<
� [ۅ&iPU��ԮP�94	��Ku/�B�����C�:\V��+���q^��|H��WEnBNnǻ�R�uyٶc�p^�3�����Y=ۋ.�]/�6��i��z�_E�d�=Oe�`��	��x�8��'�{� �2zh�[��+u�Հ��v�������ଡ�o������MZ!a�yH!�m~��@��&�$��ƕ��VB �{$X����/�ԣ�2,��rj�I����h{����X� ��{����vW?$����t���7c�,&�Yp]��͆��2}����D�S�nP�[Y@���d̠���=x$���@&���yb����� \��X�~]�@\��ЩWW����@�v���2��q��y@��o d�r��=��r�b�݌�©=/7��5j6�KPc2�� ��'���m��y8��d�`r�f_
�?�\bW�)*�A��O��V���V-�'��G����wG�\r�F�]'��b��P�rH���:�-d�Q�d�o=g�:w�g�:+]%�,�����j��|�������QE89�>k��aʬu��L�d>�R7B����K���#����U�d��e���p��:�i.a|���d��|ж{��?N�׊`rA�3ca���9��A"�;��(3	\v���;��7\?Ϳ��h�ص��\��Ӆp5����?�=���@��?u��{�������G�Z����EOB ��R��k��n@H��=���j�����ztӻ0e�ߧ�H�R&{Xܻd6$8Ô������f��'=�Y4A-�r�bz��D�/q~\H��I�%��08q�s�Y�?��	�$�'X3�)3i+A3l���Z�,i���RO�bU��o�Qq4جK&x&7f�9������g�+gy�3:]�!-��5�[����=�~��[�� �9zm$bŻ4a{�@�O�ό��L�E���֠1���M��h
yT:f���3�;�f�wV$�a��A̽�W�dWH��F���z>�S�?C�?]|�J.N���nv0W9��0����Vr��a<�֋+xKJ�^�b�Dkz�����W/:���eC�ʘ�i]d�E�|7X�d���������Ah��ߓ[}��/R�v�ƕ���i�C�a)�Mz�A!E*h3y5ń'z}-�@@p�-�ӿ���
�G~�>7Vk⭇�[)� ���OX��"f�u��η��V��ui��]��JL�1�R��[ڗ�}dL��h�ҭ�2�s� �d��x�c�����A��Q��+��K�'�B7��=Ry����U��FB��PICgYC��#�j��[���u�#܎�x$m�e�:�D�����io��G�JS��װr�Tʾ
:�]��m"	�3��I|di�:�ӵ}@��j�I;*b�j&���� �-��~�̘����h+T�iik�:/Ŀ9�qh�Y���V!�@9���=����q�tC����Qy�\Ts�'*
��uW�WhnL���>,1��g��"͕l�f'��T'o�:�ܪ}��,$��!�z>�8Ds�Z������%6����q��,���4z�9O^Ŀ43�W�.?����VeI�b�{��Dp�Mo૴/˸PT�83�����=.ѻ����װ�-�g;�o3R��ܻ�z&I��x�V�G�Kk�R,Q���m�+\��|���f���8���<}>�M�}�ir�����|�O63�M���l�J�D~G_�?���]5���:EQ
A�Ĥ#��#�Hk��2���=��u�;�o!r!��Fȍ-v�(�X0z���Wᱏ�4��;��y'un�ݺ��.� /%0��8d	�1�w�:n��ճ:��CK��W�8��C~�rmwDO�~V�2R�Ȧb��oo�>�YA���1�����z��>-�]��%_y()��mZx����D6-��L6N�+-dDni͌sXN���y��}�}�M�H��Ҏ�6��n~�>�F����*c��*�?�;\li���/iRh.�؜��3����B�*��|����zSp�T��	��y��&3�F�����v����J�~~������X�Kj�#��H�Ռ�gь�S���E��~�=4����Dg]��t6q�j��H~���՝{���$�u?=%Q�sdG?�X�k� 0T6�����7�5�G�Tc�[����9?ai)3E>�%<�S�!��|ۅpՋ� ���f�7��#q�(��p+_\�������Y�g�w�k���^�V�W��Z�dQ1qH-x�|�y_��]�(��6��R���������mGmQ��9���������a��q��,�Ec�,sT��{p�dBF*w��Т%�o&��'�_./l�S���7���=���VV\�h��޲Ɇ�k��K}GE]r��mz)3��e����rU���Ӯ�{6���Ƅ=������̠o��h�(�=���wc�[s��������Pn����3��̫s����@P��%4�� ��ݷ��q"�dn�u	GC���ۼ������̞6����C�9jp���PʶF�����A'���'�2���/W�07tD#�RQ+4t�1�d�Y^�	�~D���J��腰}7�]-�l�6����q�x�g���-G�'�VX��
o{����+���������_qU�&ݠ��Aɇ�U#;�����ņ�-�i�R�Ҕ+)@�Z�I�����!����ƿjo�A�Y������Lw�m>�(�5ȗ�ڱg���hq�?�֒�O���-y^iS�������kz���e�'�O�k��Rx~���T�ZvN�� 7r��4���e$�o��bVؽ���SC��ju�
q,�==���(�-r�Y���X�Y��l%Ng�?��c��m����6uꏗ��Sh��GfG�OB�L�
�L���f꫹���%�7�ǟ���=�o���e%�X�c:{�gnp7y��
�ܟN#�iՈ����Wc��#]	��7cɯ�JuC>Fh��/Of�:b�fy���t��B}�4æ>�{\=����+�4é��-��P8fO��/$�}ġz���%�]˙�am�$�����T;���̻6��a;���Ĥx�U� �����iX�#n�$#�7ۼ.�Y����X�S���1����N�ޤD�a����ď�o�cM�\��ޞKէg���+��`��U�� ��R=�P���tb�ڨƣ�j�`s�
P����'t	�5;_p^Њ���d�Zf/"�ݩO��|���璞��G��*ťA�s`E���Bm� Wj��R��h��)�|���u����h*P�Jo��?R-x]rc�a{�=^�ڻ4�I8�I�(`U��E���=�����yDtHA�]ݏ���
n��[��|i����֥P<^�]��oˁ���ǌ������Z��Oㅥ\���rf;
��H���0��~"|76��z��w��ZW*�����@K����ᱴ~�2-����X�s�-�ֵ��vUwOt�@UWr
��'B ��~��Z���QM�.�3E�I?���d'�ٯ�g����ehg�v�����u���ם�fJ�S�%���74���*�^~�hH�;p�?�rƱ�y����f4��͊z37M#M8��%�[�}�{�< �L�i�^������ۙOV�)�)�M}�Y�~#� _o��ɩ��?�����+��e�u�9ޮ=�gL����tb7uǏ�oJ��7\�9\֭\rF?��Pָ�
�Vw�8�2��Nڼ��D'� ]3�Ջ����'�뾉Y֬+�������0�zp���]˘���y�
��z�a��$����{�bP�0���5뀬m��b��n���x)�F��O���$���>�fT�)6������^lx��࿀4��T23}��\EӪL��, !7�^
h�>��=�	} `hqz�v�>|�p�⵴���mSZh�3��vy���O�>;�![E�S���;��BY�j�������%(VH�����|���t���K+F=�l���5E#ϻ����{�#����l��T�����!��8nr�!q>k��O�҅���.��5
Gz����Po��D��q���=4nJ]�:J�ȣ4�T?:)M��du���9�J��#�9q���O&��3[����E����PԞP����⣘8���摀��A_Um�St�6jC���C^��x8�N��)��=�"���>4�d��[�M\��zd�o7�+/.�w��������'�(q��w�c@f��-r�|����X��_����^��\���^��5�Ͽ�Pmb�-�if��k�?�u���h&1�����f��o�CS���g���O�q�>��J{�����]4����Xy��R�y�gP�ފ���Y��POV�@�?�F�j�_zC�ۘ��V3i���|�i�%@�nmS�s�%�9�q���G� N!B�p@�#�*"�>7�	Vo?�s.�FV�.�QuG.W�+|:B#`���0N���?�6�GOޝC�R��DN�4љɓ~-��ZJ�r��K�/Ī�3�z�Ͽt'��Sd:kGxA`m+V�ɷȩ��=�E��1���(��j�1��8[�L�.�Z9�%���P;�N���쵑z:-V���;���`�ϳ����m���Ɯ�；�<�]�AG���X�.���UL�<`�~�!Ѹ�:���jh�^�?b��T���n}�h<���~?��pR��>��V��O�g�����F��k�Uʻ��bB��#�lR�7ɸ9����t�l��tMf�E���qe�?3G�%��p([5<.�JtG����λv��Ǩ,nR3�+q��I�L��v�'��*fa�Na8ԭ��?*��Z}����t*�8�Y�&�l��%����T�y�^v{M"A?dp��o��k�o$W�Y.�܅�Z��
:x�Y1Q^��~�c�Y ]�H^$�y,3��g��+b�߳�����%�ָ�;�<��=��ǘD�{��d����=���[�Ԙ_�"�#�.�AE�
�fi��Tg��2�&��Ͳ��~.NT'7;ΘrXC���2�^~�.�x:ft��C��!�!���G'��-��)��˼v1vk$ k,[3�TY0+[���A��&�����u>�+5jCj~����mg?JVpMk�#r� �����ɵ�����?ҕT�1�T�:�2byK�2.���)���mRq��=�H��8O�e�Zd��Ŗ��l~��nw��&L�����4l�Y�OzH��XY�A1�.Y�H;�yn�}:��}� B�{�J��X�s����y�r�iA��U��b� =�ʗ�������B�Zx-��`��;l��s�ͧ 4_e5�<��2�g�jÊ����P]66$~R�`N�o>����`$��#��o�����m�G]�O<�rp��+��\�7]b!�x@�Z$�rhV}͸�C	�g#NE�tכD���bX�
k����X�t�xb?�ؾ/3 �3Cdx5^�+p���x�&*�� 8]�v�\^��.9)�S�Sї�z��߽vQ��̅˧�MFuA�+��"^�����}=p���*AD�}���.�W�	
�;�q�W�c/�Il�QmUf�W�ʀw�9X	�b�ѱ+xV���PH����ۏ�8��V���R:S�'� ^���ZPG.}�y�8u=̨�1�'��Y}9c(��Q?3MD�<���:UP��-�E�,@��:{x9������w�ۜ�0"ⵓ�gtpi+?b��O��k vo:{���$�&6X��!��m�{�@CʓOm뚘�WĜ��kǄ`��M�%*���LGf��J������H�l� _A�p�Ol�`���fO������>?�p��d(&���̯��������S��ʅ35Oy&G����J8�?�q:�sXӭ����$������"Ӯ�)|g���:��I�5-u�4�z 9����q)��^[�1Z�c�t4�m�v'���uE�ݡ�F�yRK���9Hv����c0�g&�FZCs|^�ծx/E�N!t��ߋk���m%�ͫ�����`a���8�o����=p��>6�Sd�������D�N����~�4f�Lܜ� Z�Y�~�f��������x��ޙ�;h�׽jp�cY��G�͆*~�����z���lM�]�2��ikxV���h��M�S,C��$�'xZ���'E#Od��ϟ���{ͳ���rM�[R���i�j�G�X��f�ML��V��$ׇm[S��Բ�1��.1��em��É�5�����$%��/�[(�{��r��S�"��%�&�S��`���f;�{�߁����~�y�]��G<��hk��˵�nM�yF�|6�vDK�-���K�2sӱı_��~L��� RBɯ���`L�Z�t����o���kF�������n����_���y�����,Z�]��vE�c@�ll���cP�K�k�����W��I�Io��_�jJ�߳?Br�/��EgkԄjT5jN���0�4!]Ya�D�5)J�+�<[P|ÿ���U(�s�@���K<���93l�;�9[�m�pҪ�N;�؍]�b:I���'���
3 ������#��)q���1j���}�[g� �L��8����K�u�!�����`�2�����'��.�o2��؊�y��M��Y���ƠE&�IеѶ��F�o�"�ؽ��E���m�$`�l��i�_�ͫ,J�cB<c�3���S;��T�c�� d(����O,�T{�Df%�LEc���1��مcJ{�M��$��>V�*K-��{��d�J�A�}&�`�{X��k��k�Ҧ�b�B5�W���h�Lh��fq"p�#��n�����EÙU&c�̠&����{lX��Ī�N����5mDlY)�u�{u�Kj��8�}l��
I���z�7iP7�YB�-�� z�q��� ����4'N5���/��!3ިcƨqR�� ��d7��r<��ʙ~ f���|vϛ+�{��,Q���dwˢ�zS;�`;	�����[�9��yMT��$aNYK*.q��z�~׵��"&�Z�FwB�jj���$�T4'�+4|��L_��QLb*zmnXl�ϛ#�Ͽ���+AF�a�ֻ'��6II��r�P+K.�Rk��}�Q�M�}�q6f��D�Z ����u6��Ԓ#a�:��v���mG��4�S�09��Ԭ��Fn6J�-�B�}޾z��L���_�$�3����������6nMj�j)�2�ߤǼ�s\=��o�<�ٹ^��ZG�'y��C��ݱ
����z����%0L��h��0LR6}!	X.�	;��9q{�[z� �A�	X����I {�%�)�� �Ԛ�s��e0�T=(����7���I���(��:n�I�OP{�F�%}�Z|�+�H��Y�����.��Cy���-ƧU�KvQ�EvC�,�zLS-�{/I@�1�\��=��<W�sf`q����;�
��!2���w|-y[ʃ����������t{��@�F.�v�sE�iFj����}�����g��$@�������l��e���{�J'�����F���v�
�Q��O�)�_��=k�z���LM�������`�T�خ�|��*�ՎP�Jb�S��Cz�//G"��
Ý���JG� ��,����]�?T,|�:1k��l}�#r�l&������>���%VY|�sS��F5�*�#j?칮���ĉi�F�C�����8�E�i�����M-1�{�>��]���:,P�..k����.ȹA"?�;��)�N~/�;Fr^Y���l���2�o8��OB�1�P>��	�N���;���}�Nq�x��[&\���.� Aj.�SA���Ӷ��q�F�����6^W���j��i������Q��t�h�n�=o�+z�ƺ�Nv�ŴR�~���J�{��R����D�d�Q%�!>=�`�9)�����c�a�j�D@��̸O����v�٘�+)5=���c���'�rC��W��gy��:ZUF���஌���Ի�aOAk��y�t�ns�B�Џ:�j�'��ѭe�]��ފ`5��\2F�:מla��76<�v<8���P���f&��-ވ�jC#{����_K��Z]<4��)��0���Nu���I�������5�#�?�8(ήTD����J�_��i�$5Q�\ ȝ.���נ2������c�,�4�5g	�n#�8�ѿ����MWu3�	��P#���^���Թ�����C��Ie�]����.O�ɬ���T'��ġ�U���8h���8r�R1��bD�ڸ�Q�#��+s���d�N��~�]p���}0"��C�`O��ޖ�u������;/0"a�7B��g��k_��-H�1���DU���p�K�,ך�W�:��l��bѱ�.�Ŏ�r?�,V��Z�G����zH	��ԯ�R���������'�������{Fe�!�]ܼp^�qz��p�٘(�&�~�'�b�"��&�"����ǐ�m��VZ�ǆ�V��Ӽ��z��͇�R��H��m��"���t� d�J�s�� �lH�+	�:3m���ðDP��Va/���<�|��2[p����,����鰽/��E�q6�o�S�`&��q�`e;?���aFe��F��u��F~n��=�\��E����G�ݑ�'$_#�!������kNH9���q�׈�	�Ҡ�r�L����[	����9��;�ʃ���ߩ�j\�.������zLzF5�?��I(���	����|���O����gHc{
X4��p'3���-YT� 7�n�`nc$�與p���'�zў��"�X@KpM�뺛b�M#G�,t�9�o�Hc�%�7ΏY]��!�D����U��-���paG�K�������$�j/dz�5ԕ��p/����p��~���+����ۓ:u)E�~n����)*�"��31.�.4ω��׵.�3�ũ?�GYŤ\�0q���h�ZXh�ܮ��%4Tjymڼk�G�3�"sg�b�r�g��i~Ƞ
+���|�iFMq[������ޠׅ��m�:���������58ђ���y�u�Y�w�5�:5^"��BfV���J���A��vc�7T��yT�ՙ��?w[�8����?�v���������;����,*�i2%/f�x�SM��0@S�Ĝ��y}��u3���~F7�V<����|u��8�J����Ԟ�`�BQp�t�C3��:E0�HN���b���-�^.�;U:xa�S��5�K[�T�CUՀ�������\׵��%�������:��er�Y��xO6N'���K��4�1_�u\��풅5��pm�{�L��%~�D��~T�h������Li_tPI�a���g�k�Tk���Wt[���#����ehR����@m5��p'r_H�So�P�-�DeM�h��V�#V�~ϠNܪ{�g%x�2��W�	�v:�~q��j�$h2�?6˥K�/�$o�r�:Xq�i����MF<��7���bf����Kmd-��ҳ���v=]g�x��~�)W!U^���)Z�jJ�K�����#:Ȼ\MG7����D�{���$��`���!iw��p���~X[�Ż[+h��ԝ:�%�T���*�	�_g	�3^V*�-�#�ڝ{���фb���%�����,��#��2wjs{4l��G��zU���������h�Z(��Y;���K :��Be��U�-��'L����GX�� ,��m2z}~#_O��O����ʒ���S�L9ޣ��#��a;�Od����zO�����RY#��%��di��k��92��"pB\��ZE�B��֯�N&n)��c�dL FV~�*׼��o���}M��:�˻��P����]���R>?�k��J��u�K���x@qж0�`�ɲl-^�FT��rً�F�[�t$	(����������	�j��� �����|�D3�R���=�9��y���i�ғ�u�,�(��~"L6ʞ8K�Q�痸�/7���j�1c?�#���Y�������9q��Wv:o��h�p�?�^�7�m��l;����,�OoӍ|r���g�U��ܧ�:.�����*(,�����á���4�)X��L+�UЙV��6���\R�<�7�b�\]�ni �]؅<Kع�!Q�'����n�����Wǯ�����C3�lK�M&KGV��y�L��7�4�<�B��5�/�B{o��o���"�?ۦ^\���״b�W�Z���Ip�`��$�X�7��n����Kμ�<�f���2����8��*�i�[7���,��z�����e��k��n'�&���4?.d��7�zL�Q��pӷ��CN���@bRd (be�o�Ѽ/\�xg�/��"��Oi����8��6X%��^��0Hy�7�8U�/񎐀u�W�w��.��Q�����B�T�'�R�x��m��D>>��e�e&|�UAH��'\;��M���=��{󅻎���mFD#����Fr���K��o�%�۫B"�?��H��ɜ�C�*!�i��-����:<��A�Ŗ��5]�Q�cm��{g�t��k�u�K)&-"���%��+`48�?�J��oKʲV�2�C��!��1ǟ�	?��$�w�F��6M���Bj�	:��3A���@ �`qV�����=�KS	����Ǔ���/	��^Q&���� �EV۟��g�Vb*7竁SލNUތG��4Q�b�[N�xԣ,��<���d��s�߅�z��,XՖ���%�j���f�bs��V�bMx�)�%X�'=����Խ#��̅���a�"b�[�J��<E�t�}�|�S���G����a���U�.�O7���{yZs+:m��(��~�Zv�}T��y�5_�ۭƅ��ʷ;Y��x���g�5��y���C�N~��<T��e�IK)o�!2��*���JG�G��e�*x�Ѧ(<�� �9?L����y���&�IIUU�zL���ą���ϫ�<��O�.���Ǳ�Vc�
�djb/�`���OqZϊ�sK�{�u���-3c�ي`"��j?������(�և�%��-ь���j�7 [��rI�.���mO�����[/d��Е��:�c�� �}}��iM������(�bK����.ǽ�MB�yq�v2�d�vY�@���� qG;��=��]���j����[ˋx�>3�￦8=l'�J�Ƙ����z� QE\���P��p5O]D��_o$a�ZMuãs�F�5�I�ɠ��A�q/1����Be1��:��Z���KU��;;��+���|5�g_��9cvxjQ�@F�I�X�
À�WS�� W��7��Ss��l�$O�|��=�� �����S?�5��s^e�r/❼m�u����pd���P>gS� w�LY�Z#N��	t<L߲�22�_]����w̉6�x�89��pu.�jՓ��J���W��� � _؟"n���z/�js�g̿QIM;w��{L6��k	�F����b>���y5��X��똍Tm�Nw��e�R$�(eR29��i�u`�0�($Ȑ]8E�m���W?D�y����1��t�M�6 J��]q�Hm>�;v�+�1�8��П�Hs�#oD�Ԧ���q~�knvؕ{�aL.rP�X��fp����9�KI��˸���g�XԌW���1���R�m�T�x�B�����q%��WopQn�u����Pfp��ٷ�]���lI���[�.�L�s�����r�K%���v���s����Ŷ���p������D�ѿ�A���ڌ�X{T������a��\���l��\�;�aE�+��R��#Ƅ�ʖGBEf�c�s��Z�Qo45c���M�mD��K��_����q;�-Ѝ~1ż�^��[���tXE������֣6뿡�D��%۲k��|(�R���]�5W��؏�i��:Z�*uX!�|�;2a�D�	K���*�U�rF4��Gu�_�=�p��$:��"����kFt�q&�>#}B����X*�N�8���u�)�� /��{Y�K
�y�Й�� >����E����ęny��y�R��-z�"+H~����Z��J���]�#�1��	�jF��gH*�5p�3	(S��tQ�G��ұ�;&��o1�{ǥ��k����uH��R�6��"[�y��i=�<��aNz�p �:=$ȷ0����Σ@m��䔸�'#�n����o�U��b�Uy����S�x�LKSޞ��L����� j��E�HWz�
�RDz' �D�t��Az�i�H��;�{�zEB'� ������ͽs�����n��f�={��=�����b �,��z�rZ�m����B�^M͋�[T}��
wh�1p��T�� �:�:]N��7�H��-�F�?l�0���F���U��hW:�e|�D�{c�M�* ;(w͒I��J��]lp9�&��$�ҼwgbX;%7��E'���� �>�x��_	-�T2��מ�3;���:�t�TfՄ�6��_�R?�iiD�
e�/	�ʡ��P���Wl_g�_[�r�D}S#�+�3��ҳ\��@5P7h�ʨy�IEm)���CDT�y��a�m���Y��ąb�]������?�,�Y;���~�L_��p��5��'7;������\�I�#]���]7z���Iļ�bf���/1H,Q|����kx�׌���C�eb�.�h�.�3�?3���*�&��\~���5�3=��T�<�T��8I�T�&���+Z�96�q8bWM��#\�Z�̻D1j��ڳ�N{I4�c�u��lP��͓>������K]�����Q�C=�Jx3��ޏ:���o�EdK84mx�gӵ"��\�W�#�3n����lfii){��K�Hwf�[�Y;Y�S��n��&׶K:}�D�܌p���t��	~��w�Y�����@� �3��VQ�~r�n���0���´Z��wXA�4��Y���,���j�˹K��隔gb^1���l�W��^hp��K��|lN䠇6L�3��A��O�:�ۥ%�%���/4ğ�����5y�,�7��7E�7|��v	OqW�R�ct*�Lz�U�#fJ���	�f�������X�a��C�M<W���	����[�����UŸ,�(�=mQ�mv�4���߿z?��N��ei����%Z����Ӳa'*Y�W�LI|N�d{�ne�j~���q݉f���R,\�ʉ�:1/2d�L=��`rw �n�ϧ�@3^�rI!�6�$m���u��C��=�ݗ;8���.&�w$t9�������8�����}AZtx"2��>�@o@JSQ/�0�7���K�l� *�H��������.f-����X����4��'�r(��6�mjlX��I[����fB���6�>���b�}IR
q�>:�B �&�ќ6D���tmj7ϓj!���T��N�/���G�����u����8�Gj�ɓ�CX����- j�������x$h��"~��S�"?) �d|�p<��Six�׭��e���_�Ec��o�a�x�M�j�E��R�䥇�/wk���<�]e���K�Uأ�Y�I�������q
���<�̛w�'?�͔�S��*�u��lx�=���L��`�e�y���Jܓf��U<��0��(��rҜq�5z���3y���$r�FpX�6�z��B�����'�+9͸Ğ89jioZ��<ت�=Uv볭���^��P���i�.<nr:H�ϕ�(��ʿ�w���)ʱ_0�!r���.��*��s�Oa�Y���hZ��~{��@I�jV0L�����g�f��[YL��FJ\ܐA��O����]���;@��)ԑsL�g'���Z���0~M>2�`�e��.zAdaшG�a ��l�g[
'U6 �01xp:���	�_���;�||��{���خ9_ч7�]٩.�is 9�iK�`�~6�]����	 ڝ}[�R���=�v�C�U�(��CP��[k� XhG��*9��1��Lӓ��e�^��=u�wA��
�"��u�B�+��Ę�/	DTKӨ����DV�؊{��ޕ�Z�
�܋�KqgT�\���@h��M5m�����S,z����m%�oo��u�;�)+$a����͏W�}b+�`���r?A�x���(�?����%�iԴ:�r\.�>���6�΋Z��ޟ���xcx/����~�
%
��'/�7	���z�[��r�Ed"\,�G�7:3g�����ٿ�Q4�nˢ~���ٻʱB�����h1́tE،����ECE6^���<�N�r�e.%d0aΒ�ޒ.���|Iwd�f�1F6�n�]{�7!�I��,Yh��j����� ]��X���I��s��ae�?�]���I��!�1eh����I��Ct;�0`�ZѮ��cڇߛTI��|t�a��_��[R��DϷ��>�4ŏ_����u��Ԉd����w�W�vʨ�ENx6ї���pS��f�.�MM��{]-؎w�1�M2�L�b���:1�����C��B��;t��K?o-�vZ��P
�B�k�X�h����"�>������r�gq�������#��k�,�ݓk�e��+�5S�.O��ϣ�=�tYc�:%X?>l֟X�/ٻ�w"3	6�
��|�|)}�s�X/T���i�i`p�:��䣫�ƽ_{@�-�=ӝ`Â�D�p3��v��?���_�;#�E���[{W���r����
|�>OA]�C���\L���؏=�p��� `�ZA�'1T��}��=���i��80�?�a�Hj��5�5�-�v�;�@ѫ��6��lvS�~��Rn	x{p1)&$�s����|;~�$��:�ޯ��27I8e���m�k�«SAT�1���$�y^ϖf�87�N�(�(��i�1�l;7L6X<t�_�L�}�*�A�`�R�kj0�c���Zh�ط����v@����G�c�\I����#� ��c �)��&lhn0c��F�.K��/ᣵ�"�+:�S�����J��/�[���,�S����'~XW�����ʎL���Qփ��(|�S��
����L/#PU1���<�p�L��A��E�s6W	��j���#�+Td<�*���)�~���<#�'�I7F}`R�f��O��P������<��1��˛A���u���:Q7��J�>3ྡ�������<�ܕ~�:[ 6��N���^��ta�gD|�Vnv�T]~��*��(��ν�� 2�B�h�}�߆¤���� ���6�K-$em&pJb�����.(C�k����t����N�B�d)'&�z��Y�m�+Ӊ�O��J�aGYa&�*��R����:��=�dv>���{wB�� �?�r���Z��GU�b���8��6��"�f��D����rZ�hm�U�����^o����$Eg>?�tZ�mƙ�J��eХ�`����|�����y���z����.8�$���%8t�Hq��`�}ٻK��Sn���a�5m��9К�}K�qS��T�ܹ;��p������^	�ܘ?��Ήb�ڕ�+r�`�P�ޜ�ؚ^c `���7��?j�H�,NK<������z��\�i�^����NLd��M=�����E�72�����Y���E_��f'7�5����4��̅�S;���eo��n(yB�E�o�#6P}RT^TB����N�d>�>4r�*niG�Q�~����+4�~�μ$&���"7Y_��r�{g��G?th���bBg��E�R`�~7��l���?
K��/'��W�C�r�$�sp35ֵn�ڂ����^���ڸ��=���SVQ�]úñEw�ܴ�t���{���e'#w�Zs1uX�0����I��~'
�SE,Զ���L�Uy����I�~^R���dx���\E�ï��P����E��Os} r�8�PZy��'�TcX-̗�;�g�`CqOgf������ր�K��E��S��k�u�����V�����:���7������S���XAXˠ���JN݈4�,
%��3���k[n�5���_�̊���/ˈ�?Il����^�����-��(������=i�W��z7R�a�c�<��ҭ�)�T��b�}�w�oh̄j�����٪s���]33����|,`?>�P�bE�t�q����V7��+�u�e˕���{� �����]ty&ម׷�d�wac��ߺ#=*%���<dд:4Z�t���U�crx!D���/�\c#�v��%�~� �0�v�g�{������Wi�bVpMrM~��!;T�j��*"^B��o�&XO�ךa�����:ϥc#s!����W�E������S,�Kw5TD�>Ú�/�H׉7q>���{�>�,Ri�'g�� �/]�����tW[��n������Y��S ϝ>��y���
^���Y�EN�(�,>�d��0T��۵Hd�����<&����w|:���=���|q�'����>G����'��c�;B�OH_#B�3�����K��*�\5v���,�^LsF���?͆�xT��6�'�)����w���O��@9���;t2�w;OgQY��9��*�Ł~H-:�i�R=�~�a��eg0�izy}�^u�_�zV�\2Kƪ�����sX+n�"J\G�s`�5ehP�R��v?^kX�����V�7��M�elhi���n�r��+]�:5�d/���:���:��y�+0�ʕ�]u�ƺ�������P��%�����+v��\!��ۧ�%��"��s�*����'�����2�X��+ؕr�\f�W5X�$8����M}5/�)�QB�;������=����;2*��<�u�����<��e����al����OU�5~V��Q/�9 �xf�Z�����5���.h�A��^�Yg�nr�$�uR��q��}�sɆ��:F#y �N�C2Մ��җv����9#!&�6��$�*F�4T���Is��,<Cpw�S��<����c����IYJ!w��Ƅ�d �ob���Hr���)
%X������8o��`�� ���3M���ޅ��^eҪT������_���j2�J�'bĬʭ�m��~&�BG��IT��_�9ܖC9��B�͗݋�1������i���L��-�Wo�?�^�imϩ����0G�DK�ۭ:����"  ��"Q�F�]>�0T��)��$�w"��^d+���⤢Te���)���6殾��9�n�P%� &W�K�K4&�S��5��d�����Z8���?+�ml�t5+�0��Xc?_�	e%Cc�׿��(U_P#�� �R��^1�R���@i���|��15��'j�6�v�_����Ѱd����-T���#E�:��c�=U������>�P<�Ց�,�H��i�1_d}f2��Tڧ��� ��~2]a�G���
-��U��_U
N&Jw��ç[a+i�����Pc����z�3:Kc&���B$��<:�g����Iw$ʞ����5��_�ט<��)r�,�ΪC�|&:�?�s�I�h�l��BVk..f�@\Gn��jFЎJ<7�3��`-�����*G�Քc���*Z�.�����<�ҍ,����*wI�n�p�[^�&p*�M��s�E�����TV�a�Jv��&��x�ɄD��J3�/�UF�zP诤��K�{\���憌a���vR*w~�F
��+�&������f1ͩPd7�\v�z8��dc%}tS�_���n��	��J���U��M9K��y����?���A���M�'Tcd�������� ������0Ր	��q�M�J�$�C!Y���L���4�K^�݌����՞�lX9z�{󛺜5�Ͱ��\��DI�6����$�.�=�D�pn�NoA�w �wU�E�'9�bB�֗��Ԉs=��	����w��Z���=O/��Z:=���Obf�,�~����c=���)���^�:����1����3��1qC��[e�i�ρA;宮��3q�B�>ZUV�L�w�y�J���^����e8���ǵ5�C�}����Ѝ� ��V)��x������XT�����Q%�R��OH�A�(%�����L���ko�0L;��G:�Je�Q/��P�m�&v�6 $8&�7-�.fs�����Q$�?XR[�1�m+^ &?[�M]�����}Q�t���Y�й��-w����4'4+~ M�G}�d�k����V�a�E��Y;Ҍ�&�O��o�>��N�\DM�+T���:���kn��J��N �T�F��b���`�P�����g�����W2!����a�����[8y97�^v��p��<F˖$-��1:���O�Ŵ�:՘E��~ ~��j�����\��jڨD�b���u1����w���_jX8�=s&/|Zs?�J�堪�dGQ�/UH�c�g�@�p��(�-����|v�
{����=�}}A���к3���[��}��S�9.`4��)�?'\Q��_�������L}�?�Z�v���`z�3�[ ��J�����-�3vLm�إ���-���l�ivS�8�pԧ�=���\��wz��:A]���k�Y�mQ��3N��>�?~�rc�hcЪ8��+�������v��'p@b��0X�e��G?φg���;����$J��}я���)��}����EN�9��;1M~�b=��B~ǂ���P��ks��P�/���R��;�ݓ8rwЅZ�,2��4dW����|cN���^���\�P��8D�~�@�����Y�'6س7G�}��~LQ]���4��!�޼!��Potc!�����5X���^誧�Dܧ����ΎR��9z��T���Eǩ3q'��\^R�3%@(�*}��l�,����44y����:q**<D�'�e���������	�y ��,U�s{�u'{��,m��?�ͣ������I �j�cxL�6q_��^5|�a�M��n�1��7vEɵ�A{�g"�>f�m���'�P+���S�	w�e���X0X�s����M����B�r6�8U�Ͻ�K�U�Ubo>C7-���K��X�.*��73���ћ5N/���:Zf�[���= ��^6����j4+G)��շ�+@���è�vƦY�jY3�����{΄�A�u>�+�|C}�� ŞzLr��Z�g�t2��8A����XŒ9��8�(�#u���]&R0[��땏�R�������B�Cjz��Z��Re&��g��;��s���
�d�DPO�%�(%�
�ׂ�w�Yf��u/��e���~��,�f���L|�۩�&����v�Rn���_X�>�H��0�,���S�������nI>�>��d
�<�n��=Q+�5���pg�|Y�A�#��W�?x�G����"}�Z}N)����3-�_Cl��قh_�W�^j�0�G4�W���w�A������1�����29>�{�W�]Y�q� �h;�3]㼯���2�"�ۉ!$X>�0��2�X�)�޲�_sG�v^�XjFc�|�+�.���pV�W���n����-4�:����}J[���ZR��a��@���=�>�vD2��#��w&��C���x���A\��ͭ�Y=Ɯ�h��r8q���
����X}��LN��V�\PU�R�1�	���[
�����L�[h���qc�M�u��Xc��0��e2��u'��?*pw�Y�(P�e�`�3�trt^�B}�T�\g6蒵��d]�����梅4�<T�Ӧ�A���Es�%+x@8ؚ�ԉ|Tv�w����F��Hd���"=.sʨ8�>8��ڴ��Z�G&U�?vha��]FW��Sx��)9��U5��a�(��h!�}QVy����.�Vg~�^T}�kL]^����Ls�Ȥ���e#�۾@/�т�wnp�j��ҰM�ۖ�42q��V��-����-߂Z�\�#!�a�_	*8�e�8]���K���4H�;�E4y*�t�	B��w��2�Q���6�gI��h��
a��zԑ�7g�$�RM^yD��gB�*�(�����,�#�5���ט�I�Ki��,|��E�LOg�d%pj4M�.��&�+���fJC��r^�rQ�bQ�b^��@�sT%�;��Jwe}��0y�9�4��Y�8}�$�mK��$$��N����Ot�OK��(�s_䲍s��"���������|���F3"�e���8��u)�,N^[Z��Ek���#S)�iR�i��u�V��̓������EM�L�_E��+��ێ!�F'��d�2�- q1���7�x��G�L�SI"���ͧ�/��V�eSO�nXv�:���̦�t��eғ��߶E��\���{�����6��e���y�Iᭌ��3/��f\VS���ܜ�\6�UR�L�|���W�)BH�u������c��n;�����Tl�3�n��B���l|(��f�c}��jè�2���֐Qv=��!eY$�C���l�^���w��ut%��J��x�t`�}/p'Cc�E������Ǐ�&s���81�c���)F�f���VGW���z�UZC��X�ā�G�T�ωk }�P�Q�3
������=��7���ƴ)
���z`2=�$~3	܆�T�^�>;:�>܍���Cs���+�TS�Պ�>��G}���g=(/�ʿ����ukX���{��7'���
�"[��Z�qj���&!�O=B#\ۡ����O-��U�E��@7G���m/�D%Kup�6�{�	r�j��~z�6�,����{*��#��ñE�'�g:c��L6c��Md�d��NU�_>����wO=����#?�lӹ9��M$sL�c,���Xj�Pv���#W2�}>P5�iN�3�~��vB�)�+�Ǌ}q&7�B�Ek��*ʲi��]�{^g�ٓRO��TWq�(�B�U����Z!;l�Ԥ"�nc��k���,��e�<��A�ad5J�v+��Ǒf$�zI�l��*�<й����/*��X��e|\{Z~����?��Q2)�EfPX�^��t~��k��{�	&���X�gu��f�~v�������S��g�!�1"P�F�(���P�{
�_��^�-*D?N.b��ѻP'�]�
\b��;������dxk����ff ��i�2�V:8RF��M��:��������AW�`I.�O�h�b!æ��������!(Cf�#���0�}�Q�Pi@-�̀S��3�`�}�7��7�\,�U{'8��@�� �����`�����*|���O�]��?żL�x�"lߏtɼ����L��Z�H�2!Ut �V�1A�g�Ɲ����hJ����0?����E]ѳ.���/Y�1F�A~�Eӫ���® �5g���3�ǫ�T��lr�����$d��KLت?>*w�<N�ڲ���0����U^?��ٯs�X�RY��?���h�����m�9=�\���=��:��$�)Q��O����Q�-�l;˫ޭg����qZ��U}��{��������:-Ibyz�8U����_R��пI�W��tz*�G��0���^l'�f���h��������Ll2�=dO�r=��eZU�$Z��fq�������`�)Fȇ�1��j^��`yzz�[]�읿�Ҽ�t��C�$����>�A 2���\�kDO��Z��O��?�m����K����?^�.e����&?�&n�=�� fO�1�ַ��(z0Owm7y�p)!��_[{���}

9[�nS:����*1V���k}��`��a4��)*�s�c5��dt�n���u�R�G�s=�韓Kh Z��<H��A%&��lbb���SL1+�R��]&|bҭ%�P=dt�y�w�nQ6Q�4w&���|)m���e�+��A�]�����n��-qj������\C�O�_�u�ѧ�1�A��2��
�ɓ���$�A�*�1���6�#a��dEmraZ�g��؅{��� C��H��Y����"B\q�u9s���g��*cf
]�������,)&:� ���l��LJŒޟ�M���Q�G�tX;5��}%X�|���Y0��^[7��k��*����E~��L�"43�Ž��ce&_�$t����|�T�I��ژ�,�me6�[0r�^p��B3}mgى���Jq���0��ιo��H`�\���w��DrR!j�霝�Wfxs�L�W���Oz�r��޺�!i[���S��`�w������7�G\�KIK
g��dY ����߫��-&<N�D���|��SCH���kc^3��I�k6O��j�K�I}�CRH�eX�p�.��nk��&���P��ܹ�$�(-�I�fM|��[e�@|�'�e�td��m�X_��L�|��8߅�<.\�6t����:V
 �m!���C<�2Q���&�D��8�њ-�Xx���T��#�2�p�J6�T��4���R�:-�D��X#x%�nw����UO���ޢ�*˞P��P��H�S���>����������-��t�k �z��/j��	|X�)7��@=��s�ϛ������uRZ��f[jN��hqQ�r�Kh���ckr����-�r0��������.�lE�\����_�"�6�k�����N��o��quD��7M��M�f���O>ֳ=�CW�7�}�/��է_@��;�,eq�?j�M$��F�*�N�F 
��%�}�#YN��/J�#����y�ׄY������)�W�[�����+�5��I���؏��4�_��G>Vr��Si����z�Z��z�z����k��`��Л�aq�/��i��Ҝ�Pk�[�{�����!fo�ˈK�[�@3�妑|�$T��G�C<}��ع!��/H�jfç�Q�x�$'�QOSp���zcOb��c�N�ԡ�-���5�TJy8%����݌�������s=�)�[�ix�2�"Ir�9ߴ��.eMƦ9(�v
_��1^Y.�������`���}��;PP7S�ud/����T�>�
�i��Y�?;B#PE�cأ�
5��y;МP��4��0�";y_༆H�:�M�;O�|H豱Q�,��C�Caa����v�l5d-�_�o��j�-��
�\������}��j6c\�:�͌�#����L�x�j4c�g��?���s�ts�`s�6�bc��"�⾮� ����-���Џ�
��3�2(vM�f��H䕪��a�Ԣ.�./�-��,ۅ��m���p�D�5�?�)p�΂x|���8#���g��l6�6���!6�����zN���۱q�$��9����b/���pC*m��{*�"��{<�3�?����ecn���K�.�<os}sU��=�<P�8��X�"=��*�p��O^��DZM��>��u��#�`C��@���6D�U�U|ZtV��Yz[��E6?�zP0�[��bRC�@r;'�GE$��ޛ��5������ĩ �n��<7ַ�����Z��3������ڔTw�:���Xh���y /�P�����vi��~��?�x��P��x����l�����]��1��G�Ui�*�lݻ��,~�>�)���l���v���6�ո�؂6Y�?����-w��c���
U<0Q�lodN�����H����F��'zҺ�|=LJ8X
�=�~چ�^�WVBk-�> �.�s��ٛ��:�T��E�K��� �쑬���FftP�"�/��u)k���Pk)�"���E;�L�Kn$�Θ����g8:?"�C	J���E��2H����B�����J�����hnr�ʶ%M�+�[,w���'���$}�8KM���Y/!�j7k>�bNEn��%�;P}p���極:�hB_YgWD��5�"v��>s�*\�R��J=C����)2�߄���P�t&-���n�ᦳ���fV��І=jk��¶�1�����>�l@!��0!j�����9��aN�l��+�8�뒯: s�_�:@g#�����a�����e�VMv4�����[D���f�G�[���:|ו|���%Ȉ��dl�c�l��ҸjЩ��oL�?���ɝl��
�z��~�W?�m/�36t�ƀ�mOk�;CbO�屠�>��O�Rv-�^y�o�Xo�����p?ӰB��|Vp�A��:��:+�\Ӂ0�d�v^n���m���h�8]I��bxe��������S�l^Ia����2�O������o\���um�:�s�]�Ҷ�T���t*�c�_|$R���j�2�se���OL������	�r�ٸ�n,+�=-De(b��Cx��v�[r��O-!�����Rt�)��rVeX�B���o"�Ҿ�R"�=�=�L>jP��0̤�͑[��,�3k'���[��c𪪬�f/��{tvrUZ��
?��ܷS��	Ϫ1"l������/���!�#?k��Rةu?��#>��Տ�q�w|�>6I>�j$�24�j�7��u�-Z�Q+�JD���5������ԟ���3��#����������Q�@�)�3�-xn#�i�$A��ag+fʗ�����p3|H�h��DA;̳�{�����dyGJB�'W��X�
�Z/����UM(l���ѯ��<l���	�_��˺2zJ�r-���8�+�}�k��B���a���W=?�zҭح�3�۩���n����&7uL���t3��>�ט��?4A*��,�d�{<��\V7���^�F�I�&�4s%�~ly�{�_l���e\SG-�ے�b*��:�,͈Ȃ�g�"���)�����MG��*":�8[b�kl��O޷ �{�	�S]�E}áP�B�|�S�"��J�"0Ϫx[hw�\��q�}E�e@S�4��g����ݱ+�K�����D�^����be��-��$�0����m�K4���f�ݠ�C�O���%V0Ǐ�P�#D���T<U����O�3;��g�l�R�^|e��oI���X_�0�|�R��A�*��-i�"���t!�R-ֺ��\F��b�M?��ւN�o�f���-�}��),;(��� ��F&9�"_��䭯�n��3f���ߠ���W���t�*˷y��J�]�A�νϑZ�@!��S�;��V�1xFS�g��N���ves�ǟ8dc>�o�Jߌ�W�cxL�Suw��/���H�/sS%��@� }�����ΌT۫���_��j������<h�r|H_�� ��OW,+7�C3i%*�r�*��ϔ���G�e��v�=�	dY�,��b�|������y ��Y?]�mx����Ĺ�P$�lg��"����i]�_gK;Z�˗�0=߂��>?�GG 
�J�_�ã&I|*��kH�rw%��Q��s���dB��ǍX�Yi����@X-��:��n��ˎ{��N���'�4��O?����ވ����$Ѳ��q�yl�āx��(�G��:��CͩC���7SN��	i�e��-��������Ю�
��U�EXB���9��������K�`��f�*+IWm	VGƔ���A�D��|�N ����T��U>w����"uq�N��T��!�|T��"=�Q��B�R �̟q�ٿ���/��9@w���i�Ԡ�Q�3�=2�½��y�
�ڕq#��I����=����3��hbY?o�ʬrS����9?�,Q}-PzK#4�q�
����<�2�i�R���L�1�?O���M*h���l�T��=I�9f,>۾f�?�vdW*i�G�S�H$:U-/&o&y0~)bi;�Kf�Аz�jg����3e�]�j��k��u�Z��b�����ADG	?C�x26�����x=BҞ[fty���3�
B���Μ3�ʞw�)Ƌ��GFg$�f�%�em��D[��3ؔ���F ^�`��-@+]W��u���&p]H�#���1l�X��D�e�Uq\�b�M�{��.kԕ���^���rgÕ�a݆�NZ#F����kʂī ��1J�5"�
�^�����?�"��da�`p�Zl�̒�[��O^f⌊E7��mC}�N9��9�i9D��wE3�ۚݠԕh^n��wI~��@�`i�\����؏G3Ʈ鷀V~�㄁Oّ%�M[;z�~���B;�~�r�-�A�($o�"�9������u��f.��lk�;cRK	�NW�J��QzY�a�1`tek	W3ի]>O�w/ ��/=55�����~����uFh)ZT������a�qH�J�Xg����Q^�0:�m���'��/���+�0��	��H��5�ɖIeT��;e|m�*A*�
��%�5w�y�h�
���JA�$��\fEzY��,� V����L\i�X@c6��#��I.�Q�_b������}�4_��Kf�_f��hs\zO-ߩ��Y*�g�(�D��1ϭ�8~O�0
-��� |�Z��ʛFA	���'��i*6m��::��%�ͧD�MB^i�f_�9N�G�	��Ƨ����j�
~�����\Jhz4���+z jb�[i�w?Zn���<�+��qC�9��Ҏ�!Hu<NCm}ns��/	�E	p��������L
|�d�;W��ݞV�����i8ctW-ӆZ#�|Oד1 I��lR�쩵��9wGm�r$Ӎ���DF�DB�8_O��M�>�g߮~���$d�=]v��\͍�'���1F�6���|�m�fV������e����d�9Irl�����K��w�K��pT�b懊���sY�;�a��_��hP�oe�+(��YퟤB�4Íˢe��;32�:$��&�M)��1�߱�X�l��*��ƦZ9������������̭��,|�����4?����8c���g{��#v`TZ9����ˤ>��U�UJD��gS�4`��L3>R�BebJ�]"�B�f��{$[����u���S�U��5 >��@v�п����������l��$!��5F��*�9DY)��?'�-��?�W�-�)M����5U��f�2��Ţ��L�R�Q�+�ݫ�
��^�T�Й�$�OϨ44��_�ڋo*v�T���>|���Ioߦ�H��ZGӕ�ǰ���dyɪ,t����#_6�̈́�oE�P�\I�.�콒a�ّV-~��C���^e�3*�A��o_�V���b��}Q\�i�)�����]���� �+x7��Q��!�+��p�}VPRX��&�_�MA��V<�w�'X�jv�O!<�F���XH*��:T�S#D+����GsIʢ�����I��|�x-L�����Y�x/*&E�h�v��nCLބ!�<=~��D(���@ 2|q���i_���zV�Z����#�pzH�Qԏ��+&�Bn�<l4_�4��Jݛ����P�,ԯ��Tv�C�c��P�A��R3����)�o�Q��H���\?���:%z�A���EȆ4S%���-u��ƏQ�r�q칧�Ї�3S4�'����f��+k��'ނ��7�z�:�C[�aVaǡ���C	�[�)�-`ܸ�ر�0�"ĳz�u�P��T�̗[Z?�����7^ڀ���*o�M�^��w�u����v1�&�x�(ux�/A�\�࿚1$].}�/�v�ث�����
#Kt���[W�͑I�2��AN�J����O#C�h��@��B��Qޓ��[ �t�������u1EJ�t������PLr����>�[�P<�7���T�{�e��/%�7��Zy�9�
�Ӄ�[�߷�k�nH?���^�s�#��~܀�ɂO�rZ�ב�mq�ׁΆ�:q�&���lH�N��&X����42��u��_���k��7ȳ:9��ݓ���|p�F=��"V�P���T�A��%�.�ڶ����T�r|��2Y�`LۨO�I�)��������{n���>����mɶ�����O���O�ܚ~�a�;�/�� �� ��?����Ma����נ�*�Wʄ���_����AS���O1k��e"+d�9��_�y^J�L+R�w�4�0�E�1��w3���n)vǞS�U��$~YF:ե���ү_"I��l)��}1s�m�fg�lI���&O-9���t�@��m�u��ލ����~rN�&�J�љY�v6.�岨����9�'�?��(���n��PV�B�{��n�ۢ�Q%���
+>���՞��C�9s���0�@I���,��m�k��u�tX�i倊���aCr@��� רϠ�3&n��^q���ܜ�/o�Ο�<]�n��P
�H��n��L&뉍#�~Ȥ���i���i;t��<�{K��?O0@�}Z�E�j�.�O%'$�jnY~xg�)�b����^G��,-�Q$$@/�z¿a��U#?b����d%����#e�C�ܯ�(�\�
������}O������{��ba�t�����L�0�,���M�������
ܢf�Ww*�s� #�Z��}����[K��-�>�i��;q�r*5�;q
������p�����/�[lj����w
Ć�4��X*�������~�#���ew�L��+��(>Gn#K�9K�)E�c~�s]�R��9�q����(;˹�E����5�Β�}N�ϕ��T���}�}���z?ꓪ��Y�U���XgT�m��q�Y�vI
��1�����L��>�cS`�hn�Z��3Q]�^��h����GI��B(��Um�]i} �Q흤��ǵl)F���q�(e�T��+�����ןt�~��_>�~PTȇ*�]�I�.$O�+U���3������ϪRuz�WB������\]���b������/p{���3��/�6��J�Ы

�{��HS�T�zoA���#��H	�wHS:�z(	5@����ޗ��Y3�a�ܹs����{��� �����<T���o'!���� CYnH�����ޔ~�KU��C����^7�J��h�7K=�"+_��<j��:ș�>�|B~$ �	[�In��n��sj~��uo���h�����C�7�&us+��c��Lk�R�?梼������d+�͈|�4�jaw��h����j��%n<���)�����N�G��e��U&x�� ��'�%�
P�q���j���g{	�|�t;^���@�b28'i��*���.Z��N�O�����]J9�<S��W��<����o����bݛ�t��G��GpOB+~�`u�̊�E$��¡����}�+Z*p?�Z��ϼ��ߏ4��^�Ke;
|�Wڡ���v��}~�77�ݵ��I��VW�C����=�ݲ�F���� $� �*��������?Gs�/��M�T����0�0���;��-x`حv"�!4W�qZ��%��3��Wb��8��O�ƅ�Q4���1ȇ�w�f����ۗJ����ԐJ�Ր|�#$���] E�4�Pɬ'�:�X���\g�����`���Om<\�=��vdo�R�.>,C�ymk.H��'�~[�i\�����d�����dݏ��v�o������?��nv���e���s���%1�u˿1_{����(�j��<��F�Dui�_���r�鎮Mjp�y�.��6���Rg�����s�DΨ��ӑ%�kY-�E�V돽�ؽGk'�=�w#��Ί[���0'a�I9^��%�b<a���\!}�n3�d>�:�o7�%eU��Ӫ�:9�k���a��Ɓ�|�+t�O)X�	�D����
�����R+VG��rѓ����3�LKz}G���
g���]�>+�;g�Pϱ�y�)�����D�B�F#��Nu�N��+t�����qo����~��j���"ŪT��Y4DY�_��<���Ů|o�Xi�&�Z�<H�^�ڲ���@_���'��~l�Į�n��^"�ɟ=�������XUt��zη���4%C���#���Oi	�Ɋ��i����y�D�!gWJ�/���I�Wl���@�6�vٜ�r��3�o��2j��#N���|��/b�-n�8�zհ���j焤�wH�� PF�F�����6��_����*��÷QM�7n�@�]q�vw��NOK&8W1i�p�3\�fܯ.�����S�����|K{�Ҷ�'����y��Qw��*���ah9��rRb:����5j��0��Ƨ��� U�y	��^y����t���0�,!��,ǁ��,��������E����SW��@�f;U}&S��e�/��/��$��&;���:���?j�w����+�;�'"��]B��+�8PQ����EH����!5�����@l?�ݸ��'T�$��4�6 �23�#������I��n@!���Ş��p�����ht���~�2]������K��=a���j(;�ڹ�@�R�5�-�±��&8l���p������J�O@9�TӞ:x�W�CA�̭DMeQ��zݽ��٣1y��,ֵmˬSr������Wn�K9Zʟ��8n����2�����nԍ�G0���65�X,و��g%�v�>��aN�+r��p�b�h.�r(Q����=��j��'Y
=�n��E��z=�UV1w(¹_���YY�!����_��<�ʪTu�	ϔ�����%r8E��H��T�i�?�jm��"/��a�^��Fw�DW�|�MET�Z����9�#QP1�{���~GC�4\���E�i�S�~��ev������b��b��S�@J~����h�g�q��Oz���ߝ�������
�7���{�H�ؕt��*��/_������Ě��H�ʃ��L�B)�ɝ�|�	�f�B9 Ow��E�gɺ&͙q�}o�8֥_�*ݲf��Z�c)��iq�Ž�'��=����7�ю����)�BJ�C:�q�˩���S:9˱�ÅB5��F��I�GE�����zH.��~���?���VZ,L�R��Z�֒�U�z��{������v�g���޿�
�Wu�Q[��]�����/>�2�0��IẼeR�����u���M��dou������4��>G GS�Do�9�ÿ;����,S>Bo��ŧ�`P".!6�;��n��5�̗���,�C��)k�1ɺ�i��b$�_�����.CRk�}�2��x�z˄��q<B��J;�U�2J�u����J�k���̹E�6Us��i��\$��5�	|>�>�\l�>�x@^�<�@DF{��5d	vJO�'�{f���� ܭ�����?�Q�6=H��MP��)�b�6��.���d���;�P�~׉G�Gj�m2o��e$��}��e����%�����ށ�{3��neK�a����	O���Ů4����Ɂ���Y5}�b�,v���y���o�ٝ��Ix�����cU�U,��^{� �mL(���+'Wԅ�Spxu��ȲHĩ��^x(�U�����Z�b}p�l�7̸��g0|	�@`�/���=�� �ox�q�ޤ�N�A0j�.�g���\��?��r�)m"�1�=�� �z��c�{NN�N9�'m��Кf�b	�~; �zun�|�O�����8o��?�%'RFh�U�[����e�5{�M0��'�Eb�p\޽��!����A���P���aZ8���k�?��b&%j������@A���F��+E���Mbs���B�w�%}&؆,WV9q�Dx��:��n���-�	�o���:���w��(O5G��U0�	��2��.��9��ҭ���j�BW�Z֨rg�/�w���ʬ}+_��ϵRܵ��:yj_�^��׌T�uY�Z"/�D��������8�/�!2媸�+�/co2�L�dW.a��i��2갊��]�� �#"��kRӃ�
�V�K���sL�̘��F��V(w��nRm�E�{�?86�4�����.ڴ�d�痊���j�1Zn���G��P�h����V�EIί��B<}$/Zz�@����~v�-Q��	��K (�Lb����{��{G��d�dvl�Ow�1`d�+7�|fy���J�����L��0�Ǵ�o$N�6��Uf���*ܿU�ƅ�l��ȝߥ2��[�>E��8����C�5FŴ`(�P��X���Ye�� 6���	���$C{���>r���C���EC���D�xufSU!z8��w�'8�/@������	�sՂa��=�y���LJ���Tvz_�+����y%�V�s��h� �R)Rm)w��V+��MX��8fw�7�Y��PI�tDkm�`�H8���?�Г�<Zٹ�m��1��i�J�^ղ|�7F���U�v	x��ӑ(���xS����[R���;H��eFxD%���Zk Z�Q����i��f��9-���!�x.#Q��bN2T��	^cP]��I�Z
oc����D]@B�x�+uc�q���s�!�}M?9Ǡ� ��˧h�A�!r��!�+�[�G�N���^������^P-h��!A9}7Vx��&�c�+�E<�_������~� ���	��$�v�(���y�֚��~8����+��hPG�wb�p�ߚ����k���US)\�Ӭ�WҊ�S�{8�w2����G۷���'ߘ�ſt��c��k[M������X[ 1T�n�sf_�Y��Z	�������܉�Yy[�靻��P�k1�-�X���������.}�������r�3k!����%��?"��!��"���0̢ٚ���![�91���d���	�8��v-���y�t}��oK�F��f�Lfp�+��A'fa�l�p �c�������7��X=�A��q�K��'���\ �g��Vj��M����d`=��̸0.��3+
s�U��!���dq1��j~=&	���Y�1MC��ʾ�FN80̦s2GAߛ�Oo��k��L��N6�V�)1����B>��y��:_��x 9�r�4���:J�Cm����g�u~{Mj?����1���L��q(�H�ԀL#=g����m�%|zd##��n����/!y���z�Ԋ,���^�lf���n�O�&�o%'&��j�1�f��
��{���g*H!�ꪊ��}�z��#~n��� %��Zm��\��b�
gŏWLBB�ր(=���,Hax�I��8qM���yc�C�4L=kG[�����|+�z�H�����06ݐ�^ViCm��{�w1��ZaU�Z��J+ň�|{�Hh���ح�<�b��������qŶBIa�ϥK ��
����u��WiK�#rcc���ai7�Ni�р!��Ϯ���"�T}2t�8�>�u�3�r	��=ts�ʅ��� F3��'Qd�+N�sḱqn�]����Ǉ��_���䊝�!��|����f�"d�G�������Gf��J����-C��w�V�,��}3�����]<5
M`[�����4m���0v�`��_Y�z$xώl7��Q���C��Ng�=�Wc�EU��� l�-c]`��}� z�S��J�� J��_;�[6�^.�^�ey�B.7}'�}ń�`��<hS�!������KtJ���u7�3^js3iJ�+F��ʭZ�m����=L��zu���~�9�!R���悰�t�]=�O٨<����p%�f������'���z���f�W�H|�l��ۅ� ky>u��S`(7��ʐ�^�NdIH.-�(h�o�V@��YWGƼ���x1�nhM&M��C^T��D� �#�F�`�����]f­C�k�V��o�aasu�7�h�K �Q�������uU�c�H"c�����`鹙գ!�}n��UKm�p�`�z������#;U� �^ބt�H_]���)5�&��F�gn�ۀ���|(Z�D���ԒP�8٤ʉR���!�S@�nl.q�ͮ\~����\�'���!6b��9d��2������j��@���qb��X�|w�1�9ny��$?�|���ۙ��+PBFH�Ɔe��G��p.�W��`���I�����e��w��?�.�W���ޮLm���T���jO3|�gH��И��F���X�;�@S�s��}+7���=`���̔j5G�'�p����A�0r��a�œ��O���h�z��4K�x.I�f�"���mK)�����K�-��ٓ�����1=�� @� ��x��l��3� �3���򘴛�/G���p�bj\�C�c�����(�� ��³I���������9�w���lx]��O�<3��By����:����_�Y�r�g�.�u�k^�����
0ϙ]ı�K��/=ݜ���m��R��r�Dt;��K@�O�[�V���$7m��?��bۭ�#���_	�����FX��KW�l���3h�#�
�EIT흔H w^$��}�s����җK����Y=v���� v�9�1��P��>����7�G��ڷ�dg7Q��@qSz���D�U"Dݚ<VT�j6׳dm�8���n�wo��Y�� �*�%�:]�}g���Y��+�jg8Dʞ�hp	@�1�O`ՐH�����h��!�n�א��֘n�ɢc�n(i�vq���d�B�76�WD�u�4z�M	E��w_Đ*d�rw��S����o}+���<���Fd]�`N�)jD|�-����I�x��+mx�6|=N^��~��p�e�*?�F@>v>N�Gy}��T6/�p�5���|T�X�)���Aoi�-H�t��[���Σ B�ʲ���^c�L���Ɛ��4��4Dv�yU�
>����kZ1�#��1S��4���z�j���X<uvR�V8μ[�1��X}�b���W���m�|8��;a���w	�����Շ����޸��W)�I��qHuX5�6��R�����Ț�q|�>�qo�m� �R�1)�|�XƳ����8^.g6�cc������G�H�5�4n��z�Cp�K�̛q���2����l�$˓7�O�#�c��B����R'q �x�e=�~qx������4>O�&�M&�O�{�SI�ih������y�ss��"/������:F�d5���Xt�ə�1�}r�э#��w�RZI�����TW7�7Q9wp>'�Gn2�XHK�b�uM���A����I�} �X��ͤ'��[0	3_O 	.����l8�r;ǓG��F��ć�@�Y(��cf�³�?������kn�-�AC��oB\"e\U,Fy�4?gXm��o�cYg�o�<kK6�r#U������� �i��gm���Ș�xg�f�)�[ל-���I��d�춼������f���:s	�bt���0P�k��kΖ��(Lq�<lJ��p{���If;�1y�>`i{j.ي��k��tIzGN;�Õ"��.
�<��ĳr�f,Y(�0�o�3[[���X��lq*s	0�W�$�9�
�=�d'طU�@0jAM�{E�����*���\͏��`G��|�����dA;d����dh��L��~�蘉m�t���<���� Y�j���)ǽ��[��,��K9�/�lD�Ί��ﺉ�?G��%Z�Ke=�-�<���ꟊL���~�>s��g������G<�!���Y��s��6Wk������@���F!�s��B��d���H���6vΖ.Mz��{*��xCU�^K]9�'�aL�qO;�'�8k�'d[�e*�	�S�بn���Ț�����g���r$a�d=�~���S���S��a,�d.�{B�o<���T>���oT����۵�{<�?�n{��f���q�{L�t?��W��	r:^�?���ġ4&=���t��x[ f�%�vd��0�.��-�1MU]�/m�*\P���I	��HU׳��څI �D�s\��Ω���疑םS��'+
b�Mt���6.�М=�}���r�L ����y�!k�.����eDe1�'�%mC���ׁ�ς:g��Q>b����<��y�4|�@͇;C1��;�Kow4�w*�\�]���jc�KcZs��wM_��M�>�GAq�K�˻1��f��H����b�{�M�
��i`�g&��%����d��$u��o�7����K��̥�f��᰸~}��/3F�L��n� ���ǢC)]�֏����ƒD=���9lz�	H�`�O����f���aT��60\I6�Wa����˽M�X)��h��'�Fp�s_#d�y>�	4�/��Eҡ��L|��ܾ�3�\������w�9Z� ��5c@�î�B�]'���v�$������g%WWD���۽�[;6��v�#%Np ޶��~?
\55�tG�A�˴�|>��#���w�m��G�;�r˭Y'��V�ٮ[Mb$�*�B±���o'�!s	%g�dSk��X(��A��Pk�Tk����	�|���?d�W)�8�8����&��~9�:�ƌ�[�$��>��y_�c�!�_F9�L��\X�%x�8�)ሃJ�.�U^t�����)cǼg,�EO���H�wgq���Z��n��R�r�l�п*���QS`�#'n�O�"0Vׅ�{P�t�/�n����,ACA�� W`V��Yc���|���+ ��Og~����+�+pT�q���
��:�}_K�0lK��ɷ��գ�
�p�醳��ąQ���+���!.G\�u"���w��LS'6��1�:��y�~;��1D�)%�p�fw����\w��i��G��3t��@�xB��7�n�]�Ε`R�gu����7��ϞDܑ,����%6���S�f/5�K���������۷Z�yH���j�#��(u��nM��#K�щ�j�8�~���IWQ�7WBI�挓�J�f1�(������M}8��[�[.?�ߓ�^�ӂ��K�$�����~�]R�Hu��GI�#��<�����`C�N�z�̠O�}�1�q�%��q�����"4��h�n��Q?j��$.�=v�Ť������������'ߝK�
s�	Y+��Q1
Ԏ����/�ӿƕ��z@ﶻ���~����l����h�$��0M�#�<��dgb�C�+:Qڑ�v�j؏�iO�K�ěL/�<Y���VY|����09��O�Y���<כh��JAuy���Ȑ�׈R
!�GC���&��B�D^_����`�UT��L�k��&��fg����cc���'�x_��d��T�S�{l`�_rSO��]�>ҭ�:9Qg���N �Ӭ�zҡ��w6/���6����N$���1��mU��?�B���q�b'��i"&�ei�o���, ��_h�9��K����yN�1��3ߜ��!%�n����3V�b9�]��*��I�PdI#k��j+��ӵ��v�T�E([�卵 �l��K HOi���\4��^�wR�ڼV�-.lO�X��bD��U5<~z0d���	��4v��74U����I`f%y���a�͜�
�߇��\Y�zE�R*��Ůߍ��K����w�k�?}��!�z�溔e	М����������#�i��+�~?�ӡ)�P��b߽q����F�#�bKˇ]q�S�h�u����W
d7����`7s��fl�[�����Zb-�жq�7�[͸�f_��1>j��J})�7r��'�p6 =�7�)���/7�IvM�ϋ�[�V
#&��v�O�����~E�7����q}p�e�c~�N�E/a�����Ɠ���ڴW��ę\(e2����_JD� ��y�F�~�:I$��� �6-��W'�y951�G�߲�5g�_��H��P�3�~;Z0.��E��o�M�����H�����Z��ٵ�O��tY^��
[b+���d+��:�A�E Q||;[��sh�ȵ_<|v���+�]ѹه�@����W�e��ǼhGA�*5��!����kk�n�&��s*B��$��Ȧ�?�,$l��VĔ)e0����5�v�2	s��L]���e�)g{�p"-�R8{��֦��#��2�о2��?���Rc���y�L���A&V�2td���;z/�3���Y4�*'��!O��%��Uy�������}�Sc�Z:R��X��?�S�EU�B�${H4�R�(M�	9\����z�xT��<N�h�M�#�1�|ӎ�*�E�z�${��Eg���T ���K����_a��!���J��'"j�MF׵g�U��ns� ���u������:@�?�����ña���}Zў��ֽz�7�2�.d�hH��K���P|�z����/�1� ��S��aW�`ڷ��+��ZY��_����7����'��|�u��̏ʐ���L@�n�Ǥ��؞�����j���A��.4���0���$Yǅ�T!�~����z�!�wYS+����S�n3��u2{>w����b�����6	�#H�]a�0�8j0)����8J)�(�I?�/���vYa��zh�vq�������t�$��d�ǿb��FA\ȹ``��6g���l	��qnod�9}��'�e5��ZF�
E�l�8� 8*'��_�=J��NIDɺgbq����u���6
?�21כK2�9a	���
�v0\�N�X�o[�SV��t���v,������J��:�C���\SasR-��o����,3�CU����
V���BK�^�C�rn<�����:����۟D1�Ai�!G�'�/>�O�w�-	w!Ry�����33�w���Z�k�*���i�V~�?m�x���̅(�|���͂;�+��H睁�.b��U���i����ݚƒ��bZΖ2�M^�G�48���Z�Ǻ^�\2�D�Y��׊�B�q�:ȤʽR��n����{�������O��kI��P��w��(ȓ��Nem�t_�fϬ=θ�汚S��Ă[�%������]��#l�&@7��~�_ǜP�<�0��޽*����K���#k�䊞^%�/�:EYB��]ϩ�����M�0}������*0_��Ϗkk��1�Q̳��c�ν�纉�vvά�elh�$�����-��������=D�T��G��C/��,Ԩ��/f�K�A�0�'���gq�d���ޓ���pu���T���-���4��BaC=�>v��I�'�͇3��q�5	��0=�����*���Hs�i����Ȗ��h;���[6&]ڮ|��bA�T~�n@��
�Ua��9H�&�./��Xdm:)�>��DDb��j�s�٦>�Ҳ�1�����o�4��6r��u_�9�8�[[7b�
i �/Z�$�?]Z�����C%v~o�l����w�Qh�劼ʯ�-���Uar��Ćꘂ.o�n	P�^����3���!�#�E�Q�)�-nU�aK�IVtv g`�D�oǞkӟ�S��q�ԑP<WI���[U
��ͽyܐ�}����jsԱ��؋�k�>�m�D��f\wʹ�j[�9�u丹L�� Q�w���7Cg٫��{�Bx�����:8�Y��ݵ"B0�:�e��C�c�;[L1����Q~ɞV:lor�dٗ ���p�ޟ�Ervj���}ljGKd{%�8/�v�8Ļ�u0t��g�@�tZ�5�/46�k}c��"W��;�&;9���%�%�q>�3�[l"���/�Z��-2*�v��o���t���1a�ko�x1�qX�xw�ٝ���ԟfu��,V�T)ˆ��4�p�C��%�ͪ�����6�Ȟ�N�\�����!~w>`i�fk�����5؉n�V�NI���� -�̣a��39��Ǎ��v�{Q���1(�Ul�$��y�-^�RK�Srb�1=D��6��; H6O��/SP�1'9���!f2�	�ס	�����/hv-�E6�kN�o������c�n�Gk��WE�87;��͝{%ȗy؎�o�����O-�� �F'��&� ��M�h�����;]�i��]������/��
�|��gϟ���/oƁ��Aˁ��q�ݎ
X�~�-ڡ� ɰѡ���%���e�>�/(�)Χ�Ta�y�[	�)݁/Kt��3�	M��J���(�C��ͧz�vO���R��{��c�"����,�4`O��1�o`*�'����>����A���(���Y'4��#�`���:��ʊ��hi��Y8��c3��*s�	�6Q�Ϋ���ц�(��-I3� �����7�V�d�.9�0-<�8;�	Ӧ�2���d[�[���2uO:�U33b�? ɡ
c�s&kN�G�v��
��r��~��K����fd�$cu�H&����޼f��ɺ���xBa���� �9
��d�3no<Xmb(@aOp���cP�Y�
o�e�T��.^G�����iY�q\�L.��PI�Y�hǱ�6�a�9�޶�%�'�e7w�����
��^�Ǎ�\�@�%vL�@ڝ����,�ˢȤѱd��n�T�.���W��1�Vל��m�!%^��6v	����a�;�WG��8������ڏ�0���.��r�D({�h�L3"��#��C�@��3�?�7�\<��A��/2�0��i���͑�^�\4Z�H@�ʸ���� �x���(b_#��b&y�BP����yt!��Km��aK��{_�w�܄�����s�q�(Vɗ���o��VC��b��l&[�h6����5u����dZc�������Z��1<U�.��o^��r�����)����A������zf�3�8Xo�׌�Y��A8#�P�c��R�*���!}zq�<2��4���G�����,�W��8�i��l��R4�F�<��]p�"������dKq�TF����W� ��G>�m�K�v��ْ���aI�S+���18��E܂p:{�c�g�g�݀T��~��(��9~�u�BE�ɉ?�ꦐ
D{��=�{�:�+ǹ��׹k��Va�����A��:��&���/**T;?�X����HY��/<,T����|�QBE{'Oܞ�6)�ÖJ����/Д�^��"�qϤ���^�!��#/|�{4��κ'�X������w�T�:�3o�,����ʖ�n��B�^�%�Sk����eڠR��l�9���j6�8��8%p�gV���3�(���d�|g��r�䶱��
���y��?����:u>?
�-�"��ļ.�u�M[���MK^Ȇ�W��k=����穡F�=�}�7�޾𐐣���	7Hg����<}�e�Ku���/���
Cy����K�/����荳��-I2a
���hhG�Q�\�	�ص\�o��� �O@�*n�����E��$da���VJ���7և�����'80��!�d�)f���{�A�XC�k�x�@��'M‶`w�ߋx1Z�J�~b��3׶u/��Ih��rg����Mn�B���w�\��
��b|��0�����p^e	�S��~fZ��K����d��z��RE������G�?����h~;�`8��*ͥǴ>�v�i<�!�4?#�L� �Z��9���,�ůˤ1�L�Ʉ�>�����smr(O��	v����^b�.���@L�U��g�qD|<e�r�J�,�B/l�>���(�!ϴ�Lh����i�}�}`8�����%}	@���ceu����7z٘l+���
�~0�������Q.�8�lj���W�b���*��q3z�DZ��qا��Yv7�x�s	�N�����h=�b����`��Z�Ӗ��Y�����Vua����vz�I,��C�j�T*�o�[oN^0?����7y;�#�f�*bZJ �ݙK�����S��������ASA��K�K�0+��T퐋��_ҕ#��p��?	���/0���mP^ΕsXͿ��~q��Hm6�ovν6n�v��ǈy�`�����{*��~��ɘ�r
��o�����Mή臭Q��gI��nq�9��J�O}4E�p��;�L]�W��ڞK��E�]��׭��H\��wz�*{��g�澅YD\����'M+.^�K�M��p��K��	\^>��Q��9Dc��K@�WYͭ�ưcpͶ�Pl�s�Ԏ���9]�97�	�ݮK ��w���ӕ`V�~_�ٸ�q���LS;o���r��}���$�Õ�Zp�9���-�(��*wC�9�9���bs�-����up�����{ H���X
)ԉXK"��|c�4��^n�;thb��2�2�\�����>!�j}�� ���@��V������xoN~��J7,�����#�[j�C��v|]��x뀿 �+�&p!Uc8"K�lӐ���K*d�ıt�pG��]e�r6��୙m�:�&j������.#!�h܏!4�x�h�^��)�>ŭ?E�2�y���ż�����  _��/9�IՀ���G�E��ٴ�1O ����O������II���el�nͽ�9(�����H��RΦ�Z�k���� ٿ�gK���9[FƆ�I���9�+K+����A�~�O�7�:��>n�8C���O�rQ�h��n�'��_���+��X�W�f�0�Rn27��kxLL���19���vW�"`(��[��$\vr��C�&Ե��G��o�$��p'��v��s���TaMj�snY<@�v����>����e���0[.���hj��	H-]���@�/��:���$����+��Q�2a,g�a��]�Cȓ����#�'�m#qD@}Y����j��`�7}0;����0P��rrq?�q������I��%�ǣ4�1WG��ؓ�hr7\�n��N=�o}d������8�p�q&��XR��9��d�*���{�|DM���8�#M��<�=mo/��F�U�%��W�t`��D�l�� 5�(6/(�={��=��DE.�b���0�����3Д4��0�V�K��͚�i՞�MF����LH]�@�X�����R��%uB0�U�7�in;)���b"8�8� �j v�9��뢁�o���2��x3����kl*���It��� ��X���AlZuN8%>E}Dp���ў�@3DKhE��v��|��P�1�n���=�����;�Q�Sx'��T�I��
�)�w`:�0X[P9f��z��▿ɉ�v�)�9N�͖�Upڐ�J��&|��P���|��=����[���sA[�l�f,�e�*�5�
]4Gs�{'��q�ۻ��޸OO��gE�B3]����vq���p3!d�e�g�G��e�gcĦ�.�Zl�>=����PkH�5���l���0�,}��ޑ%Θ� ��'ΠqJ|`�5ѹ�|���S/	�����P��㆘�B��\��	H"��S^��1��׶�QɃ��|����@`ȅ,�M�d-9+���˓����ck����ǯ8J @e��1��G���Mw\��!]V�]ۨ5<]49A����%�΂�Vl�t�ѱ�0,�K]D3��E�t�E����7�߃��{�:<��	�����~���?��mE��#���|y���,5��Q�ܸ�{X-T");b�3Xُ���Uo��g�_[��Uez���l����P���������yH�& 8�l�A�Ȃ/��sbơ微���,�G@�&�T��A��i��Z�n����7A9`�ɢ������Y�|�ԟdo�]����(�V�H���g� ;[�jG*�D�30�'N(9Q=�8��k�q��V�y�#�ɟ�\Lv�Ԏĥ������j�AKjw�oo:�Æ��lO�_�UޤaYM�}�%���I�(%���?����_<��M*H�ЦF�X���3�������"_c�'"}��?rz�5V8�$���u��?7M� ���]����Z�"Q���n;Ktxd��]��Rȋ��x�\6&]�Z���Q�W��J��yP��oT�}�ހ����wx��)Ͱ�B�6��<WQ�a\W���Fr�
pD�E�c���VC%�:Ξ=C���s�b:�OO�T��/S%|�����$.<+ΚeE�Ӯ���uW�t�z�i��ec${� �|_Y�ŻOJ!�U�l�{��ט ������!O��B�V�*$:RCV<v�M�/퀵��by��2[���Txϭ�I8��bkr�m+#�¥P��,����[ya^˕��Ǎ���S�l�دl$��z�+����`����{%B��o�=�2�_$ B?6�j�հq\����HE��)Y�R�)�fHvLq	`k�hv�Sa�3ȡզ��C$�?�Q�9�1�!Ρ��N���\�7-�|��"N8^s��,OJ�2r�e���!`�m1��·�S�q��;[� U&i^"�����~a�0�u��IA����*�E�ӈYa����\�֋Q��V��?p���-߉�^�3>0$dy$���[�W���"@�O�I�_./�0wh���J�r��B.���w]�r2GѼ�����-\�?{w6�W�3T�[P�x���7鸴�����`��JGj,a��vz�%���c�O�=,幕h�v�o����Lv��	[�I�����"�$��1�	ij��U�Y�c���'�+��*۪ͩ�2_���?�-9�����Ve��.�-A���d���r�>?�����o-�l$�"�h��u�`�q��ZpoH�������Q�y��oƹ+�'g��pC���?���-�AP�� �gx$Ҹ�E4���z��h\Uhh���3�lYh������Ҵ�Ky�C"�j���_��6��VM��B��y��/��$K���y�]�ߞh����o�*8�X�6U������ֶ�*}��Q|��6�/d����q��XazW>{	p�	��.�����~��5�[K[�>З�ݓ:�i��?I#��!+;����YC�7	�$����I���2��V�)�8q����@��l�3��X}��>��ƾ����ŗՒ���i4��f�<p�rMx �b�0�K[�����岮�j��t3�R���W�D��9G��~
`:�w'p��9��!o�@�Coٹ�R�D؟��n�B�F������"Q|�4�Q/c���2f���l<Oj>�A�ؔ4������ё��?$��1Ѕ��T飄 ����c�k��A�_ܖǎ}Fl�G�D�J�Nf�6�������e��#��&0���|�zl�C!	(��[�]*"��@����u��Q�\�6@f�eeP��IC_��+dy����MN��H~ �+ްeLE�3���ˈ���aN�seU� ��R*���t먈n.�k�}��x"X$a��u�e�,�~��>�e"o�������q?^��;b ���7��_Õ�S�%�ܿH&5re�>i-?�Z��k�3��Wc������nD@��ҥ� Hi"%(�DzSZTDJ�	@i��Mz��C�T齷�B�����{��9̇0;{��d�w}��5k�q�V�'�l6�Z���\f]"=��|��~�z ?B��V1�2d9&���<�@R�����a58��Oid��gQ]ٲ�7W���OE������UGe�*x7q
�%���6?WQyO#t�ʋ}2��P�ʠ���*�I�Л=�k>���4��?����BK(v�j��|��aq�c�*�����Å��q^d��f�s��$����e;�Y������2pI�2:z��=�^Zǲ���)��=O����C���ma�����X0ϫ:8AD��/ǀ������?�s*'ګ��}��\��ܾ�n�Ľ��7�L��{B[�s�w�����؏t���5ˋ��?��t��+�|7;E�W��z޵���ex!e����e������z���r������r��>(�y�l�@ӏ|�ch��|K��˽�Ԋ�_�i��<�.�޻tN���V&f��vr�����Ŵ��������t,�a]O�z������z�5�(0u�KB�me�RE���M�x�d����~�y�c�?4yJ}hµ�*_p_>޳�\��(�P���n�ASqo.��4$6�9i����I�g��ˑO�J�9����B����`�)ծ:6W!�L�Kb�.r?��E������gbX+�NF�G��0
�L�:u�wal�xm�cC~8�|�2� }�u~����0~J8�5���뭀>I��q4��Ũ��3?�28�0?x�n1x���z.�72�?�"���!>{im��kr�?y&~Q�2ܷ)������M����w������	�=q�K7�O�;jx��א!���F�(�ƆC�N��+�1V޷���30�Tc�*��6Rc�c���v��n��8/�/���O��B�k�[��ac	uo�o)F�4W�1�H$)�w�3�޺�d�v���-k~o����)��r�'��]������_�F;A]�Ќ�I�=��U@m�G�f��T��" ��`v��x�g}g5 R���=�mr``7����>��0��5�%�:VY�~X���Y?�d([�m�𮲣��� W�X�S��d�ü2��7˰�
���}��Mm�d�.�M?�� $��X���,?&�=��_E�*sN]���p��G��a��M�~]Ҍ�x���_�1���+���A�>�W��NFh�1ߨj9�.���=1��j��U %CL�ąp��-�̧��!�;.�ig3b�9s�bsQX�eC����v��o���B�ߘVn�!]&?�a��d s?nn�?`s_p���D�j��?�"`�,�ш6�����_��J&؎��WN������@
Tx�r[��trҔQOD)����� ���O)'�80�O�s������9���D��J;=�K�lҘ�R�eg`ք}���޲�r�<��\l���x�)��}l�o�:�v���[�Q:pA��8��괤!��6�����آ0=l�scԣ*�Iق���[�;���7GB]�e�6��o_e���y�K&��n>�6�և���-�.�R&)Dm��J��G<��|���ݹ&��M(�]Y�8|G��������ґ9�)�J�+�î|^�qD�����̚���~f����o�q�ߚM[ڼ��́�A��;���X�w�]�����*?<W�f�B.��|�Z6
��}"�����/�kS��%<��Ʋ«ѹ�P������ٺ }dֺ�ٟt�5voU:�y���V�!|����BB]3�+�����	n
cWٞ�v�*��k�կq��sH(�a�����o7ޟ�+�x��KלTȷZFX$��v���Rg�PK{��<�%]�9z<%��I�L��i���w�w���}��
�~��B��u�
{)�ej�0f�9g�{��&ѥ
��';����1c�����^M����#�B�~�!X�ɍ��+PY���<q{�2 L����]�>{�h��:Bh�wW���s���A�AO"�y@�"�=�X���2���q�T�I8ΐ�x����U��:�כ��H��������9�Sh��*+o��G���'� �Db!�jV9E� ��8��p���D�����[UKmoGG��F�J1X���R|]��Z���7��1%�9�����~6�E������j�n+G��N�2�A�+���e/��3��RD�_Q�][���Ȓ���v{��>�0U�����"x}<�l<�^1(Q�{� ��_v��ɶ|���t=�vN���ԛ��n�^O=q�����(o��ohg	�j��q`=�|9�ł����NP�;F�ulp�	_��Sw9H�'�2x�p��&�[��`�]����+����i����1��?�P��r����h!k��ş�x���?�_R#�Y��A��F}�Ԫl�Z/%9�~�\R�,��j�֚�OG+�B��'�
��ۂ~����ʹ/��[ e_!�[���k����ѝW�V��[�u�cfq���7r_�AV?�:�^���֙t��m�;����}�)Eo����3
��%ol��,>�n�[�| ����.r.������Ǖ.��Օ�p��z��cq)�Q��������r�W*w������Q�z]���k�Ԧ�J��p�[Ʀ��p�6���>(�����޴�	ܞ�v��&L�n{��C����n����ѿ�� �yC��P������5œ���@�?�}�9|�b�9S9W�UJ�?������s�*i���Ξd}l�kpL�,j7L�?7팣�[��+����X�|�#c��^�y�3-��^x������CT�M'�\E �o�L%���'��-L�e]))��U�p�$��zKz���2̆��7��&�3U�T�˄&V���}�;�q��o~�ӣ�N�2��M���Q�H��
��&V>7��Ů�.v|d 9\�j�f�ҵV�屸������7���$I�߆�,mEve�����':$a#�|"D��m�7��.���M��>a����ʫ_������I8S�đ �~<��3ƒ�������%> ��]�}�Y�Q��܅�<E���������c	��q��s�;~e�4ω1��D��w_���C�G߶YSDt��	�;O���z }�x��Q��ϩ�M�	Qd,o�C}�0�t1HL�����+���\�-S�*iQ�+� j���!ɵG�{�:���Ћ�q��U�âgU�B������UeV8�
IV�Ɂ?ګ�p�j��L+>���<z��.v��,������N<�Hqs�ۢ`�_;YQza��R�����*��~�I���u@�<��� f92�`�c���xʜ�cuی����	�8���dۍ�����k�q��������Mqad�p�J�f����|�t��B�ǨF���.�]���Є߅Cn?y����'F�a۫2�w�r~��|�����cf"<�"~�wa�.�F��DC�g}n��6lE}-��X�ʎ{�t�Pi�'�=�Ң*��x�ߜ��%h.Hk?����%���]�`	�ˤ�I��>�⁞	����C��?�ɞ.Ք�
�M	xϼq�d�en���~���$G���T�[u�eA;^>�������	�C
#���Z8�xp���`�_�B��NW�(�[|
J��+���X�dO.Cl/��U�s%�*25�c���E��+{9O{]���r����{�h���u��j�����M�Zi���UY؇T1���<xL�`�"�祥|�{ҿnAb�"����K=�{��Y_��ZC�me8��u�Tm��x</�}����U���a�j^d&?�?ণ(:�H��\�b���LK|�zc��ڏɣ�"ǇX�Lis\T�3u�׫�U���$w,\_W�m��^�U���c0>ł$��ѩ2YU����A��*��Ԋ��J�S0�Ek)h�4;�XuoU.�ԬG�<��{�Ϝ���O=I~y`L��/�a��}%��-0��֟��jǵ�,��>�̂��t��̑�퓡��Ihp�
��i����ҭtϬ�[l��7'&��¶�F{�y�](%t`�ӷ2כ��W�W�R~�Ʃb��0^t�7������0��ǆ����N=�1�W �%��{�=��.7�)��JT��j7�k�������+�lC�ŒY�}�-vlM�����ULΕVp�M��:4���c���_�h�L2j,:"qe���Qxq��2�]]�oOW��oc���Qt�{�c���`M��ŉ'�U���GLj-��	�&rUR�������k*��Q;�-�f��Y%PT��\0�C	+o�6UսT+���5�ʱ�� �B�r-:5�P}��Fp9�cov5+��3>��3��fD�{Xƾ��ԝ2@�������6�3`l[b��NTB��k(���ԋ`�.Z���Q9-=~8�BE����爱�Z�Zl��7�>&�P)����w��%�H*\P�R?��(�;a�%���]޴��=�)����@����5o������۾��n�c/�oL�A�A�����x��r�E���H�����8�8bL���=]��𜓰\S�ꂦ�GMy���I�
��_<_�V�e�7f��t^N�:�}��C=��+֡�w,���{QX��3��@���v&�@�7�!V3�{��*�v����V�L� +	g�yЕ'�
�(丗LM�0��=����iV
+���E?�U�'��u�����ڵ���VV�p����)����VKE ʢ���,"���`h"=�f��v�e�>��=���7��dNB
UV ��/��Z�[��4�p�b���ޜyT%����x�s��a�w��=L�W���ɯ����ܜ�m������a�sқ g�;������\P1��$6�ޔ�_+$D�?J��t�_={�4=��2%�G%��:b
�ð&5n���9D��~q���=h���D��%҈ɏ�ȯv�J�Ã$׀�K~Q�3���W�-b�Ywm��Դ6�6�"h��qrU���e�n{��r����^<�A�����0d6���$ �˖j����"���t���Ԅn����r�]H�'I睷UY���cE��� ��]��sJ</����ͨ�A�~�!F�v� 
�C�$w�N�s9�Z�u���R\��Ic���N�!��*|(�'y�J<���y&�H�M�3������ͽ2_�����VA�^�{&4n�z[^�E���}�a��ÏԨ�m+k�[K�������W�ka�������='�Wj���2�Y~9s����r0ֺEY����$́	�T�+�-2������/q�7�97(`���UQ���e�.����₿R��bԛ{5ޓ7�f����E����N#��; �����>��Tm6��"jg|�b;@��|!�Ӹˡ���Y���Q���ڡ��r��^k�Ņ+��\��
�f:�w�5���9�s��c)��5����m5���E9��!�_ݕgT����|;��n������d(>3prn�V��Qm���{l�c�Mu�<�:{���aa��{�4&�K�jF)-���s
�.�_�t��P�T�1��b�m�n����m����5"I�������S	��)���nd�O�_�x�6������M,�`�[=��R�!���D���=�3��0�P�xBBī_z��x�X��"�i��C^��1g���n@06��J̺>L8Ѡ\�KW=�T�?�_ ���tJ��Sx"���ٙ2�
�5 yZ��J�����j/+�p�&�$�����J���&����R��o
ekG� .�:��qy�Qۉ�D��Mv�[�Y�ʁ�*S����T{{+NlӘv��S��`�K_^��z�m¨IL��}��N1qG�����@���@K�������{����z*�'���2+
�ha�_��R��?�ü{�G����āf�Ⲇ�����{�c�x,����!�%��S�[ ��~/�}�:���_�nWɡġH�d�N���������fW��.)sߚP{N���M��5hS�W�c�K�|�x56r9����"h�ʬ}���4���ң�Z6��q����om�pw�i<I_Ŵ�=r��dA@���	�ݘO��>Zn���nvgn�����r�-�Ao1��X�0)�o�͢]Fs6M�Y��1�šЫ���1f��h�n�] ��S �����t�M��Х��M��U<��iإ���Ɲ�;�ٻ#�r0�u8��i��=�^*��A 71�i}��ވ���)����ix�� Ա�=��J�;Uz�Y_+��Kk�{�َ�ѧ֐�f�okXw���;�~��se��L� O�Q)p!~���<��=(���a�n��<��rfEU�����V���2�Y��l�'�J�ҕ^M��~�&A:´����2�9�~�C��C\�UgxDWP��F>�a�d�wn�MM�d�&��&��g��Wf�@�����&������LA3_t�f~��朧;F�̰���v�O2�Ĝ������<6e�Τ�v\��Q���b��7-����$�W�Iԃ�t���,X�x����<���:9�t�Z4
�_
��wN��f�e�{���Ru�c�a%u柫��u��{:�^J�޸�w$<�����f�<}�pdy�@�mHq���N��wq]x�����#����5�]9A��	�i:s�Nc^�_d�J�U���U��H{4����V�d��_�C:�fxQ�в?��F[\\.���M�1����U���8����>���	��P�L�[�Nr�@%k��s����>���4&*����*��PcX�[Meu�G����p�c��s8f���殺�/J�*c8�㔗�9�S7\�q�QM����t��3U�M	q��	�77��O�`q
svy�1eM�	��3��
l~��N���{��w�kC����u#���=�Fǎ�`LqZ9��2�������C6��ܘ����E�����e��_�]�t�)1���Zt-?��~:|<w�R�i��$s�7��{*c���	U��Q�?n�������b�ӿ89�V�`$���\���\���`������|%&��_�M�7�ߩ�!@7�X�/��'Ղ�|��t
=�{�4�Ɯ�t��%�r�g����6���h��A�މu�������l��m�嗗��D+<m����Rax�5S-�l�{�`w:�lф�k����o��d�J���Sly&�Lq��v$��="m/�򫛡WnJ#��8�E�;��K�,K{}POThr�np��8�"&��g˹��6��w��g�)GJe{��'>;�V5mB�ږ׿�����Bu�-~�G�u�`!0B�l�i��";H���<��Њ���G�t��Vq-M�̜6����nN�y��/S��}�F�e�"�7Pk�!�b�L��,�A��;�.!Yj�{֟ ��]0��`S�sT��B}:U�a+e�0X�Ec��e<:�鷪禑� c��"g�����K����g�s����񮯁��[�w>r�(����p�Q�9@��%iΨ5m[x霓���Kh3�(�˒���m�m�Ƣ�7X+<�����8{�HP���<��� ���a̐1��.s۸k	�&���0�G�^�L�����EՃ�#ި�Ga���ˑ���$�#2P-vO��8�'� ��B�G�Z=ɀx�\uj�,jE�ܦzY�[�-.7���r!�<��9e�uO���*��S���j����S��[��__p�й��*Β%�����?�v�M��ڊ5��G�%�5����(4��K�Q��1d8CrY��9����v�I��]��#�e�E�J7R��*��b2T��@�ڸI�F|0�����w���E�=���A��p5����9# j֞_K�q�O=��\�4��;��CpVǶWe�����eޮ����&�\3��2���S e��p�ɦ���v{�Z��`Gz���-~v1��s��
n ܲ�(~���+�%�G��i
�VD�(���Iw�c���m5�o�ݕI���h3X��B��� �w�T����!�򵿃ծ0;qB����G]�~+#��iƨ�זϫs4Rc�8z����j[󇑎Q�k�/��^%�O��	�}Nw���d�9m'~�g�>|����t�o5+��5k*b�Q�y9� ��p��n�*�:=>/9Y��+8=�����^}��
䆴C2��CyBX�?�ܰfI<���"�1�	"oc�=�f4!�9l�~�bK��@Y�9��SJ�L�Չ��UGAg�eLq���u�7����k���.����(_ή�5K��a�)9Yvlq	}۞����L>ȹV��м�d|��O�����ƉgO�<Se�ԸNrV���V����K��]M�x�1~����s�X̉*��>���h�W J1�\����2����Ig�Ȁ��5_�ɛ['��os"��X���c�����_�)��o����%4����V>��58rP�$�R���t���%��@!�F�a,���DP_���X�\u�3l/��=�� ��~���$�i�Zo�%�H�s�0�s!*��V���f�U�I���aD$=��ſ�F��y5�K�2w.��b��>���	�j��Ψ(E �aE�}����%���壹O$�8���Ck��(v�*��O�Tת�6�@�A,ћ_pF�y����sئ73��d�����J�}��Աvo��
���Nw��-���5��n:=WZ|�A�3䤰E��07'���.j5ֱ��U� ����*��Ȱ�/v2`ju�a�^:uz�����(t�ë��ĪJ<����aQRS�Z��]ß*.��6�6:^I'����Ed>�=�
1V=�A4W�T�m�8�n]c�\�N� /q�:�ٮ��?(�_��f0IeuϐZ�D�#`p�_V�����)vXY���ؔ����n�OZ�t�^�	�6�g�Mݤ�8o3��B_�D�|#�f�����/��K�`ض�h�����B��8���yqm�ı����M՘f'ԕ���6�7��b�ײ���,=�FB�G�����K�^ /�6.�l�#���m0�����^���[�<{��PH�c�6��W��)��PN��x��\"yk�8�u�2�IdK�oo�h{���eW�t����Y-�{s�����v��H�.L!u�h�%g5X�9�=��2��Ԃ��+��$^��X^���]�rP"�p>m�'}IQ#F0/��aW��"6�a$Ү���@!�zmW������9~L�׿3U���&s��y�!_t��:虋ɀe%��/�xMP��]��g1U��2П�����/Վ��,�9��'y�1
����/54�+��^#��v�章;4���2>ў͊�~��-��1�+�n�R�����0g��E��QF"a�O�?��w�*A������A���H��'`�a���k������ 0��#y����Υ��+��]7Bmt�	�*p�77�����
[����Mt^ޠYf_i��.�(�h�����u�5ˊ�b�h�����`��~=2@��ia���p
[��=3�3�<T(l�z�@青�0�n@��ޢnT�/�&:-%�$=�����w��qӗv�І,L�O���p���Ba��A#�-�r�d�����w���?ۤ�6Q��:�:���R4������}Z�H����U�[i+�������	˫��xW��M��t^�����Y��9������6��ܟŮ'G!�3L!�;��j��N��Z��=x{ʻk�E���I�� y�8�鲑�M��&,<�� X�Y��$����u��AS�އ�{�*�RnUhbT���%��τ�����5Fڧ�9"\Te]�GO����g�
�C�����r�=f��*�]�ZB���S�����qq��c|���}c���>T؁�|r��^`�*���9�a.���ST��X~�q�O�ȵ<���̛	�B�_���g��4�It������S�㷿�2Np)�R~��\�"���ǡ������z���P�����ㅍr@��?nl@e���%��f��nf�m���6����\ul��r�g��M]Y�r���{�t�h�U�qzs��v-��/y~E��s�R�v���F���p/Unm���t���c��)Oqو�|ꚮ����?�$��=S��{æ��63/�nɖ$H��!]'�����n=H������{z��^�r�n�2[�8l�7�A��/�ڲ��i�ҟo�c��I��0:�"&���yn�bt�)����"�t��ŹlL̊֜�#]��w��o	4��@a,\�N "�������<��˧ri�;�~k������1�g�Q����!Ӳ�/���KJV��-u���R9z�f2x�����������c�S�ēu T�T����`b>��F��z��[�{U��P�v@�������	O�z,S��"�EO6���wEE�[��O�kO�J�~��g;��$�38	�8`P�5�鍻d ֖#5�
����HMA������ATX��D`|e�=�`�z>t��Yu�-=a�q�y�� 
��)�jJ��G��6�^D�{&V@�=u�3S}��t�h);E����}��ƥ��a3�R��T�y�;T�	��5�� }0�n(�I�1lP��� �L�$�{������F�70�w�(�DO�O]��I�ơ)F�8�3=�+�B��@������
�*��T�0��u��Qp���kw�R��Q���nxRt�#��MD�ī3a��P���2ՂM;�I?���['���lY�:xo��H�׽y��l��ȕ����65S�Z�����:<���O��1�86���pa�̀���ҨJ4�y6�J傚f��Qj�i����2�=��ge�������G�.�B9�da�}�J�\�\�A��H�;ӳl�+ok�j
r��l�=�3���];v�ݞ�0�C��p���W�;��/��p�.�Шc�k�E=��Gϕ��N���&�Kmv���?z�V~$�Q�7��(����}��N8�$�#�)��n���(���8���	ӭ���ZW���/nE��t��Y~��ѽ��'�n� �0� ØIH���^�ڮ]���f~ �.�þ=���n�Jj�ע�Xy���G��"Q+��E*~W��W�|fB�jyR�3;�l�3��z|g/�&�S3�F�g'%%D٫S��u��
mc�õ�Kj��'oϩ���0��<��/0��@Wذp\��vI����i\j�dm����4��H6Q>9rx[�@�����fo!X�g��!��)��� ۔k1�`L���W���ۋ��O�Q��r�7�d������kܯ\���d���jN"�d��6M#h'v�)���J֨f�_�S�4�3�{}Q�d�$I"���A��lq� �g*�.yӺ���'�;N�*�]uϩ���meR���8��̕��;zT�3<m�h3$<JƉ�w½�r���^0�E��Mf�B����ݢOң􂊙�ATr`DN�K�����fB��Sv�m�m�a� <�t`�+�}�ꔎ0��s�]?�Z�U�|Y�HLW}H�+�R��NQ�#=���k_���{��d�h��T��Q��+�*�#�m�X͚ ��᫷|;�O�;���w]�
{?:��y�y�-ʟn�g&<��d�n^|����"�#6Z���IP,v�r�G��n=��H�lGpY3Ab�yp9���bw�ٟ G��u[�y��)a�D��2�F�{Qi��XDo㴣�dU2S��7w���QsH`=l�|��!�x��s$[Y+K��X���"���	��K��h���n���J���L��<Иk�rA]ƞn;c�{�������0]�y���j,hI,h�h�da8�=���'�.����/ar���Y�����D(&�����xk�m�2?�+B.�Ź]n�u���c�Or"�6S<Ӟ>����S9P�����Ƕm}�`�^*P��k��A��Tb��_x�-?�1MI<��\}�
ΝĿܟ��+��e�(�*1'�Lо�Vcq��X��o�J��ً{����x��N>�UU܆�5�X��r�f�ׇ3���#i�*�6���#_�G�0�������.���s��I���'���|x�CΓ�DCЊ�v6������Pf�Z~��%����;FF��348႙��|ɗ���d�������uЊ�a�f�k��6r��?�X3�Dt����,$� �/�:h�=g険���k�{W/��<�-7�iw3(r�q�5��?W��I�8o}� ���f�!�=�}h'��]SO�{�_!�?k���a�� 6
��H	U8����c���B"��1˳�@KK�	"�'} ��U�ѡ�G������:�m@=U)�i[��e�xL2�]���8S)�"	aFH��_��ѭ+�d��f��023ﳭ�z=~��C�H�xV!�����C�Ć��S�6��q�,�v$(��`�9~a�RU{�9z̔�ؾ71��I��>�������fiK��h���1�����M���]��4��i@RO�Ue�ru׍Y(3wQz��2یY������<�1�G\O/�m���A3�w&�1hy��[�~[؎~v%��!�P�S�3��՞M��bB-�3���q����G%�����/$��)���h(�|�Tyd���2�ˑ ��9A�!�20��|��{V���)���w��S�ˇ��$��L���%�`|]��_e�܅����W����W��W�WQ�C7V2�Yq�Tn����2��$������ұ�K��}��#���w؇��4�����.�{�4A����G��"����Ӯ��.�l�a$R������+r4����>��i����[�=�G�ϻxs_�C�{�Hl��';\8�Ә^KG���e��Rh�3��K,��qR�������ϧZ�4U�8�1�52�-pď)�#�3S>~�9���H��~�D`=�4_�1��2a��#zJ7��ʢ~�c@�F:�&�@>3��]w�u���SĤ=
y�L�h4eq*����F�R&����Q�c"�����W�OG�Ь�x��O�=�ql&M��Wi��:-k�uuJw�.���*M:R�������[F�e*��d D�m��b4�T؜�q �HM
ݦ�a 6[x�hN���ك��R>����2l�����j���M���)��&7�GQj�5ky[�5��$֦��{��wV;O�����{
6�,kT5B���v�I0s_�t4R4G�j^�a-�:��D����z������R؈�ؑ�͚4	b�>^u�6�4���r��z)�:��S��G��I���I(}1��\��P�H�^�ݢ	�2�J�l%���+�@8#2p�Ԅ4cR�&�$���(���6�M7s"5/��'u!~�dHl0�<�ő$��Ǔ��(��}�lE�%JkU��Z3���	���yA�@���J�)��;�:�����'����N��0a�;l~N��)j�y�~��::�C�r�%�Rz\*H,i��%��و������p��
����Hk�?]F!�Ti}s#�D�F�WҎ+�0(�0zcP8��9�
8n�4[��0�<� ?�Q�v�Q��0<�	JB?��H��-�?&]�u2������.��W��s9�<�:�@n��38xA&�N�Y���b�8��О�gz2!��6#����t��@M
�=��H�|�5X��j�}Y?l�4�B�؄ ��x�d��֦?M��r�y�&��"%i�zZ؁^3q�7畔E�A�@�����U�A�f�(t q��`ئ#�iQ��:#�gd�jJl@��B=�Eϝb�>��r� yz�����h
;bz{�C	�"�>!�9�z�ȁM#��9���F���
6������]���RĮ���;�UU��N� ����t�>s<;pmZI�=*�B�~#]��P��6���K5{�Ne����XY�{m&<��3n/ ���5f�m�����*��e�;�G�O7�3VͰ6FOc��Y�7����6�{�=2
\@�et�H�N` ������۵������YM5�h>M8�ib� �n����1xł�RC,>���zbw �K�3L?�ݘ0¿/;�Uz4�$�~9��,�V��i�<_���ʗJ�������i���{|�糛Q�����	������l�o����7}�|(H��A����_��ɰ�UPWV4I�v.�WT0
7�^e�/t�>!���\��lNR�x��K���c��U�=y��3����{�6�8�LF� xg�U뎥���d��L��kЙ}=҃�?uAU���	��fH��Ryr�C?���W��2;��ʎ�p�	(������z#��GLىj��M��Ԟ���;��7@=��_8����l�7>󽪢�h���0_��PB FM�B�Z�?^�"����ű|��k��3�c�u�+�t���rU;��t8�ivRb���	C� '�2��`<D0�6�qmb���P>� c�[D���q�<���\�Nz�����RJ��l���<I��@��d��(k�R��'.�]�����NU�tyR
��A�>	�	��C�h���ZR8�e���q�F2��Lr��5g�&�I�v�%�
�HB�v�k�#� l�����*(��u�w��9�"(R�e�W�R$`�� 6�G��#��3�S�~�矑X� Ε܃�SD2�sM���4SV;�ݥR�b����]ʡnI2�}��:�1؝es��"��;i�Ժ�WJ�2��ak� B�9]3p3
qVΌ�JpJɡn�R�sy��x�2��U����n_�{����GS�	��G��Y��N	�/h{�	�A��)�Ё9�8y�~`A�8h�܌diR�:��+Bu� �Y���XFl~�g`�֫��j1�>#A��ac���#�����G����u���PK   t~�X$�8  3  /   images/958920c6-b990-4f24-a78c-97ace316bd7f.png3��PNG

   IHDR   d   �   {��n   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��]�Uy�f���o�'YB�D��[��Z,� B���c�6E%�S�֧�$��XJ��Q�Z�h}
�<-�#�XD�b�f�Mv�ww��ߙ���3sw���͝9s�ݻ��/{�ܙ3��|�9�s���"��{�,W�\�r�J���[�%�2����,���"Kv���=�����F��t�X�gYǲ�����%΢��X��fy��,a�S�w!�ES�c����.I��Pﰏ��{Y�ay��Y^f�W�W@���K,og���d���_����%I��$���4�����7^����;�2K4x����7n
�1e���d|��f
z�-7��X^a��X�c����D�����3Kd؉DXַ�Ί֌���;X�IV�Hj��,��Ĝ��E:�p,�SD�Q�?G�ߨ}��BѠ�L�rEc-���s��ɸ�,+c�Ҥ����Z,
�5�_��cq�-��i\M�3l��>��Y�H��W��繐���!����(+���NQOG��QT�Ε/�\8����l�Q*&'bl���#�C��̘��g��#�� CC>A2,���d��1����"��%���Y� y�% �шF���ζ�l<�4U���<��_�9�岘�%�#`�*cj�f�}�U��S B\ځ�6�oPiq��^��J	u��{��ՃS~4��@��n�.&�0eu#k0M%��|�D9!K�(�q��5*�"3?ux@Kt�c-�%��~��2ۙ����d͈�d���E�5+���<2��)�9@>�f�X2���Y��D_���:���s4&�
�~2K������ P%��T�e��JG!�� ��5�N]�C�'���͋�'�C����E8/ЄW�)�+��!{5�Q���l�K�͖Q�[�&(Td9������;���yd8@c���k�:�J��>49+���t$��,��H��.��k�� v,H�T�ĩ����F�S�!�y��`�����&e'S�����}�(�د;!'xh5y�X�Z�E��PL'�b��?�B����W`u?VC1p�ɣ�Q�[a �e#/Q��CsB��/�۩ق�`��P����O����k�Q�΁DX���g�E1d\3�E�a�;��+�iё�zӰ!`��F+� Yy��$�p�����鲿x���Me� �`B�|����|�~�򘘩�u%E�9�C\h�k�i*:�p����h<B �eӵ��1Jƣ�4em�O��)�ȭ�lhb� �I��6ߛ��u�Đ��!d��@�������4;����!�Ў<��hV�&���E�o�v�źh�"�/��ά�Z���iJ���E�/�\伣Nh�0W�Y��U�"�@�Y��\�E�/Xl��g��!~`/�����i0��(G�f��1�ri��b�R�o��XX]O��-RO��"���DZ&�a &���ݢE�_訲�İA�4�%ur���ei�%��zb�@���U���r��t�LH�<q��]�dZb/�4[EZ@MD��]1L��J]�R�h��K���N�����7!֬FZ���*Z�@�h��Y�8��_��}b���>>�כ�t6[�Y�l�B��;z�EP��-[�;_@����}������hk>� ���I>�W��-ш�#H�Jщ�b6��du�%��Yv�-Wp�#�9/tXb��q_REK�zXC�wdŦ;hb�gjN5��l`IA3��(���!�͞�V���)t��銑�`��a�!��u�=y�H��J㿤�u!G�w��,�C7�y,#���~A	A�8�a)�Q]h�k�GE��|��tir�B�����.��{,y>�����&\u���$9�y�@l��4]�i�����]�!.s�M���G�wٰ�PGk$��(�Q"���vZ�R��zL���?���gĊu�GGZ��&&R0�J����R9/�Ē2M-�wş�|��kJ.��\O��x�J�#��D�S���l�@��I�ɫi��7�z,���C-�&̍�oT�a���)��� B"���I�&B\ځ���T|��#�TyK%�JFPs��
3�����n!{z+?í��Iu�Ι��|X���<��M���!�	�۴��w��1S:&!���G���$�Gz;��8� 6<#ܑ�;l��'@��
q��cg���1;A:�n�J��̊���}�خ ��k,�{�X�4��I�>?i�[ly������3y��Q1���4kE�u�Yʑ���$��Z\��5E �ɇ'�)�k�[-Z�(!�ЬL�Qn,�m�ܲv�A���_���y\��fnRF����:�^2X�Hv���.cy���x}��|AB*��N�����31/�ݡ���6B41�1�S���RS"m}�cڠ�XbeJ�d�:��ɚ�V&$���4� !��A��{�A�Tl�������"(��T�&��Q���8�D8�Gw��z�
Ŵ,A�$�R:��@D�m-6�J��T��ibT���I�]b��3�"�?2][^a�
�#Æ���"�����@
̗	�e��K�`��_�u��d!2>�r=*?��ۓWvS")�*]��*��C�cT��3rrh�hd8�df�.!L��,=х>
�I���>=�>I�����
B<d��e���̝��+��] d z�L©{��	���?7�" >bB�.�@E��F��,�,n4���rY��a s���h�*�T���w�B}�~�%�z^;�%���@T�}cS�i��2���oNx��1�����f�(,-I��C���$�~��t���~����D��P�㝎�=L�_�?�qoR&ģ�Y�S���S��̹�-�^����{k���g��烀�	CD�}.��d�k-q-���̖��lt�b6}y�<��#���J�.��F�¹	���` 1����4��aqf5A�>2��4�C\7�3tp"#*�6.4�-f#��1�ׅ�j���	����S�¿a��$'pWV\ �S�cV�x6]F9$�����q?��������hb��s��:��d���=����!��wy��7�+@����\��=$=�(�9N>��?�e����a9Я�Ͻ��Xu�h�WCnd9O�֍�µ2@@&_���7��$�|a��vT���
�^"�����4��$�-��h����x���&*��W�&P"����c�w�o�v������Y|��(�b�7��6Z�,���b{Y%�OY~�D��{)��E�U�A&ٟa����H׊�+*40)�"�Jk��k_gM�O<�qkȵ,g:_�@��;9��t&��G��n�ʛ�$ىN�ѨA�L��a:� 1'^�7����7�0c�3|��}��f���O��k�{�?��ڂ�l���^A�:4{·��D=1��݃[��Mz�,�x�\*F�O�^/���	�Wj� �↪q޵�)� %��^�D̿�w�޶��t�!/ź�}�t�Д*w3����0,�X�a���g�j�6g�D���ϟ�s���Y"Ok�'-σ`n�WF?W8^�q�C�5Ւ�]ۀ1Q�.r����F��!3��^��6˃��6�����k��o�lZ�A���WX"0�x���h��#٣�E�]��+�\NUa?U˥�j�Ŕ��D�wn-�K�$`��Ti��L-
����ihX(��P	�\��-\#�}i���Xb�pX�)���d��$�@:�3Q���9��v0x�b�Q�qL�����x���}�G���.Ie�,���L�	b4Y�̑!֐��"�:\N�5I����B.7�h��Q�@�yLB[����4�2�2�3n�8��d�)S�ӑ�I#i�F��-��~���/ɏK�s��Ig���7���׼	��E��i4����Q�[���e��!O�M:��pt��a�vVt��ͼeU��6�P�h���������J������"��@��r&�"�X�0��Sn2xHAO#i	�(ru%u:wu��<�>&"j�\�loG�ϟ���������W8����o���K�v�Uq���ʎj�3B�uE���������E�%�����-�5�D��JR�Yo�`��D�����bI��c���\��sڞ���7�})+�7��֚!������t������'^�S�dM2)7ιB$lxH�sN��F&��DT��xF��\�Y����Y8�(Y��T�d
�[�7S�4�tњ�s�}��i������F�g��ȣ�nWˋ3냿|j�]���V"�`-sq*:u�\*h*l�>~i��93�go�nn2��#L�Eo;9���^��$�o��(��z�^1o?|�B�B�S����dr�f��"L6�n}�B��y�
�A�>�YVd8@�W�s���W!�L����9j��j]�!+��/ [�p�]
!�
	`�'���z뭴\q�-�Ў�l&Y'��LL�B��%�V�	�ܹA	I���o��o���͉�-A�N��Du,�҂��*�!V��7J�Iʻ;�
���f&��:0�����:��[��r�ݡ��AR�`5B�@2X�w6�Aj@]�Pp�A��E�����B�@���{/e�Y��{�!ϳ\����X>��-G��"��R�� �i��RH�͏���LˉW�`sS�b�O���Hmv	|���z�<��JhZxȀ��c�I���@��X�UH��{H����>�ҡ��<��`2�mR#��i�-�of���,Pq�; %g�"Ac����Y��|_��5�-�d1�|B��"�B�X��E�;ї4)2���!%����a� Z� �8w����@���(��k�r���Mȿ���u1��R0������\@�I48/���/Q�\�}�_A���&J_`-��M����ĥ�~����� H�B�x�~��i���n����B�J.ER<��&�_1y,�~�}@�� �bї��:`������|:����6��P��S�ǂ�]_	����Ѻ��;�\2�߷o�����!�F��}ރeB<Z�U�Kɳ�[d���U�ti����r�CL�*p���x��xH���L7���V@��4�$����nr�x���B�������\^7� ���R��]O ?R�{I�邁[���ظ�$#���_	����k'--\�rb�`���5�@�FYUC<�`J�-�����I�7i�r}i�19�p�s`!����g&�k�ϊ��5`��͖�܈�uiI"(C9��b�^4L��Lb�d�Bư(�ii yU�
������X�𘁔=�``�B��TK��+I��L-�o0~��}�����빦�������@]=�炚�8 ��I�� ����F�G\� A�TGW_v>�Z� �����U^����]jl\�x=,���5����1b�D��3�zC�C�=��~�@�W�e�B�\b_�,5&�&Q��@PBT���pǼ@�	�m�b���!.��5Dp��0�G��e�B#u�}�=���B�.[P��-,�S��O�Rc�M�ףn�U^N�,˻�_G�ռ=�BB~Lj8��y\7�	I$�ϋ}�/��v881��PcktU�ˠN^
z�oB�l��t~X�R��$p4�q�h���p��nVTLn�wz%-�m5
��ur4��*�`^��DH�0Wq��)�p=�$��>B�1��U�5���P�UB�I��xP͓R����LC%�J���'��/���"��aB5OJ��?T�
V    IEND�B`�PK   t~�X��) oj /   images/9b962a8e-14b5-4317-8666-1954827ef6fe.pngĻg\S��=�2�
��>zSzG�w�BT���	�����N@z��	��^H'z �����|_�{�?~��疳�.k�}�1TS]��������\IQ���z"�k����Hg����\I�O��ߟo?���I�Е���������:�� ����������ks"OOOk[W��N�<�.��(	Z"���d��x�m�{������O��݇D]kg`%��1�hU�O\dq5�Zl��|�M��l?���c�0*M���Z�ZwN��a��j�ߕ��b���������ad�~���ޒL���~0,�Ƈ�/�7d�|��b)���_N�;��3H�xg���c�AA⿏eri:��>GB��},��i;�w���J����S��E��ٮ����G#�%�ܨ�1T�{���''=���']|޹U��]�b�E�џ?*�������W 
�_@�O㩤0͌����g��A)Z,��m��ąO�s��V��I�k9y&�+����u���58����|������U�J�t�ر�����M��/���;T�1yD2���k�K�%�$Uf�U3�W$��B����K��"T?ϗTa�:�
m�p<k$��W�����YeZ��<[
�7.�����5.����/���y�_���L�܃A����d+�̿��!s��!s
�W�B.�@�r;Ku�&bt�����4��E�Y)!S�!��,�c�����aAX�J����e��[5y���F�,����f�i��x�d!H��y7��<�_�Mv�N�Q椽�Ѹ^y��-9f�q�~�q$�W�
^5?�]�?C��5(��`I�VZ��4[7��|���H��[��S�M�_�ߞ�x"+P�
*w�M�n,5�p�?��}���y{�|y��omj��M�z���4ŉu[_��'u��}�f��!f=�J/��do���{�+��鄩A��bKw��|�1e�&V�~��I<G��t�1[ˉ)$���]w�ޝ�.Γ�Y�"pi�s���O��S���ſ�2�Ϳ6��]�F����n4JF�y0lM�C��!�ު�(�AX�o�֮�Ue3#y����ٓ��2<�`�;�C2�Q��J ����N��c�u^��a�&I�^7 BN��pJ�G��i���q��	�j�tǉ�z*�?v�_� 5�[���W/���)��6mwƌ��%-[���8�.��'7r���xћ!'6^�h �����g��NS��%gvu�sώ��.��7'$���J�L��}�S�/�}ٞf��|�kb�W�)��ء杜�>v�zQ{P�uoQ=�����d�ꃀ��b����uM���պ�X*���`g���s���㍋�G�G]��H +K��,�	��RC�T(��3;��Wτf1j��D�!�%4[l�w&�e+�:��zI�^5x�2y�A�9���7N��e����-i�w���[���P�Ն'lE��)$�ɏ���S��0�a�!m�� �`D1�װ(\o�xoz力�׋��D�߁ԫ]tg�g؜!��C���t6j٤��� ���Z�=_���c#�_Q3��}C ��$����mD�$~�-��I����8 ��Y��3( �s���6q�\�1m�Rc�B���Wu4~��Ū��h��2��z�(|+�q���9�h޷�+9[]�TS�vW��e�Jr@rB�g���/[a�W�1Z��������DeL���O�OyD��u�ԁ%2�(�����{�F��lk��L6M]��8�z��T�B3�x����Ⴑ���gs׉ߙ-�^�6/�r�O�CV�3Z)�]s�P�!:�۟����C��9j��Pa�2��l��j�b���Ml�	��'9E�v7>�o��V�1���u*!�h��ίޕ��	2_G����v����X����D^��l�I�YH����z�����Yr�I����g�}Ӫ�a ��c�Nb�wO�ݝ?j<������Ĵ�ZN�]`�
(��3�i%_�F�s�� H�U\�fz��kw6��w���fË��9}��X�Rx��e�y�d'-�� ��!��;��JL}+�����S�{9<���a�0%��i��U%/�X%��T#��'���䡚��3V�[��)\f�3�H�y�Y<�c��j%��o���vR��F�4�=��K����,�ұ��؃��`�Dim�i��b��nNT�d|@yLV&T�-<��|�K�1��#�����;�W�s�^���]p�髀K�ـO��.���?��� C����kLLH�#N�g��oE��NF���|�e�����!����	�W1E�!G�%�^=;Z�f-2f
�36��.{6N�}�S�;��V�#�A��އ�E7Hx�"t�t�m?<_՟�?��D2AkMb����P�Odv�.r���c�"�x/��|m��A���f�8qr*�����b�u�����W3%^L��[8�Y!Z³kG�7k~ز
�:�S�)
�����l�c\A}�����L�׵�o�Ε��`,���|/��K�G]צ��h�����g���s�f,��4��e2r��Z~�>�Do��6�C|v�g�u뛳��tb�CeOw��]�c���/i�t�L�N��{�7+?�pя�Y�o �W�g���u����&
F�fLd��o^����>�_>�����Ċ�/��Y9dg41���w���:J�B�s��XG��+`�<�vp� �Ê��2�&����!,��nw�P���ك�-�|���n3�{�����w��|:�n�Ȟ��i�~ʑ���;�l�}6)R۹=z��EH4�_��W��'�5���.��A컬�l��_�p�}�����'����ض�Lz�VΥ�/����ƌ���+��J`�hZN¥'ŐS�f�M�ӱMz]Ig�Y�8f��]9M�Ư`�SR�`l���pA����\����u���M��#g�!H���Sy��fm������CO�-�����y��U�&��+@e�Ǐ"R�1�4��T{{����LZ��Z�ж/��}���#U���m����:՞��g��ɫT��k&N�詝O�#z��"{!�زw2�n�r��<8�c�]jǼU6�r��r�>�J@n�W*�U,��|�i	a����˼��oB��~|I�X6�h*k:���݆�Q�G�M��P4d�3s[p�Uk���qc���X��ں���cCs�J�x�-R��tojg:wt��f|�9=�c�a��s��J~�RWs���E{"U�G�����t��tj�*��
��1ũ)��1M���ԫ.=��T�㙫�
����q���H�-u�H�0=¹@ؿW�Y1��JK�:�"��J�\=LJ*',=�g�G_{���I�~l�b��w��G�\��Vk��=�juڡq~�˪��:w�q.��&*XUz�"�Ķ����ι~}kI
�w�2�^��>5u��?5}��%N�*�@R��}1x ���4C+�c�����i�Խ��*/��3����O/܆�7�[_��W�).~b���������72�}_0������-Zluq(���*�Cb(!���G��.8[�~��ɑ'�y�#�N)Sh0��wЦ>��� 9�` 4%�	�m8+������� ��W(��Mlg��f�z��D*�-�ӗ������>t�5t�IO�]�v_w��DA74K��u���^m�1��q�6��xp�'q=%����AP^ݘ�ݸ�nt�t���t7e�Y����^r�]n�b�f��[�¡9�o
����8^հć#n�w4��*�}n(���r���Q��U���i�����8}k㟜o�ש�>y��,�;Ѧ��b�y��]z)�����Zo��n[g4�zٚ��ܖ��i.��[8��L��1�r
&p��{��2���/���k��G�I��%0R�ۘ]� f
�}jY����9�a%�2��]�0�Q�������k|�L��&�Txlʹ>��t�&[Y�ar�}˰�����F��q���L&������;���/WdГ��Z&��N��|�d(j��-b�r�^Cֳ����ܖq��V���|҉u�:>Hf*��e��벤�YZ�3BS�����|JQ��!�6;^G�#�g	>�v����L��yºL_�,N&"�����u�Q����V@�w! �������m�*1�S*,N1�g36�B��J�=2�o����/�
��L��}H�����\��+���������"NwC���-@*�+a���&�({� �����x\!���ԖJfc�ݧ"lL�J�R4ob�.��}���I�d���d{�DB\�l[A.�k�@����0� u�D�	��y�	��	w��[��^'�r���	�ƎިC���Y��B������/���P|��t��y�d��Y���)^6�{�:v@��t$��|�-�&.r��>� �L�zGjv}�	���OgFq��?6jF���)�
��::ߝ�^*���Fz��nOn^�8��W.ǭԂ��0L�:Q�7�<�~���7���t���эh�I��?�@E�?�o���v(:�����5���󼳈UW��P��Ʃ�8��~��h��YN�r�Mi��BNW\D�m}�θ��a�c���������}�)z�l�j���-��1S�;ǣ���л-�`"���$�.�x)xi׵!�rf�:ޗ�vhVLdc2# ������qiݵn��C����7"s�#�Y������lR�+�0)�Cݷj�yK��I���TgҮ�䮇'�a�׭=Z��ўL;⸕*�����@�ƛ�~���-�-&JL�ĺ1�bC�D�r�0�%��~�g\�3���=0�o���=}JEE�ǃ�3����'�/�p""mO�6K��((;;���ar�瓼�B�r���^k�����7���?�\&FIg	|�958*��Jζ̩�GV��!��8�v7�i�P��jɯ��z��p��7}/E�A�W�y����ѭ��D8e�S���1�]t�|v��w�v.`/�Un��;�U�P����2�d�����;tH\R�4l-=l��dZ��(��{��^�-��2��(���0��0��CF���������J�--���޷�_h�M��I�ޭ���y\ ��p�*a�;z�K�G���?S�B@&r��RC˟���v�Z�$�\v^��I�܈n�;[��W'n�~�@7�> �b��4�Kdq��[�2|t����蹃^��6�JRp��@XES#���?G��:�{�*/le�W����yI�u�	�~���VXכ��
����~Үk���['���1_3kO(h��4�Wۍ�$�ac�|�>e�  Ks�����'�c�6w$_p�1���c(�����~Y�u~��i)lG��k��&w��',���B#�ё������m�u��D�!)�]� �>�Z�2�>�fM��-���d+���v�����+��(��S6�X�B����"zLycC�рLm����7�U��0_��l���~hH3��N��JD��1aP���}[z�W�^x�Rt�;��<g��2kS�V�g���W�yꞶ4v�;�\'��w?e�۱�]C��{S���17�Q�L�����	�Ļ�y��\I�y7F�)�uk����X�D7׀K��
�yQ
��ρ��rXpm[[����$|<{�ߟ��:�S- ������� Pe�'|�uF�*:�"�6��h��6��w����:��=1m�ß����-��"7AՕ���Q��/��s���ve+�/JԣM`|��f'��@����� -��͎̀����!�w���'�$�>@:= ����F�Syy�3��D�\	���C�ʒ3�� ?_�U#���g]�L�2��n�~+}��ח8_�o��a*�X5nSD�w��s���g�"��~�i��ްO�mLs���l��}�WyV=�^���(�*��c�Yy� g��'l�Cl�M��X>�U�.�\C��+B���hi	��v����{:&&�[ȭ8UsC�@�L)�P�6VV�<��Bm��y��JߑXXі�`x^Ͳ�Ӑ�~���x5Ke�޳;�F�	"��k�BGJ�,�\� ]���b.�aC�ً.��s�0��r{_��8[� P\ķ���������ʠ��+���f��k�a�ݦ��!Q�⏐
�pAMދr��k�&��%3J�7~�%��f�n���ښ��.HI�U�@`3�[���޷~���9Z������{=��۾�i�9�s����k=<�7���8����;�!�~����\g �D�筕����~^ѧ��{��"�H)l��h��O4~|�n��?��d��a��HU]�A���L�k[�]���_g5&�V�q_�|��S>g뭿��a����U�����9
���vp={��O7���u�ѯrarّ��ѓ��2[%Zmk��_O�l6-2YTD�f�W����g�+�q�w5�~8���8�nD]�V�Gv�3"9�,�M1ar}��m��E����"�{Y���Q����6�U��U�,ܒ�#���t\�dU7�`f��ҫŴ����0Om�e�:77��OC����$W��=����x��{ �X[~�2�f%�8xO�X�[��-ADV9o��D��%#�G�\�3�LR\V�c�N��}������Ís�RuY�\;2Tb�ǚ)��3��V���I��
Q��'���5���F�&
��$'8�f���A��ɄD�ۑs�I'��𻛺ƵVJ�M�?��U��Ǜ'�1Hp�<�Rݠ�U=b_d���)�Rf_�L%|�`�=�]���,�+��G��&��F;5�,�Z�I_X+q�Ln��ޙ�~�|����vT�5�S���v:�P@皂�V�>ݞI,Iٔ�"��%塡ɬXNgh5�w:]ۢ��A��*�*����Z@����H�L�;Jt� ;[ ��4m���N��6y�U���kq���7��������8��3�m?l��'ޞ���j4���g���b��s�U���97�|���`�{���2�1��]L���)�6��k,��Ї�:å�ۂ�<U\*�55F@�3Y�_\T�g DD�a���ɋ�����\^N�.	���^0�^�R�����L�c��9��S��I��}R��ӭ����iX+���~�n��˵�
�/c5pgS�r���9���e2��!�=�#��W��j������r�]|��>Y7�\V����ɪ����[��m�J����u� �r��@�1�6�1�ĦX�<��`�e,2!~d���ex�b��`�ܨu.�{�h	�2�9NN?�'�S^B���wGa���3�9��ɺ��PBo�9�ae�Z�^8�(�``��e� m央�Q�G�T�a��� ܌���Gg]0���^!���k�+�U>�kvWx���l)��&�X>��j��7��e&�<aw L������>��!���S��B�m��G��>!]��ʟ�j�o/�PQxQC
e�/`jS	?;l,07P�5��a�ѽ4���o��#P��bwȂ?[�l�q7P��'H��G@���_nشS�FR�ZJ�[v�vO��q:@��u4��8�3�4�z�f�����\[S��\YCW���0T4z�-�U��J.G�m`
m<����e~LoN4 1�����5��j�pj��#j��x9w�C#SA�����
K-�xN�.�K�i4�o��(��D��٣���K �dP��Ј��{6��@���lʞË�7K��*����@������'������:�*�mp��^���L���Td���
�u� �n{�f�j��)�;�d�4��Ƚ��6MQ4�
AO �|��\ݸ����lD��ig���o���Tk�&�S�q�ǌa_�p��Õ�\����d��aR$�buچ��]q	,ݏ��4�6�5އ555��&`�@��8>�.� ��>�N鮸i���Y2�iP����c��<���p�l��;��&Ӗ��=�	�EB�C+no��Y�ۓ�<����J���*�l��_P�P$j2&Vr62C�ѱ�m�Ĵ�d�ׯmn�~��Ͼd�Y��I�w���H����ۃ�z	ey
�xYH�5AIM�<\�J�Bi�9����SO2���J���u(���U�fC����4�]V�o��������J\xL��j���o��wg���G���tL%A�X
 ��f�-�]E%wa��lq��9�ҿ[���c�]�� 8���I(5��b}c�4����/;8덧�G�џj �~+�6��?�ߜ�,]8�Ձ������U�MTd��;F �$v/?��&t�z\�2@`q�|�?�g�.����Ϸ�Y���j&�%����yԣ�j����F�Zw��C�������c�-[
+�B�aUE�S�<~j!m¦�Wb���j�уy�K�vΎQB�_2���H�`�|mh�:�^���zA�Զ���f��Q4������|���<Wj�o#���zNm&��	ͭۻ�k�����o�x�=��N�pz:9�9Jh5�=����&H��z\�����X��1��������s�S�rkF�	K4?��c����]ߜ��˝��v\���ޙ7s�\���#
I��SSu/�7V37�f��ǣ	���	�U,|'Y��8kd?W����������+ ��6"�]o:<�]�6E���+류�I�q@h���Y���{(U-�ʤ�ؗ�.��R�C��q�s�e���"�xr��/�<X��.VΞ�6�����|����%�\
Ҿ	� ��O�����Te�X��9��%��x��녔n�i[�)���El��4�����[��u��ae
�SVSX9��<�Ǉ��,��	{n48$��K�T�G.�D{{�k�����k�mG;��F��|��2i�m��r!��N��2����.��?-�a�C�s�,�d9��y���G�r��6ڼ�>:w�:�	`��H�Y����l��#��zxdZn�Ď�y��X�:/��&���%��0��<X����RW����s�yK���L[Q��/�ϛ4�6�-_�4W��蓡B�>�ΰ��۬��O�QI7v��fKh$�be�����ٺp��z�����WA�)�����vH�h'������2�bz8�F�Y\
���wv�j+ʗ��LM��K�<d��l	�j��ى��C���&�W52�"�J"B�'�*-(��tR�����р�L���5�"�~�'UjZ��j1|9o��dT�T� F���P��`���.��e^O��Lk���w^;�>�*�=�b�����+Qn�N����Z����&#_��oV/��۩���νKZWrB�A ���w�b��I8{=I2�Bh�MM+��vu���8A�ˉ{�δƓ��!I��풴| e��U�{��Z�£+��@��o��B< ���H���K�s+��R/pn�@�-��cִ��\W:�W�x����=��e�1�g��Y1~���e�$'=~����L|�d�|�~�/����/��̘V[�kmCKe���r}s��_ӥi���+�م�Z2H����v�ϒf���g���b�V��0���H���ݠ�H`R�`9���ۏM�o�z���,U��%G\Jt[�:�Ӧѣ�e5�0�{�Oj����7OJw�u��8}D�X��(?�d&���{���`.ğ>�;��Q}�f3ͣ���&.)��#����+5.�J�A=�o��o&��,V���Uߘ��5*5i�`%��v��z�;Y���C�Nf�D��{�SV9w.u�������ĝ�����f>B���^��c�����!�n���O�*��%8�UO�������S�'��6H�,uO��rG��.]�t*����a�_8����ky��j�琎�
��7�\���/����_*� �o\ҥϊ�s���xr���!U���0��������,�`�.(���A8��H��B��*<����]2v���f�R���t����*�
wqO�F\H_��I��R�;W&�g�	Cq�,|���U&�f�=�"�݁��W13(�����=����!*�z�h�I����Cac�Ϋ�m�C��3	�Y{��@]���u���������LWZ���p��Yc��;��|@l����*�/�*VC�v��[��)Z�`�ӝ]��y���׏�ofl��e5��d)����PJ2���󰜙0���Y�Mݳ0��YQ���㟀�^b���|j888X�ZJ��&s���x�P��b!f&w��a�`��	v���}��](�q��<Sx��t�-��
��*�QU˲�]��ˊ����W@��dq�]ۇ�������N��T��ap����4a{$#��ʵ��#�XP�<$���#\@�8�-o=eT
���Ĳ�C��FNx+�+֓}�)&�M��/���8�ш+�X�����!$j�=��{�G^�_ NN�~{5���R| Zvg��	��Q�3�h.X=Lf���ߌ����lQ�=��O��ٚ�/o=���ӳY��,	�g���s���3�M;S3�*�9bS�i�>�OH����3S�Q��R%�vdw�1PX�.����oD�D���a�,�g��l��U��IF����5 ��}N�!�R�V��Չ%��c�$Se���Xy��i�}B颋m.��� d�2U�m���#�)s%�}���ˏ�O=�u~�z����=�81�$�1F�P̳267�3Se��1�,����0��'����䖅����D|�(�l�?�f6�1�����>(p�.����1E$G�<A���p$���t�����w���QNr�nAY��s�I�Q�)A���������F��i��q�H�\+�wi%9n�'qU��%_:�d鍋;W�c�?�q�5Y����k���c	۷����t5ޜ�s ����H��bH���Ÿ�.���Ƈ2�x=��zV$!�{C�r�y�� \��<��{c�_dT���	°�ժ;�py��顺��.)��םO��b̊�V�Yn�Z��0Wre#b$N�k6-�+3��?��%�*��d�!8UH]�w���z�ґ�Q�L�a��$�T�A}����E�\ �Xx����?C؁����bM@:�}����͚<�/����`d,W��(��^:�s�	i�V7�1e�\�c�l��G�
�˰𓾰&��{Ҁ�q����^�48}:���j�=���X���3�ڴ޳����:l[���w�o-]�����i�-T7f�{�t��~�M@g�L���ä������+���(�u�fվ��2[^օ���{d�Y"�0����I����!(��P���|�IҠ	���R���o�~�Q��,�4~a�c5
R$�;�{������Mռ�u�����Z5G�xE�������a�/�?W�UIy�#����@]Vb�����B�OK� �/�����6�ɺ��<x�d�@ �Q��k
�Nv.��6�Ȇ�r��t�۽؆��u�*6�YU�_fk��������C����Q+����6�ɾH��6=��Ǿ���'3rvWk��x��O�.���{,��{�G%��C{.���VF����{� :��_ʨ�J�#oPo0���[��HY\��i|(d��+��8��D'�PKk�Gٍ�jl0����2�ڱ���a�C��Z�km���&�}Z�?��v2�>���߼
~��5��g�;�#P��M	+�1���9��z$?"����΃�M��/��4�{�*.�Ѐ�����>�S���W��I�wy�r���y�^�M�K2 �NP�q��!�Th��͟X);��ʗ�H�`�<ᐾ�[�i��'f^�#�R}z�(���/kE��)7��$��ׅ<��[)�
�֍CJ֖��'��5�3�j�lPs��K��V��aO���l��YO�|��O|r�5Ua; �H�-z�a&�W�sH1�	+�#&~A)�m+�vD�%�U}��z�mN�u)�z}�l��
K=o��_�_�?�OX|��ǋ�`��ir��$�c�]���_����k#��h'���	�eS�e���nB���4�&#1Vۍ˶��I��p��ں4GIC�kc���C��c��8'��b���`k���������F���.!��N�vM�r��v�\>�Ą�7��M���w�Y�f��v}��Sb�'V���͒xp�!�2xUU����a�~V����gxX�.5�S�?����r�5~)��֪%�]{�+鼘�7Ӽ?�Z����G)iTOb������������(.Y��ŋ���P��dڬ�n��{-�	cݜ3��Z��3�:r��S��G��2#W��
��jk9nF�Qc9��lR�]�����[{Ψ�z�?���]4|p2��`EMbI5�B�+7u��fɝWР&'iֳ�7���bl�����<L�E\#h^=��B�����_��;���^Y�)`��6d����֕^����r-*�j�)��p����ϔfH}=uH-����2Ϲ�$&�Y�x}��\j�F�c?ơw�qP��nq��/���P�fs]��.����ݞ�q῁Qӿ�;'�&t���o��y���6���|��X�p�1C�އ�K���9mK�����P=���}_/�� �u(�8/ƼmNV���t�D��d�ed2M�k�0���O�N�)�ք� �ɫ�k���Q���M���js	�vU��7��b��4Ԟ���#
�Gt�B]��o�0OOx���M{_�3tw_��w�`�>v��/w�it���J�N?�2���	�Zi|�:FR�����7`Z`��?���*�Zn��F��~a����{8�X����=]��#zh>�����Ԋ���b�Yj�#�����g
.�RQkB?.����|���]p�g<�����֓�׬_	T������2b!C�E���x	�^�U��/���m�j22gՕE�����]�B?�B%��J�$�j�����,�`���}�4����<ӎ�Z���&O�k*TՈI�] ��Ӟֵ�/XA�=�[�`VN��f�"<���S���ه��b�w��`2��.�X�7�Rm�V͑�Qn����V��x�G�������o����z���|��I�?�(�ܙ��¯t��OΟ/h�ǻmZ�.���j���?���*�%�ʟ�4L�.#���RVE�s)77Y�s9����? �io���X��%�-���x;q�p�ˣA�ҋ��v)?
)᧻����Z6V0��\��;k�( �x* ;NvT��_?=��^3�xЋ�*
 (��(��m0��V�1���)�G�;�Տ<���t��'�m�����a]�|�hq^�N�	8%���Q��Ur�SF�=J1�p���H�0��m���o[5sg[�0������_���^�뽿�_RV��u��	?D��U\���_i���N�0�v3�o� ��~�ɼ�
AR�;�]�n��?���
S�N�\�
�vt.P���+K��?�_�xnb��,ȹ���b�;y��f�����Uǀ7��.���(����HQ����ôh#>b��u]L��a�/��fx��"��L��<��i�!N�e���X��2>� ��V:��3v��QB<���������A��z����!!o�X�\��_hPIE��Ѐ0��}��Gf^}��%��~�W}D�v��t����#vy�Rh�?_e�*�Uv�8Πƞⵝ&1S�6��D���n�$��F2�׳�Gقz:q9��k�3�:�}9Φ��>fmL�M@�V8̏_*U���?�;�nK^��y�-֤�-�:	h>,�w�K�Z ���}iwǡ4Q
u�K���%�"j&��t��O
�6�����v=�8���]\S�HŔ��[xzڂ��[ג�H�$?�Hz+��$����÷�}yt���WC����ؾf�^E�+��Ÿ�j��d���i�]�I/j:>�H�����3�B�a?���ۇ/z�k�:M����N}'���6�<�M{�H���x���.;B/�r"��l������O�c�/�H5OqzJ;�|�bSN��#��0ʺ����z}3�6Y��y���\��:�L�Ld�O__j\W����"WWwwrt�"��3�B�����_V���bV�Rb�Ѽ����)����az,[]`���s�}��$>~E�R�=��=3�޴���/~V��e�g�F>��]��'�MM���Y�|����^ѧ�Yeoʸ:iA}l�OO���~�uB�9_�ڊ
�r����I����ݐ�<��'�w�n��?���=�}�U���EH�%^�D�4-L��NS�%�Dg�T~��6���b��rl�ê1]����R�5/G�#�O���B��vy/��K���ϓ�|+���S65m�!�37�S���S�,�3z�
4p�Q�]��!�o���1��-n�IW)�g��'�|���'������{<��W�U'���K�1���k���kc By���� ���KW��ge[ճW����=�WQ�e�M����Ǽ'�Q��S�����mUe���@�+��ѭл俆�㲲�߸qC�g�q�h��o�ݏ�%��Q}.�T{�
�6�R��|�yk#1#����c�W����.f���Qr~�����}w;�n��\$���=�*��`�2���C�-��x�:)OjiTd�"�>,�}�_H�����p��|�������~V8o�6�^�u��ߵ9�~�
m�=�Xn�Pm��q2xp��h�霺�t�-��}_�}<;"�W��$�bl�q��-�E�dcs�rb`\�󮔺����8���^B�f�.�Ul�,�>�����{���\�ԛ���U�%=Î�`w�zGH��=����8\�2�?cgz�Nã�tx���_i(��ݩ��g�S�� �τ�+�;���P�	n]�ҧ_��6N�9a)!�mu���k��{ɾQK���ڗȑ��DP���#��I�^��b���T�{�Q��[ʥΟK�d��	�h�?���5T{,L	�N�GG~�brS�\��w�xyҼ�_�����F�u��4~�	W�A>�����R)�_ZM|Y���x��D��4��C���N�>�S�ӛ���.���wo'�<[��|֥]��ǁ���<M=�[)�ܙ��.4`L|�N���U��-�Z�Bҹ:{�TGa|�e��������vά�])�:]r�p��3.3�3u=>� ��{_,0����&fͻ˞��&%�/�����!��������D��o��a���)���q���j4����	���l�u�$fZ�_�+���eRW�|�������0�����sc	��Gb&g�q��3�t�򛿼�Wi�7�E�b��$��;���r�U�b��{�*Skrپ\�m��i�u�.'>�0�b	����',>�0�E6�|W���6�P��#�[�%4�O����yX�����2>k�D�<�����uўs�
?�.��-�����t>x�h��rҴ��a�f�)HY�o���;�
ϑx"U�^Ys�H�;�-����C�<Ðk�B\VKF�Ya�]j�u��t+��H1|��i�<v$�]4��S��U�P�9WH�?sn������5�_����bO��~�n�r��jF?�_p�`ۈ0i,w���`[%�����������r�vڤ��y7F.�Ky�N?��c;�^��D����<�� �k�t��}gZ|
���vv�8����߅"���N�_�^��b4j.42��c7h��CL5��K;�ɣ8�w?�u;btK}*��O)\цBu�c��cz�o*N\�ku�������3��F4�?)���ԇM�f�D��O润��')>ʴ�x{5���뫍W�4��nL?�tq��#�6�i�xy���49�}pP��^�+f?]#u\���s��a�1R��'����x�~ay",�e��g̶�'���;[�S��{Mo�ɀ�df'���C�\ӆ}J7�����Ơ){��[߲l)4�s��'��)��UA��ύ@��JAb
����b�
2�ѓ����q�:oi^��y%���q�V���3�Xv�n�^��_��-�1�!���͸��^�P���e��V����n)(�r��w�k]|t�mdP��>/X74B[;ܾ���	@� z�z.Df�}݁Q���n��IA�Lg;�����0܀�9�w�W�X��%#jv������C�aS\�f�������hi(ɯ�Q�5��6$)4�|~��su}r����Z���<r������י-g��F��_B;v20�ߚlK��E
>.�wS��?}�,� :0Z�}4�� �\��)>�o������q�㤥U���<�fX��¨�K��[r��S꘥�ƶ+-��1:�s}����h�(>����1��P'��wa�s�����q-�JӍ��uy�t8���$HX��x�P�o�7�k�U*��t)5�o=�#���Uǘ{������^dOB`n�����3\�� �ڶ�uZ�v������9���c���w��Mn�
�J͸����]܆
��^��7��L���]�f���n���C�[��
���!K�����C�y�|]|�������ѩ�z�5�.�ů5]̆w�)��[�xa��&i�[=����vW��[�ǔ)�{�LX�������\��M{�_�=�sx����F����5��!��]�ݤ�>S~�K^��u3r69��5ɫ6�E=����mv�[r��V+#1_#7�����J�1�,�UFD�ȳ8�ͨgs���=&&�}|�9�w;�Ь�ƽ�A��hR�K-�n���E����,���Em��e͘O�>P����{�Ze��?���q�<���(���f�q0�KV��Q2�����]1'3��K24������$�*6�c"V��\�SέkG�-wwhQӒ�����xX4�,��V���Ӎ��Am^��D���_yVj����}��O[,��1%�@q��Ɩ�Aa��Q_�����y�;~�_,
/�(8�|@`7L��PW��@��;&w��^t#���,��<(��h(G?4y
�7����Lb�I��S�7��(�_+Z���F�0\�ch���z�xc�=���k�$���k�����&�A�CB���A������S	��;�����Y�ߢ���;���0�����\׉*�ݒ��ް⛹6gv���5D�bO�!OҜB�߯�ԐT�B�\߽�l�ȢW�[�Q8���Zk].�p� ���\"�G|Q>~��s���C���Ć.�tD��;����.t����\|������d%N2��4����WxG��]�7B�_���4~���ax���!��BZF�}U#����wϊ7ڊ��s��wM��[NԵ(ԤiT_��4�$���Cr;����b�W�������B���?m�/�{��'Pܕ6��~e�H��{�۟_��L�Gpۂ�Z[��z�YD µz�hT㲷]���b�v�Ma�T�M�9���C��C�@��c��J�KY��yH��x��-�h�\����˒��m�8�r&����~�ގ�j�G�*�d�qB��'^޺�M�X�y�f�Jg���-y�l��5��_���UxU��9M<�	�f��c�4���I�V�!V����`��"�B>ka�-������%LȬ�h�S`b51ӥ�y�7;�FZ\�
�#.�S��Q2�� Y�k�>���@�E�����__���}.���Z��{+�:��
!W���͙�(�r�Z�0�^J�����/\[P��h�lR?M�
ZB䑬9��8Y�ۚ��w}��E>�3����x�8�81��wQnn�i䷱u�����z޵�3�Bp�Z\��e�RP�0�tw���8�y�t���K����7 G����x����)�p��B�q� g�;������������Rg��7�w*�]��!���?��E	_��t���j|R���	��q^�6o��SΘm�5��r�(<M`�o�s�r�!�9&6��N����+�{Ƃ��K��N��Y��5�CfL��Θ�G������b��&��]������qO6��GƧ����e���U�ϕX\��>R���p�NW$M��T������>���ړ��L��@؅�d$���Δ�Ҥ:W\Y�4��m�v�|`�[�l�is��)��*�^�����+x���%<%g��{����D	v����Y��5!���Vk|>��c�?�q�J�I�q쩕�㶉%���������^�*a5h֨}u��)k�yc����0kv������ <�$-8�~��پ�9ލ@or�8�fCH*�l�]������`���1+L�xk��M��u�o����.����?���8��w��m��*.�k��	��[*�*R�������v���bv�Lm\�v�	��熥����wϖ�ֽ�gZ-�M&x��*�̹�9m�e�.Q��$��l4�Up<v�f�4ġ�"_F���-�)v֑2�C���/,��0�������zRy�ɩh�6'\5�U�V����IV��!��@�����l����Y$+��`�ݪ���{�(M��Ϙw�wk��ri
��~��K�����\���T�����v�cf����e`��D�\�5�I��z�������8�{�co,E]�<��o����S�X��]_%�_���$����D��f���̂�L�` ��?��з�����S\�d��n���ߛ� Y����*6h@/�{m�-!J��~�
5l����g�m��ւ�c�7��[|&���ה�isC^I���f���}�#�hHVr�1w��zgf�(Y����5uUf����K���q�K����u7n"�V��}y�y�}!�'��������4��p-wخq7ܬ�S��&އ]�UP�~
I���x�jC3�z'��y"9&�Lb��e�V]�]�

���$(l]Pm�ē*t����sw�ur���(+W���M��*|.KMQL�@H�ztw7R��j���mӹ��Uƹ+�K�|t
@��t ;��,'� �n��2ŬKZ�kL�=��th�L��\嶕tt������%[�������VnR,�'�q�)�̟���u(���b�/�����sr�U_K�(��~3*1�z�v��l��c�s����o�|6)�~a<�Z�F¤������0����Q��3����鷙ߪ�1�(���A~��B>�"�~2�[.onU���;~\ƭ���u�Ga��l)d8��ψ�I�Pۖt���\�3;����r���vb8m�7*����Bzi�>�4�Ĺ	�65����hZ�AZ�ڑ�#����ר��n�KJQ���/ú�1O�'F���!������ �781,��.y���F��:S�"(����8>�����''��-��3��Jv"	�k�ר�֗6�.Y�7�>/E�N�Cg�&��9)M�h����L��[e5���q����?�F! �<�g��c⡸c;>Nd|�:R��x��"�+Y
�	kƬ!�����k��n�޵����-�?�;�@�ԭ��k3�x�ѻ>��u����b"Ԩ?��q�3H:rݷ�upq��È�����x���u�`{��`���q�:���he��+�Ն�,u��c5�,��US*�Ō�=�r�0��L���љ�N�֮��/�o�"����� ^f�]�q�-f�tl���5�� CM��M�NET�Q��T|#c���@FN�|4�O7��QDDDp��gL���=��gޛ�I�ȵ"7a������%aI��2��O6���gغ����a;�U�9���Q̏If̋��|���n#�}�Fϰ�%W]��m,U\���׿�������mV@O[��é���g�����D��D�wEBӿ�/�`��A�G������K8PgS�(�}��)��..�Ws�^������[��s*��q.[�����	����ݮ�b�cB��Ҋ	�>6����]ە$���N�[�Ǽqm4�#0�S��Y�ed�44�rhY���*�"2;���	�Ф������Cea�}�aRO��a�0�F��:X?�s��R�?i^�9�����@
,{$�z������S��rDiހ(�D���50w����N%�hE2@g��2Эwa�!�n�wΟ/	eu�ܹ��_��O�+�cBvU���/��1ש�_�;�� ��<d���/����g�V���Xr���&���У�������M	�6D���.��ll0��C{�?竭b҅���G��-7:�4�?u����S�ɷ����HQ� ʄx�|Z&u$EY�TN}ϰ�CRB��]̬�ٵ|�&lw�vK�S�6�k�zʁ�r��1vG��eҘ!T��ӑ�ɞ3����Q=��!B�nZ��vZ~bL�ro�q�v]]]$����3���M^%��{X��v�������)���k���}/��z�G�Z�4fu�p���72�]��/ ��'�Xu#3�P�)/q7�6�"k*E5��/p���Gb���9�y'~IE}���:X���ڨ����;��X�W��f�p�ՙ{~rZIӷU�j��)�J51�;mo\o��R2�Y�{�xR�V�����d�YWiQ��vZ���F�]頃�UB)��ue�m���!ϚC!X9Z��3c�y�?;�r��;4���o�gN��ܔ2�T��?63���-uBu�����*��mG�����r���
��e6��)ϑٴ����ǂ�F����|���]8��%`K�%��ђ[�O�V���^'���8���w �J��Ȧ��3*��@�S������RD���� �˒6+u�����T@�%2�YC4\M��񢢖IJ��C��\��e5a��,q��]�{f������&=�����*\�/�1y������Nx�sVjZ�:2a"����A��ba���|����� � ��UQYp����r�������S���[�.2b1��;e�M��{q��z=ߟ�a�l��*��^^���׶Kx9Ԉ���W����$�������������KҶ���M+�����.��p:�&\o��e�?�����|1�?���A�|��(�ZP[��P#hځ�c_���ٌ���ռ��a+���ֲ�?��!<ɋU����D����Ђ��p˛����kt�a�ㆵʤ��R�,��H�	��Z��8����g)�)���JOx�P���n1��ف&�$)Vof6��+�A܎�?��|�P�2���ԋ+�n�Kˊ�^��/�_�j�}�S!'P!�Xϟp)�tw�Q��Cx�S�d�j$��i���㝺�h��N��� �Y������ۏ�m,�a.=��N<�XЌ0�54�}����{�L6�І�Q�^_M�\Z׿$|��;}��N�0C��,^͋�k�C zgW���5�)�j���fl-$Z3y�(tFT��k���!�h�2&{�9-2�����1'C�CE��u�|��gE��x2	"�J)���u��Ξ��;C�Y��{'|l={�,�������%7�Q�c#˽F�9cw���kɅR��/��!Rsoǹ�/�&ٳ��!\��X�#��f,z�s���/�Y���6�5u/:�[4�,�����E��-�.��d��e�J[�ߓ��܂^b��O������:y:���O�OgU�#���f���4��"�݂�|�|�7Vi���w.`6!߫�rl�m��賬�{�bI��"sB�y�hȆ$�?�����"(�޼TBA]`�X��/���,b�	=�:iq5���c��hږ I���y^� ��)�}�^���?���L^��zv0�z�DN�<{9vv��Y���u�aP�ƀ���tdѝ�1��ތ5�(\��?�h�C3g�sM�$��C?a���
��|��hG����{߿
���������w�w�fo7�<�U��d=~�r�V6�i�� �V�c�j�^#�#�C�
�ʑeJ2�r&����n���1�'`��z,]��A�a���5ݜs^U-|_�G��b�p��y)��l�4�&�B2�iQ����9}!pS���O��=�Q���Xn�D��,��o�z�[�]TRs>����z��/U�����+ދ�>�������ן�8�ޙIƸPK,�3P�#�1�m�i��=?�H���"�lXC�O��R�x��8�����v�_���<���:<I-��2J��^e�(�O:a��;$8�:�p�:h�+��<o�C:f�,���:W��;a�t]I#���A��{C�/��й\mnY"��0w[: ?�s}�9�,����.J/	����%����ӵ0\��WN״��ǿ�^q�6;D��Y���/�9����>q�R�����y�UJl9[���R�B�L��X�~%o�Pgi�t���;{Є	�O%nud�ʲdn��6iC'�c/��n��g�&^}_������8�/&���(X�����2�H�Ȼ\�O)����y�1y�|���C"��eq�L�5S�������.�����?yx�Qq���h��d�Ui6p]N�mQd��o_1z����+�vYJ�0�u�[�i����6<)���G�2v���� ��`2O�ڃ���bÎW� �F�y��&�t��DP��c��Q~2�rDkb�͞^gy�Г4Ѝ�*���'�[�"�����G�����@=���܌��D��6uT�����z�v��W�>��_�$���IY�_�~�P���>`�u�p\����&�v����%ܶÇw .�|̃9�~�cBw��U6|�,�a��ئXWx�f���(��>݄�gOl�c�wO����ݮ�&QaEY�l�!��k��?[u+O�A����Vv���%C��Y���'���1AA���^$%{�W`���sR� 6���hpm���H�m:����j�-�j��?���dz�;�#��|�j��ZAp�!�FB���z��3�
�
ae��fUb�z9�b������S�cd!ۛ`���<�v��=��g�#�.�n�f[�OΙ7u�G�f�.��#x��=��������&�*�+ⴠa�opa�,Kp�E��m��ߴr<��8r r�SY�\��tn�����7��v�@���~�_�4�����֊<���3̒��WPN��'1c4
1��TҎP�Vf�]��o�'-;�gw�p�с��|��_�nY�}0~hRme����ѴHڢ�4� �ǭ0~{H��/�|1a�X/��(��T�I�s � �
1?�k=04i@����]~ƚ�n�,y۾/t�V�f6�.<��_a������-�z2��5���SI�Zx�z���L%�0Zx��%��F<���;��9���� ĩq��J=P:K�$�|V�b��z�6v}%�ni���X '�~Bp�.��'{��e.ᡝ��{|���e��e)3�x��SY����HWb�u^*��|mJ/��ǣ빅�53T��cc"�Y�RQ�!�0��t�!�-��<b�"�]0��_.�9��^�֯'��$c�^�u$��)l?�IN�5�?��.M�S-��ȣ7��Y�H(��9�01���M��:	�c�����%��Ҙ�h������a=� �[��߽l}%f�(kF�q��P�hq��f{. �M��d��"|- �/�k���-Ccq����(h���W�A����`(Pvu-B�a�k�Hxۻx 	_��+<2B��ٿХ���"G,������>��n�k�ׄ�*�ί�0���U�0�dwz�BH�?�-j#��rr���/�C���}�&{�㵡c;hB�	��tȣ���0a���\f�L�܎�Ƈf�A:�=;=3�������>�4�9�.fgl"�f�x��賛o�ۙ�F�~��-J��F�>�6	���T�����B�4n<$�_=+YF��\GxN�L����pUPЁ����p�����>~�8|�j�,L���~�^aS4YƆ�����'�֡�Dg��3�WHX�^����Y3�[n��1�"n#+�Z��׎��H�(��d�dYfb��2	��&��u���Ls�i��1)Vzd�2�s��d��/�>͸ل���r�0��z�������������F�9�5P�~ʟ%&��{р�{�Ӣ�˥}��~�4�u�8tI�U$����~�m+�-�� òh�/�<.1)���JT���L�P��|gRAv����m���"�m:x.l�B$b4:��t��x^�K�	q��]>�Z颎�/w�g����̩U)���Ƨ#�U�17R��Loj��/mz��YG�������\/�N.����ӻ۝����K������zOd������￉�%�M}�Q�p�O/�k�����A��u�6o�g����~T�a�N�VI�b��"�Od;�Ϯ� �w�A�G��d�����/��ߠ�F2IA{��V�2�n���jtzU�{8*�2������iK�%J}���{2�{g�#�@u܋�/�'���)s���d-����.����V�д�����ZM�9!<:P��t�>=�w'����A��P�� �D����R���d�k�
��31�ܸ7�"c�/�G��TbĬ*m^�R�}y^��LL��f�'K�И�94�P��"�\��j�O�_�>��a��tbJƄ� ��Ij7�t��@�ko;�pZ٢�6�*56$�����*�U5�|�O�o���5��m\���<��s�5��n�?2�Ni����EG��h}�|�����3�)A�/Q���Ң>���6 �l�tx�1$�}������c��IsL&H�A�"Hj��5�7&��o7J;.��;q���M�2ǧ��{�USB��'�O�)� �L�Љs�ۓ7�I�����d=�.�d�����5�c����ِc��c�7�8�Kē8�\}�����s�ګdA5`���8�c?���>�cxJ�s�6��e"�_�$��ޕ����Q�Z
8u��Z�'-��J�#z{%S*�0����M���ӕ�/�6�4wuf�툦s@)I��/�{�	�)�z2�S�j�^��d��\~��A: ��$ʺ��׹��tX���l ~�]��\�}F� �ǚt��6�;�V�xED��8%��g(�Y�Puul�S�������&8�ݜm�2�0�N�vm"�V,���r�L��u��]�Ѿ�&�\�ox�O���Vj_�|k����$	'E[�$���@<�E� ��8���H6ϕBl==���O ���I+[�LAG���s�=��;��R�	p�f\���_�k4a����bu����M��6}~M<Zo��T *L����ex���gT|<+&�v���-��(��0n���$����W��"%�'1~I��bB�ܑ��/Jb�N/h�ܭ��˿�uzˊ�uS�!0qh�i&f�"N��=��5H��K��6a��B��=����u�I�͐!��X8N�p�ȳy���!ȋ�Ȅ �
)44�&?�c���z����+�7��.�y�c�x�� ��j�����H���5vu�t��0\��\�5�_p�,4U�l�P��t
���(Y�1��{��C�S�Ab�G��5{���͑�1�r���$�'Lں$�b��s�v�a���H{y��/7R3�k���ٸ���>R,a�M�8#un�D�Ӳ)ta�-, 9�:0�����U\ܧ�:��C%���M?�$M\?i����u�˛�{wD܇-���C����giX������v�Mޑ�GC�����2%�W��m�G��XnaGiޚI&�b��2^vE&�P�r�dn�A��":�u�gJ�f���q	���q��.~��fQ���ĲTZ�r��e.Ј�LB�e��Tv�C���7��ں0���|=��s���.�.$E��T��z��vӕ~�����q�=��A��v1E��[�g��\�&�̐6	F�_���Y�Bs4{/"|�x+5��R��*�!B�4�Q��l1aP�s�>@<�����^S�gS˔�TH�cD,�'�ٙ��^��ۿ�r/;�?v%	�a��Ļ��t_�z�^�E�%����+��\��'�
1�JN�R�����Ј���o���yqWG�&� �ԥL��)7[�g���P9�k���'�ع]��6R��H؀:\VD��s�` �[D+�+ށxc_:.^�jAPƅ��$��*h܁,{� Us�W�u�-�V�~�!q����G�N��{�9	h���u�ϕW*��YHrH�m�PU�I2�}���^6��m�9��T/!����o��=�0���bb7C�����j�� u��lO�3\!��M� O3uu\g����d _��O�P
��40���&���9B�P ��w����㦃���R�|{�^Ts�qb�CF�B%z�_h��1R6�O������OH��3g���1]WPx�n�JLsH����Bs��[��/~��X ]�L��<� �0^��vk����[�3��(���R��E��}^VCYi����c����N��I�(���`߬'eX�FB������m�sm��*��ݟ+�Cʃ��uSG����S��q���_�L{�����ڸ�["�ڤg�=½=��~�Ed���J�/i�ArT�_�Z34Dθ��:e��8w,ͬj�AN��p�_.�Q�㊾6q�,s9����}�>�
KOW��v C��*Ѫ�Z1"p�KK����Xz|v�����A(qݒ���T����o" ,����r�;���$$R�T��4� o��IxD�u�2�Um��ԗX+���������fP(S�)�e=�:�P�sqK��K��vO\*���#�k>�(�X X�h�?=|��O���\<��ת8����М��.�D��fV=CS����e[��e�ӡ�	���j���b��y��[�MD2V�^�����yS��-�R�V�oS�jD$���R������q�s��	�ԉ���:0.��b�\�OK�9�Z��ؖ��'�F�R���N4}�RtS�d�.tiGS����~��v�Jf��=s;��!Y/o[�����=�l���n�C7�W#V���U��Rn�l�W�+e���(1���2�ٕw9��"���V�V%1��!ʯԚ�k�A:�%j�g��J3w�@����a�5��ް1�2/�1���g�ʹ�.�KLKl�drKg1�`詸TL�D5�M��᫺��&D�&�m�g���뜀(���L�4QJ:;!���|�F��6k�d���IF閂H �'R�p��;�#ƪD�����6#7Z67��l68�y�\��F��Y[�~W��l�)<�V�9c��3}IL�w��R��� b^"pfs���Ȳ(�j~7��XѠ7OkRydP��F-����g��Z�	��<�K+_��s��av��3'6��X-���c&�ٺ�o����ς���������'��y�\�@h5��Gp.>����lO-W諴~	A.TMWπ9M��Q�yU
�%������N�+S�g�	��$s=FH@~���(+P5���8��|U���?�_*�0n�����8$�����-@��$��@S�����}�e��ˠD;ٴ턄-{�����1��M��GtK �U��%����h�
I�M�u�\d'���3Z*`C�܁T�j�%�&��܇��Yf���;�9.$oE����gR<-�}���b���W �c*(�rE�zH�r7�팍�"y�`��,���%/���I��:zv���r���?$2�6c���h�w��=
���~|'�'P�9<��]�.�O�}7�|}����̄�v"���Y�LO�J��i�����b��lL��۰�NH/�MH�GW�>�{#�G�| �;V��.��BqA��Ͳ.\��B�%9�����*f4�8�8�!3�V���p�ӧ��HHrkI�2������҂�NCۛ_w��xW6�$�3$v�ǩ��֤�bq�%!1ŽWw���Sc��� ��n�G�#veDl�縋��P��2�/ӝ*���EQ���TH *Q���C��
�XL���@QI35)�q��,���,v���C�:����Ͽ��܃��`����8p�+�tsm�f��b֦j�D�&lS��'K��MU�ޅ�rUWk�5m&��4��-9즾�oι�H�Lzh߮�E���K���CPVu�z�JG��F4�a����,q�����'�צX=�d�?�OvCY������8ֳ�6��e�~�n��A�����M���>��v���啊��SHy�Z�̈���C��!�g�KT�<%����(��I1Զ�o����˸!�4D�f�):0�(�b�*��W(C��9��f[5��J1�p�Q��Ыk���JZ��]�g2ޚF=�<���ް��4���Eڈ��'��7{��w�D�O~���x�M[��0�囩`�>�+��"�c>W�2�v�c�k��3�J��Y�� D���Q��  �ާĦ}��\��m6�`Ӽ�V^� �1�D�g�ȳȦ��+<x�(���N���W�gKR,0�d�멏���r�mP����q��.C�z�hX{3Q!R�Ik�-�<��`��Ξ�>W��5ڤ�:��˥+��U:���pħGj&;$�#^���I��^+Nr'�����Bu������o"X[x�h�iu�8̒b�eBu.�^I�k���?[h����J0�o:��h�:D;@�S �k�9�Ci5U^�D�ӻ����R�qɆ����ܽ7��\[��a��E�^<�Rj�.�u7pٌYV���mL?�z���aw�{J%Y��_��;?f�����@˧�+���uF1O����|�g!:-X���2ESr~a����.s1Ze�k�ͬuC�^�&l���+�^���Z�X]�<���D`�X^��ћbw��{�$s��9 M�xAD��~��(���)�QJ����o�
�Ǹ0����>d�E�W8�7M��#��2idq18�)�k��(��x������V: �0 4tC\�
e9R'�{I2X��"��𑠗.���"
1�a%���Lt�/P8���p�w��@N���n(ԍ��5�ڞ0�z���3	�$D�����4���Q��҃��o���w3kC�Ó����6S����jJF/�A�ɞF��=\K�Gn�G�"%�W^Gb���]<�W ���lP��F�zs��bi��e8V~��Jt��y(����p��l�t��+���Ѷ�_�k�IS&O�� �uȦ�I{��2�Nj��LS��+���W�q�\G�J��I��99�6�{�C79��&|����������/Q�9ċԂ�!Z)m�/K�xe�8Q�%��%ҺĹ�!Wx�ʴ�
8��J�=���%���h(K(��2,J�Z������\K��4���_},u/VV��!	�G�ͬ�����8] ��f�e(��P76d�Z' R[PҪ�D�X�J'�KA�\w*���+�\�@�l�\�SϻZ�/�8b;���Y���?�����,��(�R*K�6\�79�m�Glv$i!�����5�bȿ�(��GKD�{�UQ>�1Gl����<�z�"k'����i����p%NP���j���dL�RG���[�(�oXֳ�����`�6�>��V�l*m����D��J7��2�ye
X6:L	��J;=-�b��E�'����}�t�/M F����2��z�8'�Y1w5+�\����F�|G�N�"ҩB��f*�o ��P?�/�,;y@����Vڡx�V�.�]�ZY�G���^�#P�F�pL�$oI�;Mq� eɚ>6�s�跞���B?D����@\	����P��V�Bօ;&
��8|�T�?.r��o�j�m���4N�&��R��νHO� �
7��*X�lN=�
<���'�z�
�^��$w��Sˋ��D]ڼ��P��?�,Gm�;�0��-� ;��(<Ѩ�aL�J[���^��᫳*"z'�9am�.<i��l�o&x�;s@��{X-�6G,h�}w���d���Y�O�(D��fd��v-��1����!'}�P�ۂ�2W���s4�C+"PB��Y_�`i_"}Tv5I�@<���=J%��b^F`�R��dQr�Ĭ�U��^�5�r��]IW�S���v�I��{�� &��8����v�*cD��00� T(��X>@a3�v4#���KU�<��/u�����i4��"�3&��Dm���[i�g�ތ��G��3��i0
��7L�)�М���y�!��\��Z]i��b�����v׎��ܶ���C}X�:�^N�&3�@��uawyƅ�M�*��(w�]2��YTP$+��cΖ������\������]���	V@9t���eĿ���I%�RD!���>҃����?���V��>T���vT�R����0t���#��aj��X-b��8C��X�<W�}�n� A>+�Ysj��m�Uz��$ҡa�a����l��vh`з�����X�K���u�W6
&���y���M1x�.
�� (iQh8����D%i�lxi�L�n��6qy�n��^o�<�a�qA%	�
`�e~�����:�BN�K�NP4�����^�>�EӾR�ajL�s�����S4q�Bs�&�~�g��^�<�K�T���s�/�r�����aQ��0��3M�Y�^�e;��F��v[�^���Ox���q�s�l�}�4W�/�>0�p�d����2�@r���vO(4�
�|%�mdm\�;���Ck&�z��K�55�w��]�5�AP��`���7 ަ��E.�)y%Z����Q�Ʉ]oH�h%�D<3ŉU3��<O:��C�h���3�.aJw��z�s�����<٣DpLQ}���B�k٨���+W��������y�.� �q���<)�a+�y�dC�S#V�l8� �i��To9:N	l_���_�����4S� Q������1f��ex��%ۭ	��{�IXN/��1�q�"U�E�e��˚yc"�uZJ9'h��a���x3��۔�aG�L� ��ױբ�1�[Է;D���;*C��2�WUk-fM�#U��'��:H��w:�5��29���z�%�(����dSݦ��%�%z��n��� ���6�n�dufL�	�X�?gl�O��V3E?[������4/3��:<0,�l�ʞ�/�@�NP�I�-ul�L^��=dS�Z1�to"/��)����:G1��	&Yd?��bGA����8!z)
�Ue�8�%�9#��^��Qu���Q)����/~��	A!�DN�W�bk-.�[ΑX���j�&���h�E*Ќ�W��ѦG�ĵd�	���%B�D(�O�����r\�����I��%�K�RF�*�m��b��.,h�i��MJD
4�䎴V'�mp�=<b��wP�Jw����?�l1�ķ����3�?d�9kaT
	յ~P W�ɶ�ȓ d�� It������.I��3y&2"�v2�]g������M9�L��q�!=P��8bK��O.�����d�C^�o�60� ']�P��W�WI3ީҐ�mg ^��J��[�r�3ڽ��kd(��o|�$��}%F[�1��:'��^�$S:���}��@�^Y���������&�x桅��r�T��	mDI�J������nhiw��	���9ίJe�x��ퟺ��p^F6l�b��beS '�щ������?Y,�M�4���j��
00�v5�p1�����R�։�������ҥ���@�s�Tzi6�g��b��+���ήf��;��$-,�c*�޻,�]��v��%����B�h;�c��lp��ݗ t�z�R��k����Ab4Y��I	d_��^ﰱ���F�
�n���	�8������.!��g_I��\�Z���2� ���)Cwō�*\G�.)�ֻ��k���o�GF�D:Y��ը���Ȩ�BNm��Qye���)ۯ��U�P�%қ���u���-a�,�2J.�1�:��p�m�K萲�x��F\?|��L���j"����"��6Ľ7���皎��_��}[��t��M<ν$u�����ZnrHY�/=F�k"b{%QF�&\�y���Ɉt���+�a�^���"�@���כ���vX<�����<�����K;d�@�oY��<i�W((!��$���6��I"l�b�?��g��j1��\F�"��$~�#���O=K�5�ѽ%kV�iޟ��Y����z�ϫBE�jO|��$���X�S\OM6�^�Ĺ���?����r��4��_���RK�� OO3PB�d� �|m��~��#��#(IP���ܯq�FfB��'�l�cAf��)�_�9�2�Пi���6��YZ�@�g�������+�ӕwj�'�h�7\��;�3��Cv�+)f)��TBP	R���$ϭ2�t�MUV`�#�+	��)�T���/�ȹt.?,h�L�p�Z�A�L�'Dǝ�}c���+��j�*�w�DH�Z{R3�_�Tl��o���ʡ]Y_,�5E�~E,3�2���������n7W�Dw�/�0謾��"t,8B�S;��m�z�ys�M^)�5�E��M�4�/S��^<8a���pE�Z�֭.%�ac�;:�U�
���C�ZYH��Q�Rp�i^��H�1Z����֖.u���C�ˮ_Y�ב��f�+m<[���Ԇ��lk��u��K�$(��Ї�M�		�����Z��d�@2��W�TYt�W
FhxΘ�8�Ui��#����؎շZ���i�-�1D����sZ1ąm&46�g(�WkiWU��hA�N�}��x}��@���cD�����j~�].��vzL�5y�礪 ��Ǘ��H[ۀ�o�pFYG˶ėrn:^�lY&���Oj��?��!N�t�[��N����p��w�������K��]��D>�!��#jX�&���V!w�����\$�Tm���B�U�G��D�|q�k�C�j-J�%-m�W�#�k��~���H�_Q19�-�%Z9.0~�G�YQ��*8ME\��"����Q��b�C�I�q���+�Ͷkt:�ǿ���c	S��� �_���#�'�Y�B���Q<_�.IihƼZ:�i4O�E�-�-�okp��[A�/a���)~X���z�7����^�^{?����V`E2-�ۣ	�C�����,���ղв�#���+��� ����Mf�\��a�o�{�F9[Uir�4�Md�����A��*���\ӱ'FB�2�_�S�z��PF�&�O�������g8�L&��"T<���Ys��9�P$D���ANf���bk�Y��6�l�e�;�Qz+�Q;�4���@��0y��G�\V۠�JK����݉ɻ���Բr�&L{/R}K��b����T�ԕ��"�l���?2�N�>�(�������|�汉M0�D�\<���HF����*������C��'�y?�3�ѴQ�ho�㵁�n"J� ���W�����T��=�꙼��a�}�s��ى�e6���ӕ�$l����Nh&وF�fz����L%&k��6?�sgHg�	9˴��WE0�l����t��/=��A��i��n��y�dB��1i�(�9�����Fq�Z����zӾ���!W���w݆D�3nA�,�
�R�n��^��\k��t�1n2(�r-�����Roqy�R�gO�mk�!�N�Qn��n�ٳe�_�<�
5�T�������=P�'^��(k_�m�l�ƐU�� �
S��i\Yt���K�&�L�:v�/�B�4k��}��a������L��B�R׺�q�B���n�J��џrŠj]ؒ�k�g�r����*��ﶡڶ1��+\�@�����*�V��.A��f(E����f�BB�DA�{i	��f(	�zh�A�繾���̟9��^{����O��wt��И*�wT~���?%)ģ�<��m����o�&s�_p�:w��"���)����Uq�|��'�;����Lm;�ģg}��g�t������(��3�+�P̞����9IX�8���t�![��r���/BK���U̥B�0�!�����/�_�k���l�zVZ����=�Ŗ�NV�I퍊\Nò���H�,�;>{�(�������\�����˜S�?|9���ч���lR��lz|��TWd�'���SF��E��$�N�`��w�X�ٲ��h�ڼ������[G�o�U-���	���p����b&��	��������է��X���@YC86��o9�=rټV{�'%�Е���Gw��'V-ƃO%wU�z�c$�~��?Ir�4��>����<��&�:T� n��&�Y��~h�'m�ѡ�_����8n*7����B�ê����2w�E�J�3?���e6m��Ӈ��f�N�X��ֹ��~�a�p�:��%�<�%]�D2��gb�2���I�(�[�O�o-A�m���=������ܻ�2�2���UR��?��{�I�<b]f�43+|��2�@h	�q˽��uV�!k����2���G�+N�{i�I��s�w8	:T�Z�#���r@q4y�u+���Ƅߵ>�SWu��䌜�n����t�I�;�vX�U+�ǂv�q-�agQ�L9|O�c���_ͱ�t��Q��)����F�-1��U�ڴ<�s�$T^SO1�K���&Fu��&��6��|W�}�P2�D9{V��,�f���߇w�2�2�C*�p׳^w%���,���P sUw�.);���)j�4~�t��T@Xk���Fm��0�b�����S��q�3.�ذ�M䧅�%1���"���eݾ
�T�籇���n��_��ȚR!$h��xD�lZX�	t��7L�oӬ�:�>����U��������@�՚�x�=o����ۀA�f�ӌ��C,FZ�Le��?��["\V'��	��uS�3ȔI�RS����I�ՑO	}����ɑ���³�0����C�r�%C�Ig�-[p�˵��O��)�_����U�uݪ%��
��HT�Y96|g���Ǖl�����XR%���QhA�gL�T�$D�@T�MۍȊ���=DM6�~2���/�X�Y`ʊ��	��!w)΢�[1�u��NU��I/6_�қITY׈�8��ÚT��N�ea�u�ę/�����̀��$�sF���5�)���T6���w���#������z�z<R��#�*J��靸�ǜ�����|;�6��L�_Z�YL��@26̔կw��������S{(s�žT]��{���>�j���d��D�������/�u���p{+�)��w��jn���P�^���V�������<�M����
� ���]bskQ�4Ro����u��Y��A�aj���л�5�]∇�{�FB�+1_��pp�c�c'/,�+�o	&u��^���Yʻ@=��F0<Et��J��YYI��|c��S]K3o�:��	|��֎
���ur��X�9�D0�ԃ�K���-�/q���,-�A�z�6HA
�I ����$8K�� n�n�rleI��}��_,k��U��J"�6�х>��S�a��?�)��B=�J�zVNY��cf��5��v��3�b?��Cc#ļ0HqI��L�Y�vE�N����3���ݗR��uɁ�?j&��Q]T��,^�r���v|%�\�>�о�!z���7�*�%n�gn��|�'�J(�ɛ#2���#k�{i��$p�\�ȅ���X�@�T'����l��O霈��YڰJ)��H�bOBU|��^���d�<S�vZ�K �m�q�A��u�`����C{�s^��H���N".o���b�	���+y>2o!�٦��~C���Hl��K��:;�LU�Y�[��yg�귎�;DsPM�n��D���#/��/��ۍ��=.�����?�)3S�7�3I�����k�j�xP��W�}��i�;�#��{�]�D���+�Y$���6�GWa�z���
+�����z�Ё��߹ߊ�X���_�ˌ�����f��UT҉5;T��f?RmJi�kx��/@d�r��Z�"r�z�)�U�Q�o���M_O�޲�Gk��8�^���q�C��.`oeŗ	�R3A�%'̫��d�IU�����[���ɚ���S�A�9l1*÷�Ҋ8ف�{tf���*���n���q~�:k���

H���4�&i�4�׭�~�5��-�z���.���60�'������w�45B�
�n��C{	 ���������So8��n���e9��������O�5և�ǣ3ر��7�����[��	��K���;�*�q5	�\z�j
�3��R�8��Wh]DzM�����"���8Lc�����@U����^,C:,8���$��N��*)G�j�.�4|v� �N-?�r��5r��l���[M@�E�'{[��ɾ�U�@�G��8����E���G��8���G��YQQ�� ܛB
M�/�d��V
���=d�%?
jYw|AQ�->�R��ƏU����^�Y��g|��Σx܌Zޭ�и�؟+�t@�K������m�Z|�]�
��H)����:�\�B��������v�]\k�����iʆ���-�:.kT��YX�m��*��0g���$M����2�T+��S^�&���w@��L���K9��bV��w_�j�AthH��
��uȨ/?S�S�������Ϭo�ǃsk��(�1�-�X�:�p�4/��9�<?�R�j�AD����`yS,˘}���8:����%��>���(�#�fV��).�������nN�8-D�$܏O��H����+���E4��>"�5���0V�|�r����/ٲֹ��+���a�IE98#Ut]�f�2ܣ,�ʻ��ړ)����5����0�����`*2_�`7C�]m<e���F�µ��}�p� T�y�O�1U��:ݑp?�[�_e���{�շ��M�}m<"�NG�>��I��6\�c��� �
�]r� ��e�����iE�Ʀ�gJUiEnj��R��0?��  ��ef������jK���I��#$������p� ;��X~&@8˜�1#J�fMÀȱ�V�t��	��(g�XY#����7�g�E�9ծֲ�Ψ&�����=�u̲��SNK��Y��Eɸ���R���+��M�c�z�,}�zY�W�Cy->�l�Ya��AK��"O�̦8U���X�>�Qm�%�m�<� �x�?H�]f�3O ��d��hr� Ex�]��*��Ƃr�Q�۹+ �K1�'��&=K&6���l�O!����������]��]��s't�<\�5���q�^EXҖ�)���<⧼ �	T���~��.: �q�I����S�C�ڊ�_Ǽ��ʆ�ѓ7�ZsT�'�.�3	��	�&E�rE�o�nfPl��5�c��uVz��(kR�W�t��ɡm�qIx|�q	�������=x����5D�~ sAiU��b����Q��JC��J�[f�ZAx���|�	�+$l�dW�/f�����!.��5��ˎ�~�W�0����6[/>�]�{d�7]Q}l�ܺ�1����{��Զ�Z�ﭻZ9�yAݾ�F-0������!���:����t�oZ8����������Fi4L��~��:a���Jv/�Ip��UEҌ��;�7kگ�B��m�=mV����Z����k36��W�	oXg��i��?��%�b�
�i�bf�t�1h�C����ަ�uܳ�������ț� ?ǲzV�o\eǩ���ٛ䀠��:~~�����k�&=8B���E�ԩ�=K�SwUJ{��7
=:�������5M���I˛ym~�w���f
;̬W�l��}8$-Z����N=����?秘�Y����V���_'j��C��8����ZM5���#}��z��oa�r�W<�r3<<�����eHxp�8�>:�o����z�^F�7��E��}�2bbb[����V�����m��~��G�}�":�^��թ�杪��"HZ�4V�4��'>����n;L����:����!55�]�M����:eK�szr��;��B��a�a�m�O�@HC�]��0��b�����O��4��L�)I�[k�;����qDh��pD�Tk�_�ߴ�J�,ڊ%������rd�{��pf���z�
"��5�&o �AS�/bߘ=㖙b~���bs�`�6w�i;fi����(���߽u0+xC��
}��Q�a�R�J84+��A��.<���z1��c�ώ�>��Q�x�<|�a^#�h��6�w,���y��@#��yF,~�<�QʿL]�?a��c�;и71���"�20Z�K ł/�q��,}�W���Xh�{��?	�*(X�Zp��so��#wN���ޤk�)\�!$inl|ӝ�o�����`�ֳ@/��y�>�q�'�������݈�O|���	�4�<�X�A�u	p�"���O�x���k��1 �)#0�{��a$�z���e�U���D�,)ÿ�2z������)Q���7�"�?����f��\���>�ٞ�^�sQY�>���ӕk�]���R[M�a��WNT1��$0�U/qF��8ٰ�.��b�HA�A��_�jVv���<n,czP/µ�����(K�s�/�����V'�P�nڋ|��}<F֞�ڵ���og�P޶K�g$Yo����6,.U�w����	h�pcf�ψ��,���I�b�_�>m����ʻg�PC3O����7�{,c'c/�MbSa���ċ6��{c���Ɔ�Y+%�"�i}iR�X�z[yŻƟ���a>��)�iD���9�^w�[�8QIg�ŧ'F��Ws��Y��],�bB�cHF��b��/���|M��g�S�Svs��M:n&* �7��t˱��fS|���~LQtho�Y`Q$!����a�2YN��'�(v/"]-��]�0nW���_��b�@ب�����*��"�zNuU�մ�g`��:6�7���'U%����م~�zP�[voG�x�l�_�U��R3=��� '�ki�1%�Y����:rꋾ'��}8�	ˊ;��шE���Pس?���7��3x���I���>���y���tQ��"��K� ~�.1��4���5J���?��³����J�`$lvil���"B�ǳ�Om�-b��ʁ�ZIY���y���Vn�����i��;o;��=�z�t��u�d;6�I�-zj����M�݁�@�7�<A�^����o�E�U��baY���#_Bmj}S�R���u��Z6����7NW���z���b2k��B^M�����_�k�PP�A�Db|�19�A\�E��J�n�Ix�W4�/>C~�-	9�_�Jɔ�X�B�MѸ�=+�����t�u�������z���4�-�{p�ML���G�,'Ye����[��K��|�$�={Z��%�ny��hY����R2?K\r@�7U�����E��ƐE���
�t|q�����p���O�*z���0��z�Tt���@X��%��'rߤ;��[��5�y���^���=������l3�W���5�̓_�8�w6��/C$�yE����;k,BX��e�|��0�X<�T|�>�?�	�x��I�Q%���7j8���|�m��K��5������c��WG;VY�AIͥ��j�Lש�q��,3iM�SA�a^#��R�UJ_�4Q���7��K�b\�Oc���>L�����g���'(�H5f���W�)d�߄�w�ȵ��7�Z��B������f��0��`4�ܕ������;�([U�=��<�1����l���3]���g{�5�F�i���oթ���g<N��X��P�%���.���A��b��hвq�,���?��Ԭw�j���n5�ԑ�+�\�>?����|�u�t�J����U��G}.�N� `yZ��O�Q��~S�}�g��dF��`�4�Eg��Z��Iډ,�,�U*� ͫ<5X�A4P��>|) �|���>/����R~d�eDC��@ͬ{(�
�>�ZT�.º֞��-.��ao�m@3�����0��X�@w�7Ҭ���`���5:�y�N^"f̼�V���Xȹ���p�[���x������΋-!#wa�e}���]�>�z�iÐ�N�n��1�t��"%��~��u�wb�̫���r��5�7�Z���Q(����%CCjum�����Z�h9	��AGR�Whp��u�2�8B|γb�o<���,��7y�0�� �a 4�d')�;�u�J�����r�[���8�v�Ƙ�l&���=L�R��!#Ѡ��O���Gm�ҺN�����%L��Z�RoYo��r�\����(U��kk���Q0��=4Vv��D�U��0/�!RN>3NJY�h�2-]���i�����W��0V�<�a����7j5��&"��R��j�)��s6��=��~{9����8R�A���e�ݘ��Le�N���0�C��&D4۟:���e�D�ay��Dk)(�X�gj*�Vz�ů�f�t(/~#8j��C�'�E	)��2�M+�ҭ��x��z������֣;�����*�H�V�J���4�~ 渘����w��9����R��h���Z�F��&,cdc;
��Pl��2��\H=�#��i�A�`~/ ��s�|����Se=w������v����[�J�.�č�}HI�tKj��Z����2I�p��ZvW�TN]�n�Ā����/�̛9m�؉D�XՔL9�<�o�0���:uN�}�U7�i���',Pl�_MM,SU��)Z����y@��\��/����"y�-���(���y�P�~́yu� �R<�ԀO@�u�a9沦#��Td>��{ݳST�8����>/�S/,�>ƫ�"���٘!�4��
��4���p��>En�bP�B,�у=��g|�*�9ۋ��&��/�B:����:m|�C2d���l��i9؍��	G���_�<���b��փ����1���i�P��%�ǥs��;�q�M��*�K�4�5�֒ͺZ�Cɻ�}�����Y=u��8{g4�)��~�e�mVf�g��Ҙ�Uf�(��}h�^R)�����M&G�$��m����=�ܨ�{��bT�O&�w���t�ޫ���!��÷3[�X9����E� 2��z4�s���.7��4?o��+o&�7*�8dF��+c?��I�}���A.u��p���������{�?8�È���疠?�7��f{<W���9�5��*b�i�WQ�������o�!K�V����`��
x����G0������vd���楶b"J��]���J26�A92½���C7����n6�d6Ms��)@ZK$C�ᕈ^��5�w"γi��ח�1x7_ '�ZOa�y�}+3�!���7v��r�	���=�$e���e}l=$�?�Y�����\�=��l���zf_��*b-�6�Q��q�Ѻ�n�9�2b���Lc����礓
W�F�c�$�9l�
u|�.��]R{��q|W"/)���}���.T	ٳ��#�T\��1x�4='��w�AG:{'RW-Z@�v +�j5����x���2��l��e��Y�; �bnrHu�Uv���i�
��<v;;;s���18�M2;�[�{|��2%/�U�C���-�
H��f�.�M�'.8WE�uQ7��o��2C9��gIm�~|kj�԰I�hg�75�Yyxŗ�c�*g�nw��}�9m���Y����83OXG��008� �푴A���~PY�C=�u�����_�#5�yp�}�I�� ��w ��O{�����r�_��!�hʯ�l�-����qoڪHp�"zt�̴�6Mr�e�D���2J�I�	�N����j?*���� (����a��?/�d�$�3g�02�Z��b��?��mJq�}����^����#��c2��P�h�u�qq����oE��a���W"j���ǑI��-U��K�[��O��	�ond�O�&29F	�w'ܴ
�%#�+�^���ӜIi��Ȟg�~�f	��M�T�~뗩��{ g�I>�@-�B�X�߀���o�ا�븿�n?�0L`����yϠ!���q�,P될q���3Q �����F�p߈қdK��.xNA���U�aY�Ӊ�7��w�䯫C�����i
��� u&!+�1�i�F��k�Mv �[�:�IbTT������$���ƧjV%����s��aJ��0ޢ��T��"�X�J����]�k���ˑ��b��+��=j-�,;m3���-#��[�*BS�4E�L��J�n=?��p�l�����o�����p�^d�j��
ӏ�b+kk>��'9�;�
8T	��~���2�-wT���46�p�y��4�ֆa�U�6>Rs� ��y�L���F�K��}TF�c��*��$4�_���s5m]���R��c
�>�E��: �J!�:���t�2���4�.�[��mlX�.�giߞ=-G1���6�-�U�Zco/K�+�o2H%2d���u���}����eӥ�i�%���e�H�U�<m�Ư��S��ъJ�f�ce^�?��8��t^��p��0���n$�}`ո�ʣ�T�5 Bd��:�ף���
�{7y�i'��@u��)��X�	�Z�u{�й���F�ۆ����ޡ�̿6�1X�k�KH�JH�N]�<VId~�
�
�2VϾ[�h�?��g򑼅�{yF�L��D�'d`iŀ[M�n&G�#k)�e�K������f�/��=�=�d���3��>�%X����
~f晋]�ӊҲGS����~A�H���<1�I� A����������BDB��k��%*���]Լ�[7�Q��X�i ��whi�g������g�0�C���"��]�f���2���*>ˇߌ�y��.I�T��f,�U����Oߎ�Z�W1�06�\n(e��셔R��du��1N�嶫���h���G}��X��w��q�����~�l��� {���l�5[��ہDv�Az�OnZ�f���;��W�
D���ׯ�"�2O��)~*��3�U@���|����KK��I��È��
lʫ� ��	�S��h�+�Q�X�h���$!A��&� 0��3��vY���=rN:����u+:*wY�����Q�~�I�KxE�EdݑN�ܯ���>!������#�+�q����&��oԹ�T/��1�w�����_�Ft�D^����2Y�����6�9j����%hRH	Rތh��A�/�`ۛ�ra��ZG�����=г��ExM<�y��=\����؇��%�$��w�N��d�u���ۄ{PN��b���+����Ne���
�x�{��r����}]���Ayd��?�sh�������L�\1�yL��[Sz�G��&=`���׸t,;��fɄ-�M���۩<�K�^�#Veggۉ����o��#��u��S�S�B���� 0|�W�#�ۗ���~�&�+*$��ZLj9�:4�8�!G�T�S��7ٟmB&�L
�Ǆ��8���M���RE����}]�R�lW�߮<+>"�>�yX�yd!��X���
?�c�������s�e�R��rX��Q�s��9��3w��)�E&�aQqp?���� �5#omMG4���E+���%�?D��x&0}M�d?�h6G9��
�I��%'2�j$0aHj����W�t�ϓ��0���:!|���Ԕ*Y��g>h5?�̦���Ŧ'
�:Q�εg'�"�_�,0�[�@��\>\v=�,ϑcǅ@�chB��a&X	���O�]>Թ�QK˸*V�c)Z{4�-ځ�?b�m����6���tE�BD$)�_
�hmOMi�H�1���7^�+@��Ƣ���'+yv[���$�_^�&Z���n�ݑ;/B%`�%��}��UZ��ZN��k��k�Є!k�u������Ac�9�z;EÚXD]� �}�͢����Ï����GD>��]<���-f���m(�-�)o��?��t�����C���|�34O}K23^��D�;&b�v���T��E�M�����Nf��D"�K�o�-�;k���F5C^��蠲N�2�^�8�U�H6�f�����y0K���ڰ
/թMG܁�z��&����[���d[����)����.�6Vb���AxG��YKl�W~��wH5 6��h�D�L��jV>=��( ,�z��o�MR�`i�Y�[����ad��j�HS���M2b��[�xg����Y����3)F�t����eN�ZK�%�~ �w3v�eC��?�ʞ��&�\^O؇�x�r�:X��XK��u��a���3������[ʀ �jM��K�q��F+D����|iAQn㡲�ڽw�����ɓ#�1�/Mg�O<�;Ӟ��36�c���#�߻~��_��k�s�y�ʶ7~��L��u�w�T���Tt���s��%:�Q�M=��=���Ԏ�Q�H�9��� �'�\Ȣ���Q�p@���� �_o�H�n�/"b����v��*�5��>�f��S�k�V��y�:�W-�R��_�AY��qxxxZ�(�Q�Ry�������A^�����
G�[����73�3�#���7���N�5!j�z�r�󧟣�\ K�^�eo,ӼsЙ����3R�|j��j> �uW����N�`r�+s�*�Pur���#��*1�h�]��+ a;@ݝ����7�8��h�!d'�E�@\���l���On`��^>��K�42D�z��=T 3���l·">,&�Z����&b����a�#���o��J�ť�d�\J2Uq�f��jL��3-���Xz�Q��2�[��<�C�Y����Σ�*z����ۓJ11~/1�ꌛ�r�Z� Ֆhf��*4e�h�P��Ɓu�/��C�f�B�?��o���Z|� �m��M�^��)�7ɗWuum��~9���˻��֡��vl�<l[��$�S�e�+ü4�z�ś2颕�^l�.� �U�
*C��g�9:��jh��yB_��;(����7�CP��M(s*��;� �5���L`}ZќM��|��[��4�
�����* ����_�i���/�ͯ�ٺ�a��o�~[g�(�dP��Ö��m���6�0���xc��_e�Z���|��ј��C��X�4�FJƄ�:I���S[�\�z�˝�_�����}UqAՇTtF�V�l�AF�;(V���4�uǒWP�b&�&ɡ��c�V�4����{�� m3H�VW��*�ÂR�z���VX��� ��k��׊&=�"�|4r��ׇӏ:���3�$,�N�@���#e�����W��y�s������Ҝ���q�0��<%epz���+�߈]D�\�OqU�X��3��a�QE>�+���ER}�J��9���R��B��G����c0���b|�GqV�z��]�X.�0��8��Z���U�1�o��+�˃�i��ʷ��@�����Y�㖐�o,ٰ�_"����<ǣ���*�M���,��i��	EqQ�H@WH����{X��ƓO����P�U�uum֡�ݝw� *+I��9Ľ/��A���I���i��s�v�G����Ɇ���_y���.�x�9t��\�#BV�|I��R2�������!/�7�j��G����ΠoL���������8�:�%�4 ���LH�۴��SDM,���+5ni�-��8����/(A��5����,f�3ʤ�ʪ�v�����p-��喱Yl�?��X�C�;sV���N������l�] \���&أ {(��s��j�Z�ϴYzݠ���CV�D`.�Ğ��'��8��}������$�c+�F���~�����~סwU�F�w�iC��\>Eq Qד�9+��}Yh%3�/�U��^Y�Pr'�������c��:�;*�\�0n��@�d�'�t���++b}]�?J���[���j��(YԄ���k[�w���E���%H����I~��/�������ͺ숙~�d�﨏��L�d�%6%��/�*d1'u.9�|�aFS�����)��YA����d�? ���>W�)E����t��x�~?ow���#ɳ�VÊa�`��B�������>��6�9$I;������?�뮭�����Le%wq`J�~�d�E�v�-��JN>0>�Y�W�r�[��X�~O����"����l�5#G�83k�{
�Ӣܛf�%L�?q�|����~���)<T�N�J��PG��Ki3�����!�/� �[���D3ؖ#�}HL�3�᛽X�����Q[�n_|��O��!�>�v�9�ilSb�����@��y�-fI�33l�wG�;�j�����s�?6��;�bV1��#���y(ՇRfU+LJ'^"�B��vk������B�	�$x1�uy(j�`����nce�m���a�Cf��l�ڿ���2vӠ��Zm7Z��H_qZ�P���د���3$�v.���.�SU����;�ĐrD$}cٷ&P���y*x�Lw!��rlHL��a�8��>�tM;V��͍��D��W�c'ݙ�<)�>N�jk*���%G�8�4��wR��w	l!���`dR�AW��$ʿ-&��f����2B�������o��.�����_uG���o`YC�M5=��$�z�H�.bS�sC��e��/�Ї�Q��+��+�wD����l�k����'0��C���\!��P�)v�{Һ��u�S���,�>F���}�B�� 륧k�$B +�-E������>�j�A����>Þ��a[~�����ǅ�����]s��~�5�3�UpY�xw�6�	M]o>rh�kV���:w����pu�l���Hxe"oؗe1%��P'U~��4� �
��g*�&���c��3�b%`O3��'��y~��TOl5{3���wm�s񀟯$d��*���6��*��Dx@UW�*�P}�5<�)[��1����Ow��u�]�LH8ӝ��!j�%�_��ܗ�2�`՝���tԀiv]�C6%d�K�Շ�H��zt�w���Q����7�e^�.^[\d�пEZ5�<j�����IV)�ʊ�����$�<D�-��_lB��/3{��"�0��bp"ry2+��A'���K\� �jNy��:�H+:��蔳EQ�[���T��q�n1s��rx3�\��W���o���R3`��^�~r�O��5�j�H���Wj��w_����?t{0Jh�A��+Xh��L��`1}j	��5z���'�A���#�c�d*� 'A�\�f���#b���JKP���Z��9�վ���'Z�^�/.�98�r^md������2�x�.�n�φ�������YG�G�������'�)@9�����/�@)洆�D�)*�CB<��O�d��H���	�5��ʀR'|��uZ�%^q�W��N�X��n�ⅨXt/Cg�bݢVp�[Y^t�+m�A U����1MF��&O�3��-R��Ӽt7����d�4��aZ]���U�Ȧ�B�c���{�Veo�a�H��J\ȣ����oRk��s%e�[qi�%|'�;+�3_rX�
"vGNW���|��7&%���ߤ��k=11����m��:#�������?ox�+8�/}�c�}ߒ�튉����\�*��A힇چ�s�033HW�?�%F�UZ�k��R2�t����CC�({e������e	 �}�s�Gwj�S�f<�ƭ�$~��O��]��J���B�"�ɷW�O�ϮAM��i"�sv���"�yS,��=r��s,�L{�5,*� �p�  �L^8�ԓ���,B����*_�7�4��/�3����42M|���8�8'�+9�6�%�λ�/�z�k`�7���]��J;|�S�5���A�m���������u��iR��,P�&��zR*�%"���B�kfjI[����c�'����B���<A�T�°��${ǩ#s��ܞG���3�U����1w�L�x�\��B5"�mV/G�]^�z�2����o��|�g�����si����?��z^{�B�%z��]5�+��/�iXZ�T4H&�ht���ڣ |�Y��x���,���0PG;���0r��i��2�^��l��x�Jv+�O��N)����T���<��FP`��%�o�!��&���Am��ky�%�߻l+�8H�l�
�/��Uz@c,�ư5!�8���52ɣ�����UEX��ӷ9�˭�,��M p~�4i+tకU�-]#�l)�GYQG7���Uo�>}Q 5��M9�B<�J�0�d�w�8��Ȩp4�:`x�:��j#���^�A�5��Zxe�IďjM��s�ƹ�=����x�1C���"j��dk�oӆ�j��S�������^����l?��-5B�yW����KG�5)R��r�`��XxAԜ���	�����wrN? ��YI2�����L3[�r6��V�u�?^��A�a-���R)i{2pS���f���~D�~%���
��(?V�s���wS+�����_vU���c���T.)W�q��`
)��oը���ϯA��s|�Dt
AU����%@E�J�,���U�^��39�t�HT����v��<��<؝>TD��-輄�m}��Lu=+�]�l��T�
�ɡL$�u)#EZ֎*&a ��� ���?��&�'��X���D���g�j�%��o��	_%J����D667� �� �];�=��ڜ
����/���E��VÞ�y��i���~��	�u��MлFz����W�4O�.O���eӬJ���9��b{�/hxfh��)����wp =s��c��Q���n�v�a'��)!L!����ϗ�,���Pwi��6_�dD�)�5 ?����p�X��b�R��|���!q3`o�ޅ����� ��]P������ya�X�p ������SI����u)|�c_�(�7�#������O���
��zz��(���P5(�X1�.�bU$¡'T�-�;�FE2ь�NM�$���>�UV�w"��[<s}���d�=��rW����޽�Ks��V��D��{ܕ{7�h" �ń���{%���^�r�i��>���0�Hr�JM�(�[4�\<��'�-=���=�&��h��l��aLs"���?�k��~1 z����m�*l�a1���?�醙=���n�N[�k�Y�e�"�x�U2~���O������A,��G���x;��nU�����Z��˝�峒��)�e%�l1Zܛ�Ȁ���i~7I�T�2�z7"�-� ���C�
��_蕼_�����0hU��jv�� �������g�t�Ǥ#P��󿷋(dǌ�\��rU_�P�J:�qD����'�<��H�U���%�]�TUN�`='�T� �=��0�
�K���c��6e��Q��'�N�+�J�!�c~����/�1�rd،p^���"��&�i��pcƐ�ꧡ���K􈾟=��{�@�`�Z���N��,x��������p��%������̻wr��ܹZQ����� �f��aU�K��jcL3@�̟, �U0��L�k���>�YĆgTH�w����*K�p�n�=�4$E��P�㷺l[UxFtlp 8WA���Y��-��g<e��yNd����$k��Y�ӈ𻆉�(��͡|�����v���"��ѽf������
���'ݖ[�'�I/�oз��wV�s�0��u�k�ul=Z�r�u̒���	�K�O������{�z������m޻�,���j^/���3�<�}�Y�OC�ugm�A*D3�8����q�c*kz�Я��V��r���lR�{�k���/�sa�+6�t��8ӎ���ƔR=o���o�)�0W'��q�!��<�ז�-�8�,�����;�|��P�l�g��K�❱�1]h�4ԻP�yK����>�[��/3�������Mw��I�l�D�>s������mp�޳�59������r]5uuKGG�TU���|>T�U2��ꢟ>�Ud�2Φ�����Z��l�
=�K��T�4�Э�p���x8T�w�b�&���D�\��4#B]8�Ӧ%��y�A�s5.i�n&�>mU'���5��j���'ٓ>[���j��C�{\�d���a�����#��N^AW�nvv�:��Ƥ�ώp�Ʉ�s�V\�櫛�\ѹ�w�[���_s;���Ͷ�����!��N��W�P��eb H��R�K�dd�.�T�ȕ6�Ȗjk���ՙr]z���;u��r�	�&`6��s���ɔ+Gz9?�oc���L�h6��5�W�iu���1�t�Q�:2��'��:s��>��a���r+��9�OBU�n�t��m�,����9[^.�5X��e"I���)5�;��[s=b�g�\�M��L`'��ʚ�bᜂ�~�c'-��Q#M���Cb��el���?G-y�a�E��������'^����QQv�ޤtJ���t# ) � !�"%� Ҩt
HH#��J#��H3C����u�\�,������>g����~�����w��qț����Q;����kO����[�$oo�������K���"�|K�= �$}�52%�nw���;����eec���UϜ�0�;���0�7۵�����A�����,��MT��~��"MJ�Ŵ�ʮ���S7Ѯ��9�˲)Ͽ�l"���#�:����aò�sM��fb�����ô����Pl>~��S8���63H���	������6/�:��S{v�EJZ�.o,Yf��i�#`'��|�QG$J�J�'Xc��\��d5��#���) ��K����Ff>��}� �Jz�7�X3�Gk9[�"_س�E>f��Ń����]f��𴴴\dZ�Vs܏���n>~l��,��a� ���ii���%��@��̖Z���xD�R����*"f�r�b}�-R�8��}��Q�(s�!9�)�۽��ז�8
�Ƣ��.�E��A�������>�2-H`-G�tF��($���w�|Q�tGw��+a�S޳�P˭NP������hL���Ԣ�� ��Ym�Qm4�	&))��������e�qV������#���^���с�Ч �gnVu7��ƫv�O:T)c�Q�n@,��\�fJ�H=<<$A�ÙOC�i���J���g�F���fJ�ah����u&~��x%&_���}d������s�ǣ��e���n�<Z�C�]�<��c�rE��褁��V̧�Q���pU�i��3ㅯ�$��4t�G��� /��uyN��eL�f���6"�OMuup�f�c�K��(d��<OcZ�Dٿt�44;�ҠW�/)�̄3o��T����T�^W��2q���Z�tKv��6�՗s��f}b�@i~pr�����rfaNk�]�f ��2j7ˢ�C|n�+�J%�/�4�e"�+4��-�%Pn�ʆ��7���^;T�jO�trf!_7��q��I�s`�m���ULrQ���|j�Z?F�+�0�-����+��u���[�'�9���?g�m`X�O~���z�9�w����܁9]�����s�*Sh��U���|�s�D6�)1��b�[+��>Z��b7��k5����X�9��o��k�eh���0��Pk�?��D&ઑ�$��ۡ�!�S�mmquuO<�lV��D"�ūm��UU�Oͧ� |Y�#��o�t]�F�ܛ����L���_ m����o��j1F<���+yLo��Jj�'h�_��ԧ����3z��7H�$�F?�]����^<�D=+s��'l��w��(¶S ��"��5��ȡOG$���x�@ȯ`�����>�%_��)O��c��4k�D���I�(U>�
잕�;���X��,�N˿�Z�)&��cҍY?�.P�g+���Cͻ���d����_SO/|��n�c?�tuu��^����>h6���Ԅ��ޡ��u>�WCS3��sn�=�A�Y�Q�^�-^�3vK�����@�Ufʂil�3;�����9�^V�:�N��B�}8��YT>i'��怲��A�!E�x�-&F2�f02�e�/x�
<�7��c�#���u�1�����;���>�Pbt=� �� zSXD�
�1�/��X����67�.\������nF��(��<��HWF��]��ߠ{�3a��@� 􀞞��x�bjj���9�/�y��@�nY�g�St�C�`�@jNN_��4:gL��莎�]W�*L�ြħ_>�)��`~�jÇx�9�����_S��wV�J��d�AZ7��ٞ�*���~���9��b��Kk<���q��M;��(�b��%4Z+�mt��ay�ƶ�gE�������5�N<#r*@�T��.�\1*hZ�L��UiZ>�DYZ.E�l� nĽ��M[�oib�e�ep�,�%�7��[�����M���d|q��_  <<L�-�Z��@7&��� +,Je��g367ﻸ��%�>n����Y�' iMZ|(6GrPp��GF�M"����t��]��h�g����HI���h���:Z#hF����A�G,hAY��/ "�(����f���lŵ�g����׋1�x�,��p^�%�E" ޘ{h_V�;П~k��SnI�F�O��A桄 q�v�n�+8�nL���|�飈�>��w�]u虁�3������66��L�y˞݀&605���q�����z=�1l�A>B��T��1]a�Un��z��O��F�-���#�S6Dx�����W*OВ�2YŃuٖ!b3V5*;�H�}��X?��4�����~�F�ֺ�8d�����}�S��c�ZksZ���<'ǳ.j�l'��˝�J�S���������>�r{��c������^*��r�g��ֺO�6���}"]A���3O���D�f�̓�`�吻^+}�;Nd#:Q!~�h^mF�o{J�k`h�17��I�#]c�/}�X�G)����)��?��]Ox*���x�+�C)��{{{��2�T�"�U�b�S��`�Xꅗ��\̧�;MJ�j�=�o�}>��J�1�_��{�>��*�<pd�,�e���a叝��|��$~U˿���� 	~�����b������`��қpo��^�B��%T��`�=�!"��Oaܟ%��9���Qr�|ի���ᡈ��>�7��m %hii���-'-����X��ֲ$i��o�f�rC�u�K���Zo,}�����|c��t���� ��F��CEQ�FɽI���ū����l��?�y�Z;-CstAA��ј��7Y�Zw�Ozo@��ˣ��C�J�ls~N�ƚ55�2��~��C�rys����;z���@�O�(�ڐ�� r���đ�;�E�9��Z��&i�o��Cȿ������#\gD��a���������r���wAe�k?sO�M���F���1A�t����,�JMH���Nhe���/%��Á�����ttt��<�4n'V�����Gypx8o�é�M��+�N\�z�<6C�J{,����N�A�rV�
�ɓ7y7�Ƙ8	>��*��x/SD����Ҩ�9����$Zܺ���AOi�$����=`�Vf̀Q&E��:7%H^#s���� (X���M�8Qա�;�ڢ����v;��/N����^�&f  �tG����4r�t�����f`b�`j��'���P<����s��t��7s�Е��K�r�I��vO��oZF�LUܲ�c����l$^��_nk�9l�nT,py�:�ȥ{ѝ0����\+ڨ�
p�n�~|i ��hG�e��Q��y�=��WeQ�L���g���۳?~J��}�nnL)��w]�����%�������K��P�w~/�Q�E�cZ�R5��+����^6�{�ō���~h�������$Wpct����Oԛ�����f �	O�1ȀO���� ����INIA� �D7����(n�ۘ�r`�%������H�p��Wfw����i3�+i[�7V8K���F��_�џr����h=�v���	t�l	8�ep�K��COXxE�O�G��m�;a=�@2��F���uV% �~�[��%ߗ>���c=�`VL�2���)���:��R@�A���%�γI��P�/�^>MA�#����m�*����p�V/�}ח(�?�9ܢ�����H��@�q�L)/B��cJ��0t至�}��S���w�s��v�PN��p�q�*X���=t�2�8K��l�Y��H��|���^�^D=�gߓ�����[w�ۥ:��";e���Z�k��j���K��5�z�T�f���N2~gBcsJj]�Oh� T)M�����_pnb\���-ݭ��L��y9�_̅DD��RgȖ��(U�I��9��?�)#7�aNh�$���Q'j)p����Kv{7���R4�E0�[h��<?����:�Y	�u=���voڃ�`�E��������^��MlΣ�~�]��}BV����"��~#�I��%�U��6E�#�s;�q52ɳ���yG��`E�N�����I3.��Rh��8����ӿ��j�u�B���G�<[˷,�z�<���b�;ńz�6����ɴ��2f�徴�ѐ����L�&	���M�s�g(�����bk4��ň�����m����h9aǉ`T��bum^�*���XX�2jE��C�,j�S}8x�z��NAꣃ��W+�?:ۦCͱcIb[M[D[�����&5��j^����|�Y����7���	����򙥚�������b����b+���?���i�d�>��������>\����*��4����1��/ƃ��]s����\�1�����O� 	neoO@DDtv
sAF�_a���S���ښ߲�����Kk ���םD���_O�]��kQcHB�������o��\�>�]�uchb�6v9�r�=���`gh;lv!�Ȟ�i���������.�M�,!M��j$�"��;��l��j��^m�r�v��W�/뙮�����S<i�@���O:9�ϾȪ���Y��6?�9Io��u<ʬ4;���<��I����� �c'��ߗ%���o�<�n�71�ۥ53%���A��pX���ry��xԫ�]���4	{,]W���'�ª6�L��ʼ�
�^�����5���0�@]�87���Ah�ǁHP��5���M:���y�(�v�m(_�.��I-���gE��6�2���w����MЋ��vpg�>4)}����i�MK�S��fg�ox�+��kvN���>�D�ܙ���E��:�����3�U����w|p�S�l�8�7,��\��)�uF�?)DHOQ��N��((���oֱ !��	� ��l�To*���$�ഽ��v��7��-���=Q��Z1�����P��}ޞ���$�Dm�ry���8n�\�Ϣ?��%���{�������Sy��"��*��Ȍ9l�%>=�t�<c ���\ox��:�������S�r+ƪ�>,�zB���g�.G�ss}yvs��4����O�a�ێ6l������4�z�T��>48��oӢ/�옂�`�~��<yA���`�mgC5�;! %!	h����X�G���}�� &G������������e.6lm(-��dI�������^�0��c����uO����tbYe%��.�ٿY�u�N JK���f{d&��!ٹ?A�Tvd{X�_f�M�������/��6��cjhW�||#�)#���`o��-����V3"�55��)���hU�Ԩ�fF�cnݐ�MG�Ю����V�ǩ���?>�=�yJ���5Ɔ.dd@P'Mz�#/3�s�;�������W���=��3��%	b3QOڭOV|��4�^dț�i�"�q�,�������Ht�1Q�y^�M@]ԏ�����M�IK�E���=�M'<�<�	�~Zi����1�gs�L*��� B~ڍ�d���#QMMM��.����=neee��b�;�+�-��5���OK��Ùە
��W����hB�>CJ�wW��
���-�t3]�	������Q�zf���{LWm���ee��}t��}p��'9^�����@�W���N~��g(Dk�j�]�����]��W-7�,��⻊=Z<�����떖������E~�������#������c�LXO���� 0us����=�~KUU���5`7�I�T�rc����;��y��&���m��w������R ���Xy�G#�(��ió4�A���c���x�f1��Q�tKU�^䞴IVM�7� әL���1�K��ǺW�Y=����wa��G�e�I�ʪ�Q�sjm�vn��:uD����I�O1qh�p30�Y\��)C�! LЮ����x����g����	�o1���n9���Y��� ZP���g����Scs(x����"��-&��-�7�u6�����k�h���G�1�ЈH�,��!����s$_}q�}w�Ҕ*?�����^�zD��+J�������@���O���ݲ;�+}(��\�����!~��!���zB�k�Jp�S�o�L���Qd�U���Z�*���=�S��f����L@�W��4�w�_��-�`�����j��Òq�h-�Ǉ�u3,�{Ⱦ�w��r��q����޾I�AO!�M�Jr�%C�D�?���_�-��� ;<�7��%���NH��=]N�����8x���c���ؤ?fXnoq������Qߚ��gU���L5N��7��\����6A'�Qu��x���9�w��F0]��oZ���:Z�̇�U�D
�T�o�(��w[�gp�@��ΰ��9҇
���#���.�'4w�s2e����=2b�-�^S:Y'��/�Jg��7l.�cuɞ�kP
U���s��N[~�:֏�}������1�T�y$�o���_�l[��f�KZ��ze�6�[	~�Sc;R�4h���@�����L�o�R�p��/�`����eHN��;�ݐ�C<w/eCC�ik��Y.�M�6��,�!�Ŋu�J��ٶ؟���G������~H\t*�_Q���ґ��n�R>��!�h�Od�W����^�\��| 9y'N�����F�Zb��U`�i�(�b�Φ�T�������_��my���&|P`�M�P�K�*v善�yź�er��&��9���}`��z�?�!�XhqĶQ�fc ��Лr=<+��U��
����Ϲ��N-�M�+��-�y��/��}�����ѫi���5It7�(' 
г́W�uF��U�q����#�,��L[����e�%���NP�'֖�.���FKԷ�͋2E��O^���z���XI���T���GL΍�&^���yէ/,A�z����ux�eAv�$����{Ƨ���"�~=)ƱE$�/�� ��|�(2&oo�������y~o$[V�%��2�%��A����[DOI�@��8����j�H� !��C�a$Kn-r��-�t`�.Y+�_��� ��������ȘC�;Nv%@!�o(ۯ�11DEE}.��ai���R7oeV���њ��Y�ou���ߵ�v�����Ԇ����o��-����k�5�Z�F��#�����g�[P��{ň5�u��� �v#Ka��L%������њ������r�痊v�	B�.6h
�WK�Q�`�9�-����8�D	6�|���@���_mH�w��Q��2����ƈ����ux��e�E1���K6 A7+7�skq�f�����)o�._^�1ږb�l�4����AK�z�`���0�rn1Q���r��)J=Օ��l=KM��&m��!��b������	$�.I���QXT�1���w�i���V�j��x��B��rR*�'z.��H�9��U@�`lQՐ!8wKWՔ�$cN�+��'�uƨa��ɝ����m�ݚگ�.H@Į}Ք똚�Cgv��C�㱗g[����f���^�1_S�^{]���dw��5W��_��)���#������[��xv��T�-&7VT�Qlz4�]f�vA�J��{Ԯ�G݀];��<q�u3@����!���U����:Me}����C�B�l�����J�!ᛂl����G!*�(�fe#*��{~��U�(�����Ct����� �HH�k��"a�B33�������0��m���ɼ��Cd�gJ:<�kP[n�����.�!e�y���3�!� �}tg�8F����%*��b�����7�zfO�]�cM�>�-���ϩ:-8a���~���CԦn�1�f�*��z������p'?�ۀ�Ҡ���oNѷ2 >�)�zoQ�;�ēT2"J����|���\^b`��Yf��J����7�5:r������*+��+�F�R�t�_a߬0�`��&��|�!1�3���!�,��n����G�o���V���\�{\`hi�k�q�K�!Ѫ����j��:"j3�BT����cv^�.8�H�ǌ������,���$j���[[���������|<r����Cd��ZE�u뽚�`��/���}'�)�a>��s��v�����O���ؖ���U��ꎠ��z����N����b��_���J��"�J�W����m�)�X~��z��a1,��[|Z��-Z~�P�̿9Y��ߪ�Ř���P]�R��������X�3iV���{3���āWk������o�))uW�X��ࠗDd$:꼠��O̬�u=<U׉u�d��Meϛ�&�H��T�2Ƞ� _�ۉ8�MU��*���#�����M�E>��Zܶ����I�5���G����E"�3��c�]��iJ2�o���2?ӟ�\E��ߦ�q1O�x?Auv=�q�U�dUעd�G��\�r��/����M���5i^9^�ݟ��Q�̖ `mq{s��E�o<d��3ݑ����f~H�� �I�����*�sw���9��$�O�x?Ӛ�;�S���pU0�J�q��j����O@rm�$�J�8/m8�����Q�i�|G;#�L���r�� F&����Tw�Ӝ[|����}��lH��
6'k�\�p9ܷ��U� ��O'��c$N��'��Qc=5�(txS%�A�X�E-��`.}Ukn��-���ڪ�)r�~u��C����ׁ�����ؿ�b��x���>-�����KA�����q��.�+�����)��U1��Sm�q)��;�����4;�\��d�a%�Z�O�hꊒ�֗�Lx8(*�qkQ�R�2aΙ�>n��I��ק���*�r��S�����+Vt�b��� ,0�R�s��b��ѱ;3i���+�'�]B���� �F����?�M�W�E!�~������֜�8���,8+=X�P���L����&=M�j�^�
c��I��d�t�[C<w�H��g�僕��[�z�����x����ߋ�����HI���^�v�7To��#\%������SD>�1�5�hee���*w�Cs������?����d:�ު�W%6M��g~��ڢ޹��9�<�8������W�j^\��)8���G+X�����H"��ܶy��B-��rEz�WL�	�,/6��9�R�rM�_��� X�/�^�:n�j����	��7.j:W��w��`~��f��'��[-��������?���������(+4e�8mgV�~GCm~O+�.T�w���a~�%O���G���ˬ�Rߪ�N����3��̇��z����dy��&�k����I��FF��IŜ�)S����)����.ϵQ0����`��f�ă�����?m�}�S�uj"i݋�����؟`"�'D�5�1�$��<:�^�( E����t�d�����b��b�5f��Mt�������t(�P�=X��)���	6�����T�=S�����إ&�
),|lx}�xs�[m�C8����3���C
�Vf��jU�M��[���`�sm��r��b7�*�>�_�EY^���w�7�nj|�Nl{X���N��i!�ǟ�����s��@Q��F�[�f�`�e��b'��L�P',�LS�R#��)�"�����]{V!d� !���_-��+:cF���u���e:��Ԝ�ِB��s��@���'�f�^��J��ճ8?\G��/�/ ޛ���I)�OX������N�����^x�-��G��(��O��@�X�����ß���f-r�o�`�'��<�+����8���W��Y0���u0WT��%��ή8�f�4>WR�������ä,Kه3�ey��F?&��(�JwB�I<g�Ti#_=��Rt�Tx��v$�'�Q��	&��������P]h�����P=��~���?N��I}�X��5̻���J�f�V,r�l�1B��yx,	-$ ��'d��N�$�y�/n���3l�	�M_�M���,�ݼ�B1�W��'����D�.���p���T�C���>���J!�C�v���S��(�Ɍ��7��w�2��u�5&��Z�!?T	���;Bg� A ����[�(?i��Ӣ)����Z����s�:�	h��0�c��~��&���zc�<ztn�C<zi�����c��h*��3�'���/:x���T؅D'�F��Oʹ���E��^E�,N��*=�F��p��k���^�.2�݁�V³(��oS�ܶ���A1!wi����1�=c��x�j�:�C�Z��x�^��������9a=x����A���X��^7���#g
����0=�	�H^Ϲ���ִ�SN�M"�����G3*�Ot�L���E���!�x��������S�z*�A�bl@��a�-gb(Ѭ8�Lp��ޠi#=��B����_Qe�3���#��,.�`TŃCD:�!�|��(��o3K�W�>\}+���K�G��+���_���B�tO�Y[���������B�Z.�p��o�yƂ�M�����WxC��"���xB�49��W�W��<	mEn�����c9=<�u
bQ�����s󌸼�v��n�%�*���E@�����̋�D���co[
pCX,��=�����=#k@'zeWT�!p�� ��܎3//�y1.��&��Yl��m�Q���oi����ʳ���߰�UN�#����bhi>���_�V�f_���Y�U�t]� e�2�9Li��9P@`�A5V�Y7��Q�����O��W��Ab >)�h{�8|^�g����Q6ч��n��f�lY�Y��IIP����d(�fe��P����W1��3/��y��o��rx���apOQF�{�D�ë̇���Do�����N62\���I����g�kS��ëv^�*3n /T[�1��%�D<IUQ�D<�9��!م�Te{�%�CĽ	`�o����hR(}�B�����&�
���0q`b�×�"��ԃ.����#
�?��/�ݨ4.��"o�B�4���^���2�:�Y�1�|խ�6�B�/�lE�˸�┲|�~D���{�Q� �(����lO�ݙZ���Ns�I���یc����*�~N"�z�=�sj\O6�"���=��l�9����T������s�w�o`aV������ �R9cD�a]��)�n��y�L"d�����&_:�8���h�N@{���Yp�f��ч�l��(�Z6��'��3�:�N���(�Zh�K���A�t�j	 �)edḽJ�X�(���16?�&j�
�n����Ҋf�<.������N]~�\�u�##�`q��61J�܈.��I:|VY�-t�!��c&R/$Ȁ�y���:�'-�<������B�XxF��$^���_,]]�?)�W�w� �e|�l�xӃ���}��	�I��Um4�U�LC����߄�H
��S��D�;�u	ݫ����@:g��[KII���� ������`	���ѭ�����_��U1F��J�0@��)狰��|�E�:e	��Df��v�����������E���]�&�e�mMCj����d]�"�.=�mᘘ ����N-1�YHԛ������vG��w��|�SE]os97���z}m����sP(��f����yU��䫲���>7�H��Y,��6K�6����V�����u\Fi韏��4h2F���C_y��gzD�k��K(R6j9@2�/�����}�A���͵�%����g��XIrb$i��{���u�;9�b�����{%�%\�"���1Z�M�ۊ���� 	��� b�XQ\�Q�/��͐�[��j�H��U_<�e*�����+++�\گ��]c��A��!:�������쏄���O����-�E�bh�.4�8�W�>��m��=���'�����c��L]}�|�_�"�<o�/�8��J5���&",�H����:�E��@A�'tP�	Ff�}����+��J O���p�[���4/q���	]7�3aq9��"T�g%��d�9�_���q��R@�چ���^t��ϸ��z���K��i"��l��q���%�8B�yYZ�C0��������B�{���Q�O����bp�(�p=�u ?�Xd b!fIf0=H"׾�aW� ����љ�=v]�PW���ʤ��� ����$}�;,��<�ʕ.���*'	�XL	�T�*���|�T2f�T;�����ڂ:f��Av�N#��s��_@[�M�m��<���*8Pox'�U�4}����O^=���Y�{��}́)�}��Q0�vƓ��4�Io9K������<�"Zm�#kV@
�?y���矼�AT<J}˭wjH5�ҙ�-����ᒬ�8��ae�ǣ�B]�ʓ��R��K��Uy|�����"D6�fsW���g��j����%�?C4V��P�&��ԥ�Q:�O}�@G��}%�K�m��b~x3�nl7���MqG��i��H"H;s�"Jͯ	я��F?�O>l.��<^~28�]���"K��y<2�t�к?\t���Gz��mY�ٚ��R����/+�s� ���n���!1�!�̋�}�5��D��}�o�4Xib�f����)��B��*�� b�$�
2<�3�_�Nt�d5u�e�����3���="��sOW-w�%ۅ�g�s�(�mn�tSw���������x�i�J99iD�����-t�~s�95��I��:\pRs��XK:�w�T��2��6lyJ�vt��K/�
���+�/�����/�|Nb�o|�'wO?d���"�C�=W_Ա�jpt�r��[7��Di�����eaP	ٴ�T�V���2�jD�??�i�LU��Ej����?�����t���Q}�We����%��@ �xcw8	����X�\dJ(J�cs�����h~,-�r���r\�~ɍB�'FK`�gK�A������T�h��`��-'X��(���\�
�n!�)��餪�V�QV0x׭����R(}u+��������o�wR�_TD$���FIw-�0����-�«��W�9p�Y����ӉZ�c� hP�����5ml��T�ת��v��p,��z��l��&djJ���]Ĥ�yMMtCCC��'�o9Ҹ#-Y�8�����3��)�k%�lm�B��n���))5� v~�Wݖ;�0Z��OʉE9}^a��䎚*|�Ӟ���z\Cq�N?�X���Ċ��y�+�Ԓ�hP1)���o}�b���h�m�<�z�Ѽ�F"���O��|�q���&:�m��#��o������]*�ݒdz�O>P��魂Vg�μ�w}�~\j��d���:v�s͕ţ��H�A�*c��?Y	HՁo1�sBx�^���c����M�x�������:�"BBA�x�,L�׭���Y�'�����r5�B�Q����8w�_}�r���́_u���z�mN̥�{D�ſȟi��$=e���I@v!��ܮ��dN&ޢ՜�fȪ'����m�\�
�Tl���nu�?�tY%p�g4��0}~����� �R��[*ܦ�\&w��7a�����e�GO�f�c�48��+�>��?0�Ls�*aـ��u�,��+ޛ6�Y�4���d��7p%���¨~�������	�zKr0M�ރ��]K��CRF)�R�
����?��4�O�o�9������o�n��n ��!�9D�+4��4�)��G#�a:�I���	�r�H"��S|=�@z=��h}cv.R�؇r�0�1��I�k������0��M��*�������������)�M��J�er#����bI�&���#�ϋS����K�b+�{Q#_ԫ��\w9|����w�0�V�d�wުW��@�j]0��7������&��oV�xk�4�u����_�I%h�_"Y��0w���~�m��b!�K��1C��+��e`�3���E����|�	��5��EP�B�ʷ�b�`v�������H"�H2�p�p!>�S���~��z[��X�©ߊ7حd�W]Be���u�7�T#�Xs��X#��
i�Vc%��a�\�X�Vթp������?���Tx־�P�?i� 9��9�'�����/�
����ޥa)�G!,ϒmF�P?���$�,]@�y�+�eQ󡽽/0����-�<�l~��g���57�q�s���={hm�}�`}Iz�q��#4"�K�������T��0��u����/ة�}~&�V��N9qs\��oq~��~D�X�.Ǯ���A�kĒ�*������&�V�;�:#�cTr4���܍���ɧp{/����e�УR�Z��h\����7k|0�ü�A�H+k�z���S��ܦjbX�S�KK�����X}\���|.�T?=M����N��o a��@�7�&''Yi�}O=6�Qf#]>�t0V|,��+�y��>�������18!?��Nӵ���d��n���ɮ����2�Gy1��۝�d�t�m��}���s0+���v�/A��}B�mx��JZV��Jr��$i�W�9�u�,��K\��$�L4���bD�Q�,}�Y���E��;��¬l���Ȓ�I����NLFc2���c~g�B��ɿuuu�0�l�{����_L��͆x;~T.��NON��lc	n�*<����\��v��{�G�[��<Wko�����w�`������Eد<l.:��GjO��J����o5q!�m��;~V�;��/�ޤM��G8��#qv�3�<,KE�ȰC&����?Yu|?D�'#R�����Wq#�c!�� ��f��T�a0�W�0�$�)vf9�:ڕQ��6�� p�+���@�&7�5?O���H#Z��WGe��|���؅�lC�n^__ch3��1b�/�.!PEO�\�l�ͷ5��E+o��tf·�"6��P��|��5���3��}�:Z�>uͱ?�|s�:���|���E���)fg�<��W_�z�L���	��'�,�	Z�sף��.�`߻�#"ʈ��!���0�~.m�9�ß!y�c�^m����~Չ�xO�=Q�Z銨���r:瘍�
`4�ߥ�x��1z�����H�xT�l�V��w�k���ZO!akgf�A_է.՛\��'e�B�9^8��b�l:���U����M]�Bm�p��*����^�
e)�o�ȹo&�~
Wj�g�K�h��[�z����aP��Q�@m_��"͜��I�fi��w��	z��t\ ��#q�y��)��+"�x�V|*@�;��~	>�iY%�[%����ͩ�7�NՏ�k�3��hk�;U�5�%�5dv����N�b�737'���`U�wed�m�>��e�m��rs���ZT�'�v��n����Z�%�M���u����c���u��&�z�,�:6�.a��8�nاD�JL-e�uև���/¹+����̷�r��h�غ���C�j	=�Nt��]�ga�ں�v\�Y���.�骎C�GՂ��3q-����G%lI��S�
Y�4�ۧ;�&%�Ƣ\5�I�.���<З\�ڣ� D���ZO��� FD�iN#�"_5͘_�$u���(����0���\T�G�lX�+�p�/Ow�Yņ��s\��"��|�G�/���Y�"x*����j�>|���Ŏ�@�Ȃq��I� �W�o@�������+�~w�� �i�7�%7�A������"�]ވfM��\�>�3�Ưg����ZIz�J{�Rأ��g|�4�UQ!���Vz�2n0�)WT���������P����/�ƃN"�D*I�!���DX�����m%��eX��Z��� ͻ�ܓ%s�%�u��d�u����|��!��aј5�jF���}�E��H�U��^5���i��UY������%%�L����P������'�x��8�� Ɖ��ts���1}�'T�E���Y|���͌\#��I]ގS ����g����E��-�� [u��ۈVl ��}7NN��1|�'���,�}I4L$j�J�����>mM���ʋ�����B'�T�ah����`�$���_���^o4#/�g׀#�~�A"�n�~,1�2r}"`m��fŒ:|�
Zb9�>_85�+S(���#\��0퍝`�pVT��%�w��
��)H�H�w���ZT����Z�Ԣ�]���sV��yGϠ�������"cX�%�SEf<��ۈ�M���ܟ1���|}�]�B��Ƿ��>��}HKf�@�cNW�o����E�������#�ǆe�΄�*�b���^δ�% a费��:
=ܿ Vd�����(��h��H�qY��nYW�� ���L6��P�I���9q@~bs-!xm���*�e�Ͳ���~z�����7%�ۛ���o?�6��=�o5��2�0���O�>�|�� 2�b��1u���W��w�m~����LC�?���Q)+��r��|���\�f v�$����������>��֍9�6�v2#�?�sv�-�l�ڭ����`�7���|Id3I������z�kGߗ��]��7����G���Y��K8�#ސ� �@Q��y�	S#{p�O^>�!$��r��\<�I �U�������Q� ��T��1�r�̀���f��,,*)�	D��۷yVU^������C�
�� ���������ڹ���2}�c�����V��	y�W��k�&��4���j'�x��ဤ�r�m��">�; �-t.h���c�#G����; �*���Wb��ϊ*�c��?��#��G�u,/`>-H�1O:
�(�9��(E4,~e%�h��z���X��B��l���%�#,��+�Jņ�f���8�� ��ԩVV5��
ִ�V��p���_�2�\Q�ٸ��Q�=�򱺥z+ ����f:�)p�����|�eTUa6Lw�$�i�n�C$�Cww
�ҍ�HHw�R���Cá}��y�o����u����{f�k�����e��u��y�(��<��d�X��Np�[�E��T�d	����?��{����dƮR�q��S�\`@4�|m_��ל����=��6�S�'ϰ<S
-��h�<:2-�%�>��Yu��?Q�������qw�i���q��_ՙ�S1�j�e^���%Ӻѷ�D��9M.�P����}��ul��FX�\�����GGO�V��,̟|�HS�ϡ*�Z�2tL�<��'�}���_�����5T$��E����'��[n���i_�o��9�h��<�k�6�3<��6U�%5O<¨[V��s &�<�`/\
�i�b��� `��J�߆�K��$X����y�fo��7ƿ/���n6Zs4�3�6b���Z�Y�+6�Ǵ\�C겋���umC��0Ye
�镯9t���я�tg���k���|:��]]��JA�t�LYbf��n�����W�㓓h^y_�����BqN7�*7�0ާ7V�X���V��T0{:����a���	�D����dm�wc��%�7�U��їgU�	�
��p^�~<%b��7Kx�x��_'���{��U�)�X3M./��x]��ml��W~�՞�[e'<焾��e�dB|�|�����*1 &x<%$�]	)���|ݴ�AZN���t��)����?Z 5�����묢��8��0�DfX�!���kV	��SQN���A<3��"8��5L5�-1�|�b�^Hw�,e��3�l�c �q9'RNx'�
u���X����{Eϰ�J�a�h����.�ϔc��EVJ?uCGiIJܘ2���3Ѷs�ul���M���%����\�=B~U�� ��@V��B�wM� �P|ن�����&hy??�� e,Ff�.�u�<W�ܦ/OR:bY���xqY��3|�o���5��b��d��'��M�rmP�d��>M&@-Ԑ�I�G�|w����~p�YKpӄO,|g5��TA"A��y|y�!L���k�f<�.�͗y���gz�w�����n����.K
�j�n�9�kf�7r�Q$����C�O��φ<�(�3C!f0�헺L�2��R��}ۓ�o>�0˜d��֗H,�� ,��?!PYE5$�3������js�6�ߔ0v��~<��Ҵ/��r������i�1DU��T�Ř�#�zBB�F�o��gRBn������ƽJ�Ӛ>�'9��Fq�'�ѴC�˼���ׅ*�>�!����O�+2&Î'��<�ܤ(>{���r�V��,�q��"�>��Ņ��`[�D��7!���ϓ֬�F��/)�����l?��g�}N��v�K���]eP]��GP�q�~ܶ�I���M�X�c�6�Rŏ�(����Ē�����)q'�Ii��X��ؓh	��D��W���~�F{w���W2?䙂vĻ���z�Z�������V0�!��C��*�u���J����za3��}�����N\��&'�����*|6)��<i�V�2�"�bA�&�?8�� �BW���~lm�+�\6��o2��V���1�<����/�o~繯��|�+��,����R��g���h�	L�\7����8�s�?o7���|��� �+�`��JZ����.�Cm>��/���kI>�n�߳�7�������Dp4�/�^h٠�� .Aclhjv*u�K0N(A?�5��2�u����Ӝ��J�zfJ�vhZ���f�iZ��nyC}z�����^��Pf-�w����1���m��b0j�K��������t���v��{ގe��w�	7��4Ьȼ
߆�OOs����	���n���M5�@�=?3Y�ӭ�&������kc 8<r��*�(:����Bvp��*�
7��혉�4����ަ!oX�is�Q�\�ا���n� t.��Ǟ.����z2�u�V{�Q���X�i����M��=�����,GD����d��PB�f��s'/��v�crjj��l�P{��������w�U����2��NF�1��Y)L_t?�69[ȕ;�`aDQ��:��G�^�����S��U�ݣ�*��P��dY��G>9��}�����>X/O�����͛����Tv� =�7�}o$]廃���W�B��w7��Y��> �|�n ��f�{
���v���������8aݞ������z=��0���b[�\�W}�1��b��L���_�߳k����QҐ��n����sb���X� Ot�^59����#]�T���߮�k'�|.[�uF���]u|����Ng�����Q�̕�},Ƥ��>&�������e�#�>�E�3*�^�-.|����/��6h�������OK�_���K�':�8���p�nڨ����Q�z�(�h)����!g�$+1ƷL�o�5�rot/ ��'[-�S���2Ja��y�<���XW�V���^�x��҇��q$�d� �=j4�|��-��|h=����c�����kjhl;d����CS��g"��D�_�/G�4=���j/�X0�(G^r��]5<l��~I�#�P�ipEiL�����'Q����/
2LM�����%_��C��OG�4����+��B����TM����P����_�p�a��!5�>�N�W�⿖��4@�.�󫈛j����Sm��?N�GQ._~�kyĲ�����p9Sd��N��?�U>]g��	E�(��dJ6$,��ǫ���/�m	#*Ar2����r%^����B���Ɍ>U�>)�Nr��� p�L�N�{��lrɖ*�����2 @
��d�F�qu����'{(���Y{ZW[�rL zr���b��t����:�D�"����t/л ,s`�6�#&�+=
φ��D�'ïuy){��0}��, ��WP��@��?wn9y�?�#8���/4� $M���{�/歎���eH����?�)��7x�޽�o���g�	O���z���+��S���䁐q
D݇wE�0x��NBp�!E�Y�O�c�N}:�E1�g�$��m�1͸5�
ޤ�Y���7.��Wl��&����W���D����������z�5	�c�m��1g�c}zi~>�~��t���ѕ/��{���Vo�D�K+����',z}�v?o��,bwdќ�N�Y=x4ǮI�le�4�5�~�����C��֏���11����;�s~����"��|n��J�� ed%�Sâ$/yO9n=y~ZF�X\I�齗k+�4-2!W$�´�A�V�G*~5�,cY��ݙ���{�*ġX�~�+�����G��3D\�P3�����/�$_'��#"8��q��� �i��ܰ� �1</@�VMc��~T��g��jy����'���g;Pa���Y��%�Z >30<��i5�����!kK���MUt�<�
�]������9�h��}
נW�8��qҖＫr�:�#5�Xb����pV�U?5i�ʔ,��e��c�y?�����}�ȉz�רZ�'�2ؒ��?S�
�BZ��w��q�߮�-U�(F�+aӶ�E��5&�����|��l~�M�Ǫ�vz�<ն���&��3>��
"��������D��p�a,v����iA|999p=_�/�B�,��- Ɏz����k����O\�ݧ��(����&�t�C5�A��%9fb\ae�d�������-�R���r���ѥ<:O�V�u��N�z"��}�	�*��bλQ:�.�����`ko����u> �s��u[�[�׏l��wg�MM�x��O{���YV���ވ��SfYw�P.�
�v�w�)њ-�ּ�z� �X9f"�:� Gc6��N�T��Z�-S��b_֠Aj;v��h�?�bH�B)D�`f�u�p���M���PT�D:DM1�7>(�z@��kX9�76�wjD?o������ԧkP�HxJZ�zݫ�%|w��g(S��O������x�}
4��#,|��@�`F��h�YW6"����Q:_�ji�!�ó54��l��;[�e5�j]<...��#S<<<�}�"9b�.f�]�#D�������1����(�O���OY������ƯS��7麸�u�6��#������S��)���F���Q�Ϟ��U����&�L;�̼u�/:^㼱y���jX7 ��,�X}�m�}����$�;��jm�X�s�8�����ln��'nSv^V@����vӧ��l��;Z�B+%���R��z���rX��C�����7��%���,��x�>Z�Y����A�bWۗ���2j]������k��rzw'�޸������x�\=�d˧F�3�s[t�tg�q���9n�,q����D��:�����M�l�_W�#�:��<��ӴD霹P��`2�u||iyYE�n�sI��Q2����H�+���:�nc{P��~RB0�w�<2=;?��?�U@'��s�m ��'ͦ���XQB �MTj�y���<;�s=��k���Ч��sP���v��%/���)�.ki��-��>��r��WZx��
Q0N�����=��J���zF��hԞ�|��ۭ����^@�6����O��a.��Ŭ��c1���{0;u�e�,���5����$���	��䋋�T;��n�]&-�*	�L�����ځ-�j\Ѫu�*�� @^��_�:��P�����I�xv�>Z���Ug2�l�f����/��Vu2�[8)�ql5����8XX��s?֤Bcj9կ�6s߆e��|�_��;������[�BH�Ȅ���!���e;�~��O&ޚ�;Y��c�����/?��퀯���{���Ѹ"����t@@�¿l�~ߙ�����i�P�ceXJ��$>K� �,~v�T������\�Nt5�m,�0��f���q"z,��X�K��J�y@���`��!�J����Aw���6��tt��,�j�Ƈ�ŋ�r�[i���zE�EnRw��P�D��=�����!_I�d"��T���""�<#��WBN��=Q�eN��X���YX̴7�}�@�*li��FQ�#��7Z�o���#��W�-�u,�S����D
�<�g�no��`�.�2�5���{R�T�V�~��9 �Pf��3B�L�}zz��qjq��p�>auJ�=����w8^�6�!�+8o���K��(Q��ag}R��hk���c�`Ϟ`�^�� ��Q>$0�*�>���:1AQ�W�q}}�x2�/>6��������8yT��୭���,<||��Ck2zUY�[��<U,F�q	�導��Ƴ��lܰ�.���RX��Y��<��`y*�RV���%��}"�D�׺�|��R�b���qcXl�-���k�w�bqryMMT@�;�,4�9QX��D��/��}��t�@m���˼O��s���&TP.oL)�a�C�;��h,�~�6�Fu
���&�.�/�O)�����؍��$�D_��cK�`���4S+0��y��Uf��Q���h�l���$�҅rĽ��uR�w���|B���lu�;�^.{@�p;�:E�?���i��V�ߌx�U�1������I��1�j�!�)�]�3���YP���#I�j��eNV��7�#�h��Ԏ�|���5��h�t����$�(a�u��Ky����`_SK�ʊMTL��r������p��r��lи,�_����F����YX|��87UU��Xk�gՌ����Ja�f��|���סMKy�������aT<�V�T�L�̞2ΏB�?���[���{�%�w��S`"*7��Y<��J� ��ayy����6y��/�)�ttt������:M�A/H}��G�T�����aU�x�*!C��X����
~-��pՄ�V�20d+�@O�Q\�M���C=�A��D�&�H(�&r Q�˽C�|��NH��7Yx�I�F�D��k�v��ז4���IDŭP}ʲ7x���`w7;��K��S��H"��|x#���N����$p[�o������b]�"N[Q?���Ґa�z����"���Taʜ!H.�[~�6Z��P�c�>5��m��E�Vu�5r�8����C���9o�����t�p���,���Z�>|�Lk���T+N������ؾ{SW � W�Sq��7�`[���6��r����N#n�ԱAඬ�`��.V��ÚĮ��>��g ڃ2~��f�U��lB�iM~�(<~`�#���<Ԡ��+A�C�
�2~�st���f,r�a�=gDi||m�f�;(Ң;F�f�=�~�K�9|5ۼ�Fb��Q�(������3K*�X��&���[�%˟g���U��#�-Ǜ���.w�R[�W�H座&��===��n����Z���Q���;t|��Xi�9��/�䲍�h���~���w���>%e�:8�ޤ��"a���S�
�u��5���WGK{gUXD��%��/�=z�M	i9Vҙ���P	ƻ�\A�搰n�k�>3k�rhXߤ���������;�V�*	F�����<���iI�䪢"�Uf�[OmV�1��k+%��Ye8��ȅ,������g�T�Uϝ��\�ŕ���f�:-(�s��(y�jN|������O�UΛ�b�4E�RE��em���0�VnK��ػ�s��=��S�ӛp'A���Qt�㭨��jِĘ�����;��_F�j,���C��{���;����N��^���^��
|�w��x���V0b��A=Ekձ%c�L�b��`�%318�����@m����i�B�%{�ZZ'ڠ�����̟��6o�����UNN�%s�J�[Z2��.-UӚǡx�P,�.�}��_��S��wA�pX6N䠡 ��$�V�;����q#f�%��n}C����.��ض��u���g���w��bi�jo3 �c����I��("�/@��s������6�^ŭ��8�"/eo�g6>Aa�7 ��ir ۃJ@� �d��_2J^_��]\h��v5���9}�	�{+D8y0��v��+k��YO�8@׾�ӾJ4	�u�&�I1~{����-��s ��y�U��C��\��@�T�J����3Ȏ����^��yE���L ��lP;�8���{�i��18��Ih��\�_y����DC��`c�7��<�����[��@G�򖊜2= vZ�N{�4���E#>�O�#�va	�ܜ��]�Ki�=+c�/����w���ވ��G�'�7[��
�{C���t�/��E\@>Ń&{yw/��j|�W�xL���ϴ�e���ǨY�P[;����Q�Lu8��A�C��/�Z�E��y.�,]��ea����Y�2n���Z��хU��/�Cn+���'��8e��m�A��3�F����IB����y�6�x3`� �;8SHw#���Y��Ǌ��� ��ʢ��<b$�At��2�K�!� ��D��OȥNt aNP?_~��qj;���d���Ťn�V�ex�A�Ņm��S�����j�s[��橚�� � ��n��=Vs�ws��Ǚ���$Z�K\^�[w����R�K5w����˼;a�vc�3zS�8�룺r�wZ]Q�A	�	���Os�L����U�q5�3i�h5��Ldx����G�ֺN.5���+�����ݠ  Z�Ƕ�ܷ@��SaS��ٸ���O_5��x�@�(s̻z������43�Z9J���+y�u�rBڻv>�/8�VDx�Iz僜�i0�r4��l_�c��0���WTV6�u}�H�R̪�wĿ���9<�����W����,�`$��'RI���1}p[h�UǙD�lg52U�JdMud98�t�	}�DQť�����ag�6Y'�+���P��d=��\��&����w�jp�=8��ź*?`���:v������t~go3=������=#��4>�mI-g��ӓ������>"·Ԇb�X>]��z�O[ ��!�M�f�"�����'��KX�I��u%U�'?=������V�t����d�
��ހ�a�~�����(���\`��l����IC
m./��ס��3>>��}�~����x�?5�.��S��8߉��8D�J�]�[��0"����/j�P�֟�돊����W���Z�TXi��Hs�w´�N�_����;u	�	��LLL�������
a�AT�/??�*���B��
�w������_D)2[��]Bf��>h3�ե�r�Ԣ�E����V���um�Qψ�vS��U]��i�KC�y&�5�� qͫ��" '�q{��@��o?+�Y	����8����#�'٦�ǲ�4�ػ����^/����.����3l|1��@�!�~����n޲�� R$�f���?c�}R��5�;�Yis�8e�݄M--� X�ˠ����6�>6��5�P�?r���S�<����d��p���N��H�U�Wc+[{b�2��߯�(M�^�Ri:��3KL��R^4�H͒���(�~�9B�aI(p�����wz�!w����4������ [!s��m�_$5M��Ѭ � }��QIĞ(|����g� ��|�p3yp��w������Ҭ�,#�E�dZo3A�ë'��e�֭�������lX姹d*�b�/�ܧ%ˁ=z�����;"I,b���*�����P�{�!��8��b���@���ǲ��w-��6%']�b�(#b�=�V���C0�����w�o6~kѭl��O���k����v��WVj����bU��Ѓ���q&� M�Ծq,,e���.�'��$+��6��CT\�¤�V��l�
m����Րq~[��6%�X~�I���d�/�hx�"�Z�t��{�y�2I����@Mw��J6A��'�����j��Z��p�)��)"��KF�[���;R$���X���ς��*U �&2���8�{��C�ZZ2RY��/߼���9=}lf2�)�r��tn���=G?�^�G������א�8K�2}�Zf��ld���X����"�2������S��wD��ˇ���T��k8�3�����cV�(����y{<p��s8Kj'E�p�e��G���7ԒW�TQ������<!b;���Ō�˩w8J���xv�g�Ծ}���?_L��;��Z��8I�;�bxz�ȥ���I	��	�(���k�)>^X
��6?������蜌jS�Z@��U��@3�!iN8$*��o��-+��\{�p�c�V���y��ț�6c�w�qO�^M��%���r� 1D�J��&3���^��i%<�:~,���"�.M�>�A䲬�|
�>~ȏh���7и3��jҼ�Q��|ںrm�!X�Tӹ�[qY���!�߽�� ��n!m�� ��ht>�'%�F�L������	�����:F������WxŪ*�N�+��D�e��VNn��WD?��M��ʪ��J,�W8v�=��ܓ�2��u��]��>`���6"F�&��l�=�xd�A3.���˚Q\$xd�
F��8x�__���}%L���H����Y�2�f�tq��J��GO(�/��L�$/'��ʞ��z{��v���z2=��wY0��)m�)�P�X����D
��.��?+�b$��~��������p���������K�ȭ��b��#�kh��[w3Z~��-i�-��V��{G&�4C�۱J���j{�*�NE��j_��2�t�V�XT����_���|n4��۞ڼ���Ӆ�w���@
T%e�@8��]��*(�Z��e�yYM��)`��I�r�8����Z��JX%�9���DGl�y짬��[������ʹ}���H-�m����ɷis��{܋�}�U%���}d@e�9��۱��XZ1��2�;���0�og�ķ2E"F��Ix}-�T����F���޳`3�B�֓WM�(�~������m�5}'����_�߱wO0qʓa5�	�nps��枞ׯ^�yq	{�X�|~	�U���J�h��V�f[���sa���w��y����]/���Oe���P3^(n�Ɍ��/�6�`�u����&X��g���)	���`�'�!����v��IMg�$����	�5����O-l�R��U��1��f>�Q�w������V��f���`)���`�&�����v�#�q
����Y1��,z}W�I�.�m�Ky���?l���*2 V�֣Lx#s���@��~5�v�W)DFG�GH��H�_y��L��ޟ�kq�=��p��[[Г��>Z	>�;<`��d��"e��|V,�y�B!Xې!�Q���>l�}ơ����,�l�uܟW��2��� �"��E&ZSb�/�o��V�9}%�Q���S�����Lq�����t�@��1/L�:D,� eߵ��|���YZ��f���|�_��9�����;7���zn�~5jN�0_'�b
5K����i����T{�0b�o��v��@�*TB�,�1��2:��=��hɯ_�x��5��(I��zg	�?�ZS��l�4�j��Z�ɗ��[����d�1�8)f���7��?�R�r>��=ف��3)���������\��W��`���Ad������w��/��w]�/:���għݼu�B{��w6c��Hr���>�*����}��$s�ٗ"��{ϣ�4��@��lFF(�k�Y�D��u�s�\v��fZBl�Sm�wpA=Ϸ���l�g�hOо!��Q������)�����I���*H�������D�i��]�!�хO心��F��p
i�� a�D�W,B����P����2��Q���R��Q�~d~{�e�R�Я�'�ML1���-��z����؝4E�D���(T@J�<v��<f��#��{�kr�mK�e���&��%�4�w�%�"���	�F��M"r�T�gxʸ�?|ѣ�3���Z9���a��.�b�U\��������~J.� 9*g�y��q6��K����U��2��&�G���9biho�����?%���!^Aˇ����^����lu�4�YO`�����O��
x��������ۮ�:󛗟�2�ajR9�ͳ���%�
��SL�������Ir��k"Yc��\���`6~����κ�U	�,4�ʆ�c���s����d_���M��|�����X��/�J���բD�y�7���۸ﴩ���أ�Lux��������x�2��l�j{^������(<��R�@M{�a�QR�/z����l~�|�6�����>D�	Nb@JO��r�ui����S��Ə�P������<�&��oL0���I0}���>{�U���K��31�_@�3ʓ�v��-I�%�#6+���&�U��j���a��/��\�*���J����m��\t��T&��㏱pL�vrc;�Y;���#�c�2Sm���o ض�K�����a���"v`=�=p�7���� 8+~~�z=��V�А�a63P�yM�sq(��ny�Z�����=;i��[�?�����Q���h3����q���Y���y��$l�֔��_��L�.�D��M� 15�ڽ���bd�ǿI(�^�#�����\u�e]9xr�0j�3��LG�Qb^�
ݤ�dt�ʞ=(������&O@�==�߳�`e��?u�mߛ��~�iCL�}A݆!��҂�Q��	*$êߵ_LX��4��6r���Ծj�����H��o
�խ��6! �*#� �N�5%WM ��	�
���_w�/ہ���f.'G��|ZBhj���������P��x����{�ygۤY��{�G��he��Pr�^�	AKK�q/�*x��I��^++㶟f���H�;�Z��f笭���_���Q6�����3D�'�8�KR��X�4ʛy�CNi�wEE	�(�x��>ʅW�����t� ]q�]�JR�ۺ�"��qk���-���f�<�dg�j���?����4˗�R�n�?UA}{W�p����(��o�����?��F|+`DRs~�o�X���;=��k��+�?M|a�DGVf$^�\�`�=��0,�%l wQ��b���Qr��-[h,�!�����������-I9@~�­<'��\��xț��ar������"��G`[�W~)GzFF�� �/��qO�^L���_bk��&�
�������H�Fx_��]�i��9	��}ۯ9�c�c�pK��@={�8��K����~��v��qƼ�ֺ�Ož���-|Q�a��~qʭ�6������df~�A��^��mR�rQOՙs���'��x�<�!�f��ID��<]ӯ����tB��nq��Ч88��i���S��$ �2SR(Q�6s�p��u� ���Đ���S����yp;hI��ܩ!��X�U\p�ξb��og����c��l����1�J�8���W�Y�@�Λ������/ځ�Y�b���VdBz��h�,�HX
�B�/����QY��+�=��t�K��tUܟ��&^i�ݣ�j�.{�T��b7�	�}����O���N-,v�z^��u���u6���:z�ôs�����A&�ǆw�%�YIqV��=.0���(�� g��|�����a��foCO
=X2C�5ɚ�2�YP����(�Vh�/��$���!�!G+�1@(C���9oX�n��:ID)Iæ���X�D=�m|\�����s0�2|Z�� w���J�p�a����� �(:..._�k���̓�j�]e���W��Nt�t�p�P��?�����Bi�S^�0�Fr�d�y<p���a���Zn�X�*,J�����ʕ�T��?�O���y��1��+Iw�j�ņ���?��>�եd����WUou|�ۓ?��p����)�!�l��1N��o�\��)1�m�M=�±���ò�4�����Gp�\�@a
�i-��|���PxӨ�c˴x�O���-�-�7�^=5%~.���	/�QW�M}���	i	�����ZD�缆
-e%�C�m2C�ƺ���6]
�<_�J��ň��oU��@�b ����ye�G#/����mP���E:bø��L��S�x�1�e��is2A�s�U���C�@	j�vɺ�xu ��1T�E�E�5�����$����$(5A�؅����������������p5M����,ȏ۪^8��h:q�:Y��&� ����b*�{��Sw��xCju�xC� 8�N�=����SO��������1p�S���,��G��6~J��V�k>m���&9���ZTbF�2�2�V%miQ䖼����Z	}�x4i-�����I���8W�3�&���U��z$Qh�7�����TY��n�Q�"��<��Yl�A��G��M�l��_m
o~� ��&������<�4�����	U[]�G�_$g|E\���EܚF����*6c#%�)o~��f��a���l�7Aԋ҆������r������̗�@�=�Ç>qj�+I���M1YK���W#ÉG��
��m�&k,�9n�9����5��v��X��"R^hԷ�v|y)���:�>+�R����A��=��������y���z���J�y.�����0Q~$�s�����>L�F/`�!���l�E2���ѺJ�JEӌ�Cǩe�����D��$8:�����͘]Kz0~�)��Ŭ��?�����u=��CW2�ه��G7���Gϰ6�/�o>��]��j��%��j5��F�M����]�.��$�u֠��c�����K����j�7�2#'٢���LIK?��g���.��@�ՒZ���c�5�G�HV�J't��ilF4i��� �5�����S^B'�D��/Bìv����'� ,���m&��m�C7�9mgy�X �S�Qh�p|���v���쬫G-���X5Ҝ�5G���$��2���D�l����}���)$�Ȳ�Y�\;�(�p:��(�I�zx�;d���<N>ȋ�j\}�_<}�z����kQl�8e{eu���!��5�$�׻E�9A�D�����j�^λ$��O-�t�܅<x��˜y�~���R��[\c#��abܧ���+42���J��/$��f��<P4�e���\�8ON?j��S�3*����5׳���z�˲�kNpCQCC�Wlu�@�/Er�U�p�l�lAf��SEd�o��f�q}<����H&ِ�Y�6��~i����mg����	-:_w})I���dH1i|].>'��h�L~<�x�J��� ��UBv�.���z�1J��q��]t4N��q����v��'�q�ol<�Ȕ�@�v����^s�<Ӫ�KM��-��2@t���[8/n���H`鄑8j%�З����(��]��P̖d��ِ$1��U3[M�"���<�R�"Dr��}��I�u��]:���\1��%���1���sP�Z���� -ʘ�Hw_̼�tZ��|�Wj57� ������ ��M5%�BP��s�M+��&΀�)����V�S���=��a�R�{`i)�ŝ��-:^O'�u��?�[WGfhh�4(�ؘ�4�ǣ1��{�e��W�Ѵ�&c�Ke�i�D��'���Wa?��_�(`9IczȾ�V��1)�L\�B!���*snQ��>h��a�]cJRkE�Pي�D?�˦�ٙ�VQ��>=L��7�W[���9���!6Wz���'�Z�wM(�j�7s�MٕRY0��6|:9p�Y|��O%?n���Jg���i>��<���zB/Y��J%�,�缁;r�9�y%[=;��~���῍:��5���I�|����A@��p�����AnP�<�R5(���͓�G��.\S�y�H�f@�����L9I��8;94�$��ˁ�Vz|y��r������v�	��=�L?�cυ� �Fi˨���^x34j^@�o��!�G�j�	E��Ȣ,��*VV�N��z���q9'�(DL*��v'X�CJ�T��G��SW���Ō���U���+6Y����[7K��>���k�iT� S��t{9\�����^�r��r�0"Q�!����ͧ�$l.��3�E��k���	/t�2��"���a���d�`z����mL��(�{gW��~�l$����>Zխs�U,���(�5MQ��g��wy�q�E)������F��Mt��U��|����I\پE
�	L����N�zB�{��n������C�c�M.;����/S;;<p��1)|6<��%:py48F961�FL�~]8j3��փqW˪`�|NTggKv�T�2^=�8=����������Z���i%$�c���G��v=�zihq	;�k� hs��ݚWE�S��5����\?>v�q�҆�����J�*��(�"��������C��3u���|���!�/)�5�q	��[��VJwf�s1�1�,��d~��Y
پI`��2�_M�Z7���!7m��V;��%�F�m/�G�0{����L[��@���{��;ѕ�3��̵+7����vA'8��'ײ��>����4�� }V�RC"gjH%~��[c!�nX�xρ���q��B�3�n����̺�ϐ
��;�n�i�1�E\�����I�ͧ֑��@l��^��	����L�I��88�[V��l�r�]�BZ�.�*C�h��gK�6Yn��,:���O��=���l��\<F5�)�=�g� s�����3:8}6O=���N��?&՗�����*,Ϳ�lӪ&��I�Ƽ!��|ꑒ�W���I�*J94OS���.d�R�5m��{Lo�;�h��X�,#)M*i�i��F�頛A�F������Xl},ON��l⭁��Ėo�z�a,0�1��/m\�����<]��6i���.���}��d��.F�&팸:�\���*	J<�-��7��D}�R���$)�A6�FM���u%����Ew��.��+��eO�:�&�V�OjQ���=O~���9n�Y1A�x�R��/2�l���ُJ�Fڝ���$Ɲ�;��;�g���A!���q.
E=�A\Ҕ��(�mp������٘�m嚻���4�_ȥf�/F�jx+�����\�졿�nа�����6���C�#�<���v�ZX��ɯ���U���l����D#�g����i`I[f^ףl�=%�Ɍ2a�_k%�ӫc��ݬ�mY܅'=����߼T)ר�0���9�yg�����%/9����%d��*���7�no��/jrVA}4������V�e;lHu�����1L%z���$��E%ߝ,5�bU��[�T ����c�~%���-c�c=Q"��8):��ğ?u3��AA�f���⦿Y��9��Z�Nt��5�|��8/��
CJJJ�'�7$Ǯ��E?��ywV0�e1I;+�I	��V�^����{�5<���Qy���a�=�Fd/��o��Vv���|�1��xo𔺯P��Q���L����y+D]^��-��^��S���V��k�:̅��ւ���l�`{k�h"�T��@> @�UP�XW����G{:���#�3WG�Y���{p8O��K��?�+�W�R5̻��;�X��-�X��_���Z�i*���ݝ����jqn%���	('.��M��2���FC��FÐ�u.���rt9��ye"W�:p�
�UP��~w��Ck����VB
_Ϧ߅�
?�B�m�eQ�0R4���r�,_���@2��S����}G5\לM�1>F����6����X��6ʁ��V�w'�M���z_�n���i7������n���Sb�����n�Ut�jX��1F;���b�����|��n��]�s���&�)U��piƬ�����YB����k~�����<υ"�L�����ԇc:�}#-�d6ߴ����fv�h���ܹ�Ff�P�HǑy�v=��S���h[��3uR*-�����i�J��5r�J�}D'�	���d/u/�j����(��v���3dد�ã��˓�[�*u'^���2,���A@J����	����$��n��e���A������������.x�㬵�>k��z~��yI	��C�iD�RY$�bu��ܜ/"�/����Z��e�o�қ�lM>l^i�,�ޫI>�ն�+�ǭ�����������6�j��o<=?����\���dp^��쑖Ο��]]�0���T�z"D���|pP�����5�^��{w㔜�6�@��8_T��
�����=<��p�f/����u��;�U�Cv�l��\3:cxؘ&�B�;��͑��������na9ws�qG���J��bٛ�e��n�0/�(�dqG��H�`iǐK�n�����p��Y�I�L�XV�2�}�0x�Nm<�.rx�O;G��;�j�!"!�k+�~݂�0��xU"Y�E3�kx��81���ȃɹ,"
m톶B�1���C��s]�j�|,dh([��<�:�7QV�CQ�k��+g�$O'�.*jy�]�1�t�1	�_x��߇p��y5�[�Հ{G��z���|7�oC���!�4����C�H,�a�kļ�V��3[*��J��~��3a&�����7s3��
w���җf[�!��YL��kD����ܛW����i)�!0�r��is\pMNE���gjP�ýV�7�}�U�|�]��j��&�m�˰`��u�X�ڱ�G>Rz+�Fc'8ϊ�:s+ۛ<�8p�9A��ڛ(���Af��畾CeY�zw� 0F^�4|�N�{�y�T*qlr�%{�V�q)�:�(=����yzg�F�G��kJ�P��K�>�v�4Xd��e`}6X�Ou�7��g���7�VĄ�����&=�7�����K����<!�'5�a��¤���o ,]�����C���3s#���7�{i*���� b���[b���o���hW��PZ��_G\#&�̺��_�/���mh�6�k�}�	�7g���`x!Т2�Hj��!��൤��m��+^O ��E��$�y@@@���F��y�ݟ�rQ>�hiko��Nԉ"��<�����R������0[�;0t:�����ygR�,��W)J�rka�?�lq���+��������T��"9����o���xB��j�sG����ׇWs��U�4���HJ&��E���:�E����w3�#�c�YK-d9j1�S|��[g�J�w�֏�t��!S&�.H{5�'(�"�r=��D���!��4po���͇�=�]�q��13�aA\��.�;�����>�'�e�k뙧�� ��uE['���7
B�X�"Ja�3�1b�pfWB�p��p����Aw��rS�k"�˽�$��r��;^�Bu�2��h��f�D��ui��~��C�B�YI�i��@
# /Evx��Z߰WlӪ��=X&|���d |4���9�$U���W�Zi�����I��y|� ����pv��,�0h8�n�.��n<d)ȿ�����yJ@J�)Db��lw����o{˪tX�8\|��C������4A\c�����Dm%H�Û��%�y�*�<ǌ�<*`�K&�~��y���L���Q���j�����|*iG�<��H��E"%8�����C���	�	��G[y�V��C�����,P����4�O#~C^�(�7��h�q���Z���a�I�)�(������c����ɼ�ɨ��-�W��pW����ڊ�_g��2r���|�� �*[�����7f�c��Y2��e����If�c���T�-�;
ƛf{2���/��2�-���yuY<,�Y՘�1B�3,��y+`�	�e������;/�xx�N3ws���h��B�,i��c�\�;;�&! ᇱ{�GS����[�j|u�Gǚk�};�ܦ�<O�
�F���=vRh�)��M��ᱚX�kҟc��PжR�CKn�2θ/�Q@#}n��23�[�G���A��68��b��L_����Ӫ��d-5�A�2�	�Tϵ߿��ՖK>V~LđQJ����<9�*{�^��|_]UQQ�%�� �0���Y��'{)������Op:�����<�����ú��y±��)�W;��Î_#Tn�:Z��t�
Uh�I��"+������j��$LZ���\j��� ����	��?Ə�9�kMn_�P�+k�^<�r,M�]�_@PoB��qR�DA�b<�`*Lb&|?00�<H�^?H����k���h�:\9�k�e�����z����p���M�Q�����v�ͥ����Oz�K�ٺ��m�׆o� c�$�AdS'��qӰ�&��X:,�o�A�IfM�F�-������%�,�S�!�`����0T�T�Y��D(���'�!��S��ي�)y+�gA��ݖ����hH!�ċ����Ra��h����$P�?C~���Z	DX)w" %��N�*��H<3n�A��11nƑ��k9��[P0��$Μ����#I�]vHcӳ��a�����X���E���<����9 K�U��I���r!ޔH��n�4�+S@��7^?�q� �6L����3��p��ǌ�q��aG���F=a�r߲��2]ei�ql�1s�	����v�>��"���s#� � �,�YYs���������dU"�Wo[���WRq�L%$n�6��xt2��$%#no�`N�yq�!<�Z&z�6A,���jc���
�%��+crAf��V'�͢^j<�e=��_���P�Ǵ�B:���d���?��o"1�/q��q��ҹb��kJ���{$V��ͫ(z����'O�J�M�[��*'4Ī�� ��� Q�BlT�i�5���Ս4C���+��a�>�k�"���S�P��ZւQ�j���Q��y{"�����w	�B���n������SOS�(SJXE?��iy3r3���3�a8���?NQ(�ԝ(�YW���������"x㹡�Y��G;[�F�y�~$Q�4�5[<��^����'�������ٽ��S���x�S�����K}���X�����܁�N�;\��:��a�#����<-M��,�E�^���^��Z0T�����= ��ZZ�����֘rYE�cȨ����&������@4����������;� �p]���oL�6�8�q4�414"��\y�<6k��yjzm���Jy�~6��C[��B��~�8����ʸ���{�:o$�1~��k���®�D2�����!jV)��Z;�KNX��Vȼ��x+��V�)���� ���,� >���뵄�����(!�� |��u���%��?����^��¸�6��P �ڋ)4Ԭ������)zªG>JL�SR{\{V�2+�~,)9�65��{��W �lEUU��"Τ�椮wt���H���Ep�cZ����z���f�o�+�O�9�\+�ΎEI}�>O�'�e*�ij��Q�P��Km�� KZf'5�ہ�'���π�/z]-�4R`	m��뛟e�b>�'��a��|$�u{�X/m��,A>�z>���f�<ޟ|���{;tN� 	����Jf�ۤ��UV�,�窫���<� �NkV��I �5�E��,Ņ����x*YR�2`vG�����me��k���0��~ٛ����-�S�f7K:5o��[�:��>8���p#K��\���~k�L��\w�1��
�����4��$�|q��D�S��2���m�o�TaNE%k��]�eҀc+�o/*�]#sSѣ��tF�WO��<�&��b�>�av}���<��R��E�T����q4b�;<P�ԉY���97K]p�e�o�_s-T�c	�}��%��b��8����,j����z\�?<�?�����y ���sv�"�b���;�8���;5Z���a�w*�f0���"#/��8
�A�'�
	�{���4
�������-:��I���d�(��M�]�ɦ]h�Q��-S8~u�(���ʓ��Y[����Z�L�"o���I��w���ʾ.`ބ_c�>Q���L6��!�c�B��+��3Ǳe�d��w�4��Z�Z?'�3[�Ωab�j�zQ˄��d����>�gK�43ߥ�~n����d��OLrk�(��ȫ��I��ׇ�?�"������y��x	�;��۵tXt���f���$<�D$|��s(�f����v�roez���)z���Sv^�败�ʗpv��=���+�%��ǭ�h�KLu��c������� Gw���YB��|*
��N�ҍ������q˻�S�M��n�dٜ;0�P���;�:o��9��<��*�Zy�:<��?�1����H�Y����mM'w�����2R�D{�u#����\������B��n�w)�zY�/bu�3_�Uy79'�{ﶪ���Rc���������[Φ8rb�$���'W�~����P��q.*R�����c�ڳ�G����Z��2h#Y�����=��T+�Õ(=a��kzrA#	\�@!�z�[|�^�60��~��a�f�"hL��R��o�����>VTT(f�	�J�m�B��yr�/�\w���i���G c��nC׈���ν�M���B{��X��ޯM}j\2S����ٿ��_�kcd�:��g��ml���S����T���qS*G�v*Q�j���]�q��uY�;u A? �O6kDA�j��ﾉ�d���q�A7�<�ڜ�Ja�����V�i�Y�Z�:�]��+�S:��Ӊ5U��S�B��q[l�Ta~���B�S��_�n����|��5cK����j ���f/  �5���3ı��;W��ؘF攽��_������YX�d��"�˸.g^��n����ŋ�{����{F����xi|�Ъ��m79ظbXo��V#W�����1^�=x�ΰ�N���O?uu�C �2&-��1�i�c�c��Ăoo7����!UUU�Qr~-�_)9����s|�"zᣅ�
f~g1&r\D��_��ߥ�w���GC�'02�iǽ�^��K�ra��Ҏ7+q"W}�m*�@D_DF`_�S �si�J��R%���Ɖ}�,��e��u�n^�G/�åN��d7Oם	r4�tq�}�j�M��­�0��-�I�����7lQ5�u���D��lGD��2�p_�0r�Kԯ�+��f�Q�e9�v�-œ	m�6��B�����/��q����ty�\d�Qo���D�r���s�$��ڔ��@���6	~������Oh�Wh4�(��0С��}'31L�깋�����[3�,ֽ׷�O��Sb��
�m-��B���O�||����g�2tL0b&j������f:ݲ�۲�o������o�"G?
ƅ_T� �_^!�P�h���S���>������ήO�Ϩܡ!.\�2|�+��(�����46�k�⦻���l�vG�VF��0ț��gu1�^��0%BR��W<ؿ6�ݢ!��OM��L���J�)΀�.V���������A�'�� 9� ʇu��!��\Z�Z�'N�.�$p�遧��Mmq��}��U��"��i�֜_2�6�ܓ�x�,���C��?���U���������V��Y�2�K<��NM ?���.\g���7��R�Q��v��h��呭���Z$ֿ����un��[W���@��T�q�|���-��=k)�C*�|���")�G��Y���9�3n��z�$x���D�o�\�]e��fQ\L�g.�}���(�������k6A��R�ǝ� ��ϭ�$���hVu�&��V�#�	��A=yh��`�C�/а�����o&��-�!��b2�Ȱd�x�.!hJ���o�ı~���nL�hg����sQ���O�k)�j���>\�b�lki
+K�٫~L/��2T���=��Ǘ2����ug�Х��6-q�� go^��A��@/����q�9�2_���f�Ӳ�� �ji��u��v3�=���J���Np�����-c6�K3�_t����R��-�c�����7FU���Eh��K:��G4זS,F����DE:�a�3a�#74��}�b&qR�N82�š ����?D�wR�&g��-;;C���p�e�h�2vgg�V�"l�>Ss���s�S�r�y�K� ��:B�����R�ps�Z������!��_ݽQmQ*����u�����Qoc�J�e"�(k�d%���r�����Z[[3x�������r4쮞��D��S���I<[�e�d�1���������SD1l�LΌ}�
�|c�d��˗��Zz����	?�r�<׸�/o^��c�r�F���f@`�Bg�$*�[>#e{�,��"��U��Q�#�5��"�5Z@˓ �`�k㘽%�NБą�cS��N��[��4��|����>X\{7�D;%��8W4?������/���B@�psC�A}��7�������"�N����_I"x�yP�>��!1�������ڻ}JN�؟�ڐo:S#�u<�ӈ�h�ϵvv;�L}�Bծ�66B���k�4P$~�E+zM����9�2�f���pX�CW���V���q�����gX�����NEnw����90^��1�2P-�x����Q�8H��ژ):������bǉ��;sw�^"a��ʨ�Xm���-ʳ~� �GB���.���d/�)|��I��w�}h�gr�g�KF��;��=��t�v��ţ4�W����DI�B��,jN��B��Y��Lmv���kd�=�W��T<C"���/���@�# -�y8���1su���t7R�8�+�����{W������,�,��H'�:ﷻ��w.\��m%�a�T����g��n��1{�f�{I��v�7�^���}^�z|*& �t$����hko�;����bἎ�����Z^�c�,������f�'��� �*�7,�d��)�!��$�@b�j�hp��L{�#Xkldw3���$�..^W�C��L��e�S4�h���	�����{�>4�gS|�SN�M�{W�ۯ�[z,�[��8M�a���>���2�si��F��.v���T�5����$V�k��a�G�=[���͍��B���V����V!G�W�؛��e�a|�!�X6!l�����}�"���!�hgWU�M��L�-:��F���>�0���t�2��~ReEA��|��C�w������:��!+�qރ]6Q���Jn-:�2:�1��xa����5xm�R�R���_�/ϕ����St��W.��G���֭r�_�quD��u���`)/�A�����ۘa)�I���������i<��q���
��e>i��rvs]�P񥺷L���(�:����3��B.�������T��ܒ�	������0�����`�~�˼�S4dG�5�!��f�b�{��ƈi�r�?B�ܳ��6_����4�{r��;,.r�sw�I�K=OѦCb��E$(�&�GT�Æ+n!�dF%'�ߋ6�L�<���gӬ�ޟPUR����򰯷^�G��I��1�<���a�X��>$g����rww�o'����SV��½nlM�~I��_�5*&��9m'�{��C��|~#I4V�'P|�J�G�'Bū*�&'��͞�ݱ�,����%��G--�Uv��PL�~B���a%�&�� �,A �h�EԷ���h_g�MKT�ط�:������`)����Q��l�b�k��HdT�+1@|��~��"��c�}(�S5�����ڷ��>�n�\�7�� �HI�G��{���ú�SJ�'u���gJ�.а�����VZs�Ke�)�/�S�x�_�s�ׯ�~��c�pcL�ٺ�\�:���!��%�ʋQ�@ޯ(+�����V�<�����V���f#����귡Ǹ�l�nlX�l��lᴗ�Ƿ��BB�����{"X_��X�T/'����Q��DW) �O@��H�4�^�0`�h 
�^Gou�P�6�߾�@�9f�[ў��(Híp�&���xt2�b�>Nrņ�`�������m�k+"`h:�g��{����)^��w���w:
^B��?�0�M��K��0M���r����z#�)���ڢ
�z����c7@*a(�� ��K�A!Jȴ��x�W��w��M�}�ABѻKP�C�r�������*�{���5Ӂ�J������ی���"V��;?6^^.�$��;vgz��X�/I ƣ� ����Ԑ�f��q7|�|jRy.P��}[�{/r���(�p�];�ܓ6$�	q"gK3,<T�0����7�;0m�u��_�
�ȇ/",����N�l0�0:k����;q\Ee;��1cotɩ�L'���[��.I�8o��j�݀���#��� �h��i��@-���y�>K�}g�D}��Yʟ>\LZ��"��/�;T��ϊ.ERC��&r�M�-Z����O\���uAc�c��:�U�fNО �jɔ�W�P�~7��������++� {��gS�ѥ��s'S�hX7q�s�ѷc6D߲��(�뭇��A�Q`*�Ok^����.�����!O��2b����<�)��U��X��#����|��|��e�@k�C���ڏW�C��X�/���ΎM����`f'BB{{�Gg��]at��qk�.؉}��~pX��q�s��B�] M&��Zo��;B�[0�Z�\;�nDo�#���E4��T�Z!� zS5� (W����ݽ1�{s�
p������_���yQ���;�1Ҫ�fqM��3|��+y��c�fs������NMc&;On��_	B>��sc7�T�VJ/�5����zD��f[yw/I�����9dd}S]/1^�t��8������g��6?�1���8�b�?�2�Fp�l�V�$*JI?��SW>�@ݶ1^��~O���q~c�Px ��ʲR&HT�GN����vbS�8~�^��qBH�qr3Il�B(��"���޲��u�w#���mO�E�P��� �å)P ����׃�?VgR/�j����d��`�/����Fr.cC�3�d�V��~��}���/�8��=P��g�qQ��k`f���<�Fw�1@.������m���  �<��'y;#��k��.�L�����U̵�UضC�t�v�_/�j�XTG+�c���^4���ͮ8-��o�� ��ST�y7(i��̇r!�R ;A@�E$���w��W[)��^����9�f��Þc�,,~�߬G)�>h�yO����A���-+��D	ģC9�l�9��!���/�V�I�vq⦩��$ߥ_�ŕ�fT�-�R֔iJJ���M-lP�@�AF�M/IU�[/����ҡ����M4x�\U�x:_�&c��6�+	���VX-��<�厅A�����ֳm|&L}4h���0����ȿ�7@����.�~�0z��ɸ�-��}�#��S�k!D���U�A�G�^��$D{_���W���<Xm�=d_����YsYQHdx����v�&�<���1mX3�=r�'ԍ�������@��@�=,O�����`��l��&[��7��\�����+�����M��X��k������W#���ND�{��O��P����7&DO���p9�������M�"���$Cy�o�m�Rubw*�f����O�Rn����z�nY�-���&w9�A�3�r��_�<�gf��Ty�"�=n!�N�Q=��d�:2�����5[��9I���Z�&����h� į6�s�M�:`!v��� ��{Yr|v�#'�pq}�E
7��3�z��tE���^x	�L2�~�,���k��Z3Q�(�����->�,[�0���,��Ib�׭jq��yvb�,��
�rkX�r�x#���z���e�jKɉ��l>)Qd$��~�]�rp�	dd}�s4d#�Oe��`)A�@'��t��B%K��d��������,N���e����%��ϴ�O3(�~��Bm��ײ[������ʏ���5Y�x�J��=�9<��sk�h�9�)Sx5�7{�C�9�]�ő 'NS��O.�g�/Ц~F��i�2��%���Upv^C� ;���a�k�
��6C[����}���od^|=��m)_-G�[���ԍ��Y��� �7~Y�vNտ�mՀ��X���cW����
�L���Y����FR1���b��b�q+C�?k>�$q�������4��si�E'��g�t�q�:*��8/��vYEMU_ki]a19��6�JW�b0:���b��w�S����;�!٪�9�ا�$C��Y��1P��L
�� �fd�VI��7^!�t`pc���!�jf*������WjOS�7��|7���ķu��2�� }����qMg% 9���4BZ�
������+~SD������k51D�4��W���&Uo�Z�K�;U��4�^_�C��=%I�]���9��5�OO �N�X�A����y�y�[�=�B��E�'�|5���J����O�u
uN��l]\��Y�p�܆�~)�W���C����;g�?�d����Ӥ��o�1�����qۏM��ͣ!�mϵ?ݢ�c�e���յ
HT"��*�B���Q���FJ-�ӵ1�N��#��� fc�?�(�9��ΐ��2Z� �,αςxˍ���2̽E�|�0 ��D��`�1j�Z�y���Į���=O`�seU��ҫ�:`�O�^SZP� ��Ce~�W쵹��`���M�����M���\o	^�'u��#M��p��ó�%�?��W���3^�SL��~���Ϋza$�d��zv�ʪ�X��^g�*/��$� kv�#s��"{����Jѻ���I�Wº1�3�d����x�U�w��*.|��Bճ�����	��e�7"��G��q��wK��b^�y�g�1^9r3r�?����QϿ7���N���R��Ԕh(2w�\+�Μ�l>�OI��a�wY�?U�;�R4ZΝw����ү�;����^w~��j����ZS!5�;�k���Ǣ���&.�6�P6�+�
|���:ZY�w��&��zج����MT�mrn��Y����?7M����E�M�/��~K"~X��8�"mx������k*g��~�~+�����^*m�#��,�pc3x�抓?��\��(KC:2L�\�"ٗ�&	�x��_��'�5�͈�_�ըB�㊘l�W�wg�BܰI(����Z���t�;��I��~�W.�Jb r`���JQ��H��^#�����A�ǻ����%\�'ܾ�,��b�6U.��uD�ǝ�g,!�G:ӓ�/���.��se/11Zǃ�1Tw�F~uPy:��H��9�;m�{#�����w��cc���(�je9�����Ɋ(�~{bh��1�3,1�(�N��d�JV�#伎;��i��@�
��M��c�`9���8�ٌ�*�.m�}���I��*��P�~��q2gex����l���������C�\�!��x� Xp�� E�Sp����q�����Z9���&�hW�_7�.&.���`揁��&�/%,^|��"���Ûw8��!�Dԭ�Ж��Ϣ �f��:��w��/�Y�
0��>�%���@�F�W��|w0Sto��bd����U�Qb�������N���F{B�����4D�6�"�੶�ٓ�"�W�Z�m���b�޸�v挿��w�����E9@�n��9�͔�A[8
r��&��fdl��I�Z��Z�5�Z��jj��*{�ε��am�^��H<*�Ύ[-NT�F}]U#;���2� C����(�]�z�@�W�[��MPT$�9��1��
s��1�i����?���w�� �J^��Օ��9��۔�:����%�2���C��F�d~=����QF�FE'- ҉�2��&nw3(�����P,Ρ'��Z�v��%���/�F:!3�B���]^���l� -�002H)
�Fs�IՁ7�6���AA��ͥt�M&�z��g�L¶$�����σ��Y�m�I��%?�t�ߕ�זFG���'����Z1s�
Q׈s��Ÿz�n��+"�W�E*�uSN�1���S�>���X���gѬ2���_��=Y��τe"�W�����G�p�Y��]�����I)Nr�:S�(g'�7����I��v����)���y��E����nN�pZ��?�D)���kخ��p4:���TZ�'!�3)^s
���z�(��H�$;������4ڊ;mȁaͥDR3��a�\����yU�=4�	�_�;��I���EUb�����ԏ������#��p3�0ȹ��0��������O#-֠��`	V_Ԅ@Ehv =6�:�f��p�9W�ܑә���o�s���G"��ɨ[�_V�^�3���q�^ܜ���ZZ�RWzzB:o=���o��3��=��s�6r&[��	_J���vu%�_�!���x)3��,����Ah��J܊�L�)-��+�p���'�}i�:� ~��0Qd0u��<SK�_�Z��SA�[.������[�"y/K�����̷ii#�vӐ�e"V��U�!j�b�)���2]��~��=K�tE�����U_Nܗ����o ��_L"�jUkV�)����P�D1����=�_�	��$��Rm���<X[[���ʔ��9��'\�z���S����z|+CU�S�o~iS3��ia�O�p��V^��B��x]�(����)��ʏP���z�q��[���+�}D5#�v������Y�T;�K0��-'�2�l+��̻!P%)�oDP�{B��҂i���ɗ�"?Z*I����ň�u����E��:�-�@��C	�H�:�,���D�1��s%�y�l0�|��o��<�%����9w�y�B��I{z����J�o�[�<hg���"|Cq��Zr�f��~ZQ��� $�nĮ�� �m�������[$�MEQ�^��6?�}�o�I�aW�۰<T�`Q�ݭ����M�L��p�2����ͬ�	-ނ[7UQ�v�-��\nߔ;�5�W��a��`a�8�PL0���y���ֳb�5"3���(=崋uc��`qL�*�	Οͺl�p�Q�6*�́�lqq9)��JE�y���ZX�0
 =�xB�:$�ĝ�xyy8㰙/..�/&D��Ue��nS�{��O�Ue�/m
ѾW��ͳv0\�\d��?�4A&�^�k�9l���g��I�y�3φ�����CT,,,%�U�ԕ�n�>JV0�ݳ�n���e:�Eʽ�=���0X�_�f}��g�yߖ{9ݎ<v�]<�����Ł6�0ʌ��7v�W��Ύ
�㙆�+���F�@ddwǦ������tj����%�!ؗ����e�,�ɓ�W+�{��lx���ht/��J��~8�	�_�ۜ��60���{�2?n>q�7�w�wR>��D���?}�|D`�?o:�=����{A���9�t�յ�h����"�;9�%D4ז����Yu�?S|\2Y�Ũ]��y�ͻ�*1ۂ&)9������[��h��]��|9hf߱v�Mf�8�[����l�Լ2G��S�P���NEe�j���׀KVl�x�`i�#O�@ET�;-���L�f��֛2���3����l�B���v�m�_�	����y�'��o��}��P���&�Awy����qj~���M��������m�{�����׳G|{.|+Z��j�4��ןx��>\�Fx��A,:�#���>e��v"��n�FvW�ju)*��K��& ���`��S�k���zy���$Ņ��ԕ���ӱ��k��=!�h--~2x2�Z5'h����V�kgGO�|�M �t���X�d�,��Tu�����9+N�����c���,�����h��g�2�i�`	sc-�N}���\��=xk-bo��BY����*�M۵�j�uN �]y���o�В��L�����-�i�]U�/�`.�}K��gR�\�Yk���7_�����k�Zy2�X���04��.`o1��ϭ��.�.V�t㵌W�hQ���8\S,QA�*n�3�.�)���b�+`��Y`��A���~�ҫ�G���Q��ˋH�ڧ��Nf��\pw�v�őd]Մ&Z�Uqd�^'����t�^7��¼mg�q�������������ü�l���-<�F�/n��&�{�B�Ы����Ij[�����~F�7u�T���a�d��B����`N��4��6���'�oϴ>������A冐�~�<p���w �ͼ���,��zaŹ!#u� Pc��	:��n`�?�,��6]Q��F����^x�Z,׺Y�+�E��/��N+�;4��T��B�X�T �*���􌚨G��UDp�5f�7�|Q;s�<���a������W�$F�q��7�4�@7��" �h���*:�<wa�G���۶�k���=,؂Q�}�WL�hp������a0"���y�߭�r���7A���e:�5��$�~�����*��Z���=�K����(�g^����l����wD>�x�Y��l�6�k]��B�:��α��u�7�<�VF*63Mb���n��B�m�%i��f�BEz��	���� �ls>#X� �.q�Ր�)�ul�kʴH�s���Q�A�&H0��;���=:��m�pQ:�����^?t���޷�N<V�l^�k����EXٺ��;.�o��zYwƝ�0Ư���DK&
.{R�V0������b�ܳ�N�׻�{���b��v�G�Y�B7k����9���/���^�	��ԉ���os�����0����%��Q)�vF�/��wY�&��WlXu3�}8%a����ž,�?��uŹj�*�'lN�.�U�,zKֺ}y�ݵ�?��<(v[IjRc��a�+dY���	h]m f���m�g�^��?���-�Q�uL�yBb��޹���O/�����&#|�V��=�hb�ǡaK�g�ӎ�Cay�p�O��Mg�Zb2�n���}o��69h�����P�S�lFlk�򿾕�8ϯ�8�5W��d��-�<�U�����]t����"���yȨ�^�txx|�?�c��p���Fق���ך�Sކ`�E��:0O�����j<M�u%1)�"S_<P{7�O�\������q%�aI+��<A@�0q�ҧ��W��a1|}���C^z����uB9N2����Y�əq4Y�((�54�>�B��l��l�se8���L�x��+'RZ{�		�Fp-��|��/��?\*y|�A+̅��GQ{����"���'r{%�zX�6��#x�E�c��J.���@�[���
���}0��-7��T�Yj}-A�CNg�NX��샩�%U��X���ȣ���]�[;���x$/F�BP�?-��4������v�����5�y�C�nw�kg7�0� 8\%���	�+Q�W-B*������͙�a��G��ԛ��!���=_M�h|h���lĐ�=T��Z�ج~t��sJ��D.���S�_��:<��E��wO�����uU��0b/3���+�FN*��M@�_��|4��o�����l���2ȱ��\�}�kE��	Z_�k�{;��3ӿ2F���%���Q�C�n�/ևH�!�26�{������Sù�	a��j�w�T����Pi[q����45����i���Ј𝋑Y��2;v��moo/���s	ƖT�E*��r@\^�a��kF���b�K&������{	�o��}��ct��&�g�-��1=f����וUj����y��� ��u�	y�wp �(�/9�\R�������l��ԅ��X��B��k�Z'r�8��Ki)1��e�7��+���ѯ�>vh�����Ha��ϋ���$ߧ�ׁ�K�V���r��Uч���/(~ⴇw��Ŭ�����@0z������w��k_o;�&�<8�i�����?6H.�L�_���򪱴��e���M��?�Wr�S_f��� !K�	���㙁۲�,��,���ѢơL�'����e��Z��0��|�	�(���5�F����-��j
Paܵ����r�^�x��������=�U_�������y���M���ECx_��к�]鉼ԃD�e����o��W ���[�0��Z�I4X�b�WJ���t岱��}�%m5E	/�
��m,�� ��jֺM#tG��������&J�K����� �����ɵ!/uQU+�J�Û��l���S��O�<�I>Y�O��{�छ�<��O����=X�g�7;Sl$s��Zd)z� Ia��ݢ���=ڸreE�~x�Ǝ,��$Ҡ?R��q�}���1��=?�x��6,?
0#�h�lԸ��y��
��R=���8'i�Ǔ	�W�]��7Ҧ�Lr�t�\�|���;3.���1ki�E�F���-��O��J�*O)ahe�G�\-�,�6��51��S�Ŝ���f����9�b��D����ﲔ�~j�=���^��9i��f�~���}�a��K	`���	5!�����-�{��vU�R�*H��M#w��C�i��P�)i��ςDRqh��dm�R�7��'��rOk�����o��,��o�&���3���v�Z6�B"ǔ�F��I�/>S'�����n�a��Z�q�����|��x墅�ؙqx�叠�Rh*�NQm-&���eF���6��z0*�QO��;��[�f�����o�מ
zi|�|����1lƳ���|���[Oi<�4���v�GYd��'��'�:�xc�H���݅��*�^�iS���
��:�h���9$����wdN�Jg���Z�����Bx݃��Lm8�~c��v/<���X��O ��7nUī��\��$��*���ϲL�M���b+�Du������m6�Ҋ\v�^��s#��)�45&,��8�*T0���*N6Q�k�YM4����{T�����h
��\n��pJW=5���4��C����Q�����Pi��$Gǐ�n��nD:��F7��g|�����{;�9��9�:�h<��� ��z2ֽ�����������/��z4�� �&�۲�@�$���D���]4')�0����x�Ym7=�E�
p �.����/��^������8��WSߐQB�,ꛖF�D ������zM��b��/K���;>(W���N��-��������d>1s�R���lIŐ��.9�Zo�	)AHh���h��<�	�c4�TΤ�7�7z�����)>��z���[,�npN��O"�Q���T;l4�<�c���k|���|��Q�[)��QpDI��Gţ��%b�3�y��e@/��������;;g9:�k9�D5XƝ;D��@��5oi���
���^����:�6�r�QZ�܊����L��7 ���V�V�.�&]�{J�s�2$��ʊQ�n��8Q����ߗ��=���F���/%���Zjyw(h�p�PV� tƙ:�p-V��o�� �"t{�k՜��ly���T�n��y '�R���u��!�I��.��d@��hY;������ew��T��ڏ��
��Ga���������{4�I��׊Ȧ�}�(

hi�%�o��N�6q��ݻd��G����2��/�'�^K~�"E��LU�� _j|�X����$�<��K��߻S���6cUa;2�4�#��{~�$�Y�?B6��v�G˅���^h���!����7�&D���"�_qYK�}B�ҟ8Ű��I$Y�z3�W���~�1��4��	�$�M%���e>���8����{Kfw�LR��������ߝ_;��Sk�����'��ӳk'�1WlLQ��l��`"�O��m���RHY\Γ���ۼDZZ�9U�[�Tz��p:WO��ܸ]�<��7]N;?�����GA����x���(������H�y��Sx��nw�S�Ŏۈ�p!�C4I�(��q���Ɵ�	P��.� d�$1����B�����^j3�	��9K	Q��<�=:X��ځ����������.���֪]V�cum�ϋjG����Z-ٮ����Ӷ;�P�PiP�<S6"ȣ��(0J1Sˋ�=.Dpn�譡l�>ja���3��m2�dJnL�[h��G�yӯ0u����x�,H_�ҭ��;����x�);W^
�T:�H��~��%�~�U��.�h��Y���ɍ8�|���%_h�P0��a�Ƹ3��!�Ci��b��ۜ��.1��@�����4�]R*�o��$�H�T����p��*o�x�)��}`7�������㾵��6u����@���j\����d׏C��QZ�n�/VO�ev�t�h�b� �w�I�9����+����:�j�*�Ep@��4��N�	�7RL[�z��x���)��FQ�č�8�|�P��S,D��m��m���q��ɥ���䢞�X[���� @�mB:}��[���y���N.�/���P�����3���'v�qye�����щ%h��V00�Zu���g���_kC�̱���
��{ ��������n�����'��g]�M\[����O7J�CI�nF1;�rQ�U?��9�S�������4q�����^��B��dyy?S���G�t2�:(�	�+�[꘣�+7�FtfgHri��j��]m�[ I)��9>���aJ8�����B�b��@�
$�G*r��L�ˌJ��S����}?�0����sc퀧�ߣt� ["�L8Ե�`c� v�.�H��@6�5��m��v�}�����y&�8�d�}*S�=�7�1+7�2�p��?u�=��V������1����\���P7�RHvo�+I)��~%�|؅�M�%;M�Oqnɬ�}36g��׳�����a��+�ԫQal��a���$b �9ݻ���6�
�3bn��\��:�G}�m,�u��܏)L��bQph9����y��4�
����AR��yR�b�O�\���,���6�իv\�r�=�=y�/N��f$�z�]D۝U����D_�����sZ��E�M����0ϡFg�N�#�����ԏ�[��$��,���1���?*��U%��>���e2��7�����S>�6\n''|�c�l�A��z���w>�x�{6�s�dax#��V	� �����M?��FyQC*1 tb�Պl���h�<6Jz�im�񑟷y��%
��؍q��H֌�����Oٛ�vE)�6��"�\5 G����y�T�1�/9���J�2�!7�}���2��Ä&�qU�΀,��&IdT`�����Q9~�xXZ^'���ީJ��R�25MX,͎��1�:�c��~%�995��°���Li.�F���{���Tp|ݪXc�7�,8b�b�Ѕ�UȤ.�s5�!b0S�� Y�w�<2af���)�HPET9sP�5�7m~(o6�K�@�m�#Bû|*�RIQt�<)�|�Q�:P[�A�3C0�&~й��?�>��͵����U�%��w�f�i����-Q���<�=Be�{�_����:Z�m�*N�{F�����V�&*�/{Ѯp��)��M������ٺ~-g�����[�V�ǿ�� ��ڟ:��w���DU�ǻ�ǗY~b�.vr� ��	915[P��Ɨ۽R�Ao�I_�-�t�sQ��O�*o��������D��16ܶovVôԤ��Qy�%bN�8���y!غ[���ѽ��I�+���.9�_������qE�rA����?3�j<~�3DAe^zڳ��-|�W@�(YR��xu$Ő�"���.�z��[0!/t#lc_��F6
�2���r�~}��t��P_�ZB�r���s>��j?��c��WtD�
 �G��Y��peN��ii)�PA ��&�[�p���T�M�
�Q��^s��}`��H%�d���f|��F�:�ܩO�T�e��ٶm�N�h�.�F���v<��ll�V�k'ӭhDf�Z1P�aZtX�	���ǝX�'Ϣ�KQ�f����0Ƨ�ُX��ߩ��}�w���ƺ��!:�t	"��2�Zw�G�=~X�ܜ��j-��{wQ��Ȇ�"��תj�ܞ��|cm�9�Zz4���!��i����[AIH�Ц&2� dD�n�U�_̪�Irg&�3�H�Q�)f�=��?�L�̟��6��
���ȤDϞ �����8����Pp�N��T�椧w��d,�;B[g�s��#�5���V^�� �K]G����r������#�o�Qj�.y3�N���w�鐹z��S�� aV�R�_���b>�eG��������Ʀ�Zo��D���Z_�Hmb�k�39�[��Uv[�����

�K�&$��?ݭj�K��3z�����4sXUh��a�����-�k!J-��zQg��k1�p��`Y�ͰM|$at����XH� {g��%r�h{��FX�C����}����h�`�L���IJ���WJ�
M)��7s��̿[Z,���}�-1yg���S}��g�0 /�H�*�R�RȍH��'�ZU�9# ����X��'�b�ym�NA+�P�)���`��?�zh?���{��8�����Lwq��6�O��$n~X���|\[Ӕkn��=4�?$�\� 8iE�шY��ƄtcB��}6����%�����Xi�L�D�0�3�M�D/ϼ�F�-��f����b��.�7�\�

�N���3��&�D� �D����HBq�B/��S����3W�����+�s�}�]L����*B���Y�o���w���:E���Rk����l-B��O8H��H��Jpv�y=�&��S!��"*)��':��2����kW��	2p������c�[��m�yS��r��Iu�GO2�VC�h{K��Pip�p�t�J]ڱ����vr߼
�1{s�@�X�ԡ�����#��)�3d~s�B[9ݎb..�L&�<j�|؉0O�۫:#��Ol;Hx���(���j�_�ڪ�8��U�̃K:N����h�B�~uy0���w�nG��E�U���_����l'��(�X" �ұ ��k{�q���}�U�ᩛ��SSS��<����@i�:���μA��G��<E�ؘ/�sM"�����Tr-�i'L��?�'4��R�3�y�.���a�_y���6���&��JR�h��� gb�\����-:-���V��������r��eZ�#���0oT9��#�����ѵ[X �o�_|F9!a���|����<{��xĖ��䊹�����;@�@�LJ*��.�6Ń�)5b.o�-_�=���W�״�i�x:713e��Sѥ�X�5�s��1~�\R����5���n��E)4^o���;�c�:ZL.���r�ςikk�Ꭹ��i���V�c����trt�ˡ#����lua=�����%�"r�x��\Ѭ����u1����e-9��Cm��(侲e9�ޚ��O���4��<܎��@_�����k�#!;#ؘ�o%�^@�*��]&��KO<��8qi"'UY�zS>�d�u�la�_�����<8���׶v�x
	tM3�+(I�;sѶ�)Ô���P�@���{�]�(gYk����h�	dſ|�O�|g|I��s�����:06_'�_5Dqs�d<G������ʗtB��ۯ�Bt�̄s����.���,��͆'=$��Cj븗��b?�Ln�u�{�|�2��b�m���$���;85ϩ��'���PM��L5��I��?Ύv_K�w�m�]�7������#n}=e��p������6�"�F\���B#�"C���^��!K�SK��Pf�"�%7A��Mt��
�n���1���ƶv�=!Ƹ
��c7�W�X�yq.��M����Ìٯ}��3����i���Ѣ�z�XBؽ��|�?�������lA)��(I����vS(H�e�J�rL�y}>q7�VJ�-��1^�
G�-���V:,����
�iqs���|ԑ5��da9g)_��.#b{��4=��������{�	��6�ȅ�����D���(�3�"������223&�4�@HS�2�����Bv�M]Cչ	��Djs2�Z�s�]�Q9�j�9vFT	�<X�Ŷ�����0���c,S�A��T���72U�Oa^p'Ml:��������*�����Dp��pI�"i6�)e���@��˯���&��8�p4�^]5���xo�F���tp���\?|r���D���V�s}K����z�GP����~Ҝ�(��=��5���Z����<��/��g ���I6��h�s���כ�6ܲ�o�ݯ����qT>���C+�u%Y9���)�Q˛��=5u���E"���[P�_҄;52��F��>�:��!c <��*����hLK�>QE������;��y��W+~�
��O.<c�ݏ�wj�n-��{(����^ݷf��'c�ZBQ�T@���r{%m撥�MՓ��ذ�ھ�#��y.j�C��5�vA�b$���m~$�4K�T�>X@U��N��d��w�}n)��{��/�>���.��*%/$7y�)�{֛��#�D�r|�K���I����5݋�9�.qp� �է@�KzO�>-I�ܠ&�H����S�y�ܰ��!"@7_/�MMO���oPe-�]!0mZ��ir�6"3��X4�#/�AU�v��l�&PF�=}�9�=b��~�ϙ���LM.��ۣG��##�5�Տ�,T�� rh�)X���p�����5s���\�÷F�
;:���Q��2ܬ�열��~,� �v:g����\�>�ᠷ:��V/�O�p��"�yil�X�Y��Di�~�\�j6���&�R�Oyi������m!v�]�*;���0�Kq� P���[n��EV�Sc��b�ge��V�`1�r�	љ^V$K���#��f?�7`p�cI}��[:S(�%���1G!�D��%����j�����綧��Oq�H���1��m��~����Rh��d���p�{��Q�7��7��n�c�o�wdJ��Rmh�w3^�:�:���jF����)����P޶-7��P٣0��#踀���z�$���P��-f����\O�G0�#��JYA����]h���f�S7�Hi|���Y�>\�p�-N�����b�ddأ�d����2�A��:��/��vM^	>�Rj�b��Ge�e��u;m_���;�`�*�@�[<��3%�]Y)4N.����uz�#����ww=�XRKl~��6�q};��k���.��y�[���ΑG�=�7z}�=	�E��;w�CXd�r ]$����W�T���E˺3��}}�Ȇ$��n��Zͫ5Z����t��,�=#��sMaX�>drZ��~E��jp*j��
�Зu~6h�߷�[;�%&!y���QB�-�ɫ'8P����M�ҝe&U��MR[:���
�b�5����*QbO.`I~{�t�bY:�na�ǘ{�]}���J�U{��M�- 1R2����G��_�jA?���X��U��t`Wbh�v�S@��҃է�����nՒ'oH���nv�}w� &���g'r`��x��z�eN��}~�^�\?<Oq� �#���bgM�AAv��6s���I���]�'x�������R��!�(�W�*�"]�	S��8�~K�%��5y�GAMT��s�(f���͎�ܦ):���9�{���~�׮���[�G0s��G[%G[%�����់l��,�iYqW�+�p�#�g�1%��y�`�P$P�d�s�ģ�Wn��4-$��^�	4bE�>\b>�U��/�Mhhg[A:�o��0���hWz[�����*��9w�]���]������VÆ�Rj;Se���(�Lz��?���҉d�/8��(�&�j`�~`΋+����rnG�u���}���~衃i�>`X`��m6<��;���N��h�MmZ~�����Υ�h()O�]y3�rVo�p�C�	b�>I�z.f@=���ԩ���t2ep�*̐7ò�K��h�R+�\��[�ݝ���%��b�Ä�y������=����~�ط�����.!�C|���r\�x���zp�72`6���/~I6rJ�������&�i}����)��:�C�Qs�W��[I+�7�`�_1��A�?رJrn��.�{Zr���<����Hc�D���׻7�cUĝ	ɳ��͍�*0����w�U����rm=o�8���?���~s��,����}�;�W�6�s-�'�.A��!l��m�s�y�ؗ�L�7�l�\I�ѝ,w�kF�`o��mh��Ѷ5,R�x�D�wi���m�Z�=b�#6�v��j ����{k���$e���k��kV������B��ŁNL<��+$���D����1qWK3�V�,�L8�߅(��m�(�/`�IZ�P�ƙ����̒��I����8��v}Ӂ-�*��
8�9�٪�{"����nU�w�2ЍC<4GD�(���J�i��j��<J��o��ٙ5�@��.c4�_���v,x�~�����ۙ��R�����鹺�	�����	�tAH�P<I�u c!Z���D"�LYQhH����I��@+RZ2V��z���J�����蝚�ob�-w�T��8O�y���|��=a���͹��?��d?� �М�<({��F�_`��u���#��(�V��g-%�z������j�y�-�;
2Z�p�M������a^Ͼ���T:�3�����r;_���':�U��"iW�+N�ΉA��lƚƨ	�z� @M��Q����81h���_�ܣ
��y�Ϋ��1�`�>�� %q�Ƙ�����p���d�a˭�K��Ki�7ۣ�&=�5�jƒ�d	��wzS�����	�?Yv����z�E�f���0G�[x�H3���}���q�+��Zq�	U�*C���f<�{S�3�au�&�l&�⇒`/'�@�:���q�A���|�K	�H�D=4J���^PT�Y`��D�O���{}���of�Aj��*ڇb�ڹ<��������Gҝ��U�:��@�>������FLە���V�d����8��GKf6�5���<F5� eBN��;{rW s���4x&~/F�)b*N|���M���p� ?g�o�F���糮�J1ny��ȕ
�K�h4J��n}Hm��:��2���S^ac�!�{q�B��#��,;so�'Q� ���5B����`��/���������6��|#���2�՜
�;o
���|�[��xF���К��A:?�EI�������)�q��ũ���$W�~Ŭ���̐R.�$�:~�p~�\שa-N�[�7���;
�U���w�pU�O�7�H*`��9��Z�a#�v��D�6,u�v�i�f��y����y�[U�yUr����y�_��?�VɆ�Θw�]l4�0#�12|ii���k�l�p�!h�)a�m�^
tB#�Z搪�1��X'M���;ݘ���0����˞P�<X�Q;4G9������ N5�h̽�q�R�;Wr��~wT²����̅��q.�f5����b7��-O�)�x_�iMn�zA}��@�Hr����r�*c�3����f��sH��`�2(w��9�������;��ђa�f��u���F��<y��O�K���)�۴JW;�D�|}c.7�M�rn{�b8��,��x����;qI�?;U�&����l�H��MUu�<�E��Z�X�'<����	��I��Z�Y'�r��KmGA��f��8�|^�N��I�0a�Vޤ������u��3�7�P�'����yX}l?���g��[��X��}�t��b�����V�~"�P�AD�V�^N/�Y�(��;�ABۀ�'N�'*�oP�N:pT�W+	���sK�q*���D���Ò��1	��Z��@����ӡ4>ʔz��/
�^���k����|C��nM��8�7����N��?sZ�5����S77�:)#uw"�*�`wڼ�gb�tF}�b৤�Ů)W�Hf�f������.oy����sH�ٕ���*��DI�bRk�@(i\��^DZ�D#r���(_s�f�8Y�:WY�y���qi��A���/��'�6�s�QM!�3�A�vP�W}�AUN��MF���ت_�pQ%�+����|M��M�7��XVU��[)<"����BK�f�G���Ό�Y��w7��y=�5�=˨�p�P��P�|OuyЁ�m������-EW����&���z��9����9HpAV����a�aDޕG��:.s����TJ�ރ��c���Ԙ����� փG����h ���xKZ�.���s�qO�Ϲ�fN]7�#��R��@�J)�s�����:�qh
��:�������\��\�O5E��S2e9:cZ�������	U#h���3Q���T��A����A]�|������#��ű�bf�n������bI _��41���}V�� �_��>v}�K}�6��;kO8{|gDnp�q���Z!E\U͞3�uU��ϙh��)��@i��% A	q/���t��U]7"�#d.%�6Sn��VL1���0D9(m�$CR��s���?��l�u,N��m�=뺈�I���E����/���W�?��|$~�\f�k~va��Q��E
��(�JT����]�&�n�3�9��(#$1��
i�eH��Ǔ�n�v�9�5l���&W��|]0)���n�N>Zo���[lzZ%�./',>$�.F�׬������ߔ�&����s]��ư��tƀ\5�9�P�DK��i�V���R��\.筎M�kX�EV���&$��~3�B~,N�I�~©/�:c�1�6�h"�I�'vU����g��o����x@��tD�*�1I�a��w��R���UE�W*�I�X>Xn��M��PW�N�i�5�<BH�����ߋ�5�6�Ct�U�b'+	e=��d��eB5�,Ӭ�BڈUR��9�}gˇ��
^��`�d��l?��}�\�1�#���Al�q`�/�N�3���Ģ��6�8y@%�@����m#g��Cc��%�����˷������`Y/JI(�Q�f>6��	��͸Uc�\B�\�~p���|x�+���������D�S�(����k
�E�s~�������ZBCS9�@�K;�`���!�Q�_ID&���$n�4�
ۑ�`Ẃ׉��+6�d�͵%��7M���S���� o$?�EC�<�u���N�v�j<o
�V!�t��O�𑆰���Q�>�y.&71)Ϥ�BU!���=.u-�D��Jo������]� ���ݫe�M�;YI����h�܀�>�lZ�;���X�6c̈���f����yxr��aD$P�z�ʊ��&n���� ��*��Kf������/kA��~��j\�D��^���{���ԌwX�I�\��rF ,�:|��!�1Rٙ����~��Ap���o#�tڲ������߰U?��'����Y^�qI�P���'�2�	`���Ғ>�J*�F��-9�2j�dU��f3=�@t֍9�Ŵ�<�y$�p��jӖ�ܵ\��^g3Y|7B���i_���xJ��h�6����^P���iw�1@�Zs�d���P�͹�G�w��{H�9ʶ����%�M1���_���?�*n�o|� ��,/v�˯��r��\�qU3i5+�5ńo�[*��V�����������-	��)N���#��Ž�n�D��.f��z�<������ϔdIm�a�܄޴O��쫤����o�4qG�Q�J�P&erV��	ei`�&z���M֟9��I��(���f��Hdu�}[�0ź���>4Z%z�l�$bg��gjs@��Y-��ר�g�B	�^o���7.pO�4����@!ta�3�MSj��1�5��j�]�V<2k��:Ǥ��j�?ЌݐK�d.#%���m̃L#:ڕ������[�Iob��{��uP"�[;:~ �%lR��mtq4v^qл�-.a�Tn���d�5e{u�6v��
���|�g�z���\�i����S������ʣ�p���vr�$+wzr��p������r��WM�Y��]~M�-!ǐl���%�?(n�}&#l&���`!D��$�W��S��L��ލ���z���#�,�
<�M{���1�*�p�׏��s���i2<�M�j.�Պ��d�.<����K�̉�nY�Y@�4�BrTת�j�y�1�`ǣ�>�s�D,ICȶ�ф�
���|؆��߈���=Oڏ�]��ZE�K��j%��(~UA:H?94��p��0�We�&�8^�q�֮��� �Q`���%�T�U�$��rt\� ��������ee��]�c��*?˷��*ꎪ�H|
5ܭ�� �oѧ�'u��-�[��N��?p��?6��/��o�~���oG
���6������>׿9�#Pߐ� �Z3��ꥮ-
�Yݟp�@��6��-�/���y���zˏB����%I¹S�Qk��9R1Pp�x('���d{p��N ���=|�[p��l)/ے��K�r�I�{�X�m�H��[��ɼ=�P�M�<�����h����4RQ�\����SE��-'����7�tl �:VCx���s�0�o4���~Q�+.�(�u�h���+��2/����eP�7zʤ���:�y�C�x�ɾ��al�[�^q$>�+�$��ƳԎb�}Wo��^�&�#,yL7�|Q��1��>'�R���&��/d-��e��ݞS���;��ށ��Լ?�K�^p��Up��ņ���AՉFآ�L��7ZU�,�������=WU�&p)ɜ�p�	�V���cH>P2m�>�^{�P��.�}�{%�M��{ji?������tUx�]� ���	��:7��!��jIT=��0,[}��>�W|:L����1�)�˽%� Jx('ח@GI½������Z$���͛ܜJ��<JY�Π/º����@��ӑ� %�����Q�G]a�B��R�C���&��"�咑F�����딮kT_���D(��=��H~FE��� �5�5�lt&K�M��j��]=��M4��$�N<v��^�)����LG4�	��]5K���m��d�~��:�;D���u�W�Qȍ� 1=��xL\'��e�j>F3��|�&�Ξ����xm���(����H�'����*��v[N�X,���7����C��T{������T2ސ���D_D�ꃁ܏��}?|�6�M±��~�X��i�Y]يԂ�=��FN�]���s��R��R}B3��^�'�eJ=��n�����2��_Q[���S8�֓�%_H�{M��o%�2tAa�F�^�rP6c��h��> ��������7f��p�-�Hxc|�/Sb̢f>�|r�����:���x�|!��cK�]R��d�_KD�)K��r���/P���zGߓs�؄��ȇ݊l� �҄���@�çU�V��&e~�*Nk�3��ӝl�(�O�A����~��7>���~k�_���&����	��GX��1��-��Ĩ��R�F���O�I7k���)�ږV)'�evt1�{zi�Q<�{!VX�P�ӥ�J��{������iF���O���!�+���V�6tRh���P�!}Jo�8pr)��=�R��Fה����F=���j��5B�t*��|k~�-��-�\=%I�T�"B��'�s��wG�C������۳�.M]�n"���W� �dC�ħ6��͇}��W��\���+�,�lH�����d�v���|"ؒ���Ʃ��n'��*!������Mc�Kzѩ�"eҜ	!Z�KT�{<R|wWf�J�����@��{P��ygCХ�R�>��#���}�lA��l���p"G�;|���W��Ŋ�Q�[W���v��)�ݯ�L)�5��v��gB��d��]y�t���P(4n�\o�8�I��W�|� �9�������p ثӕ�{(87������d�2���.+�0Kq�)�r�|\]r�M}␘vH��q�[��&�"晐�SFq�>�/U)��@W��f?�H�H����(^l���T.{�S+�8K`���b��pr^�dW�lQ;�::<U�?�^ihH�<�@���0�U���R^�bB��M��v�=*^���'���Y�7������� ӭ�6����'G������_$�s��*�v�vs#+�iHm�����a7�X+��2E��-�P�[�����g�����-��e� ����=K����:c�V��r�͔���i���"�A�,۞n�]�f��X����uhd�{�[�#k�2�zD|�4��_�h"��YD˯��9B9]�(�.r�J�{÷6Mg��+�:Yo���3=��z�N��$��2s�0B'O�9[��������%ȁ����*�覦T�̳�?9~�l&�C�0}%Y�C�_��e��<���qgn�δ�O�W�q[oV�$|�1܎��l�H�pa*1^�.}'�&f9�l�eM���
�R^4ԏ�U�.m�3��˫&a�?��Ix�*<��FX�����d�a�.Ȓ;�\�N*�+},0�JGC `{�u�2
gt�[��	��Z��+�T������[����&��@7A;���<P,P�3�ٞ��U=M2� ;V�B�	EK;���n�V��+�C�J;�Y�0� ���$w��"4��g���R����/-Mb�z*������/}Te|ޒr��pVw`"��H��@�%�Z�W����"�Zuז��aOY�:�9u�J��ih(b3��jo���E�ڽm�J
�o���e���b�d�'U�4t���:�U~D�I#�<��MjG��������A�~#-D:(�L�ԾW��ۿn�k�dy��X�j���;EQ�P��/��U�ē�6vŚ��a�^(����)�
�%��A�zm��q�)}�3bF<r��y�9*�����W�6�M��߆$.�*�k_"��"1�MeH8AcOy�BQ�FF�����|�3�bh?`�-[Ce��� ̎T؜˵��Vy��$X��;���3ᇗ�-6�Yw��2�ѓ*�����>�:��)�^	��bs��)4����<uOG8�������/���v�h2�M5��&��7�N��S)l��4�{m���ԣ���]觖3j�� ��s����/���@C�����2�(��n���BC�_[/�M����Z�J��in*% �+�'
��̪'��q{W��,�J~ji:_4zR۟�Jͽ�m�Z��X�QW��JҖ9��d/�u7��u���hj�P�D�l��Iv!$����T����E]̸��/�����2�#�^m2o�?U�q����Zn��=z.���*dODW���;hZ�&�S�H^8?ޔw�-z�$��I�._-/����	<[��'��<�c�e1 ���ͥ0+���<`��0ܖ�U9���б�Ƌ� ���CA�Ï~`��\�f��P �w�'1������ڙ'���w��|�۷���S�A�Φ��|U�e%a2]������hB�w����0����ҹ�^4�*=!��|v�8�k]V$��3��W�$��w9I�x��D�&L�Cl�T갯%e@R�+�����C���y�n�ԌO�h5�s�扶ӳB5�d%3$��8;��M��;�=�x\�+;QR���-�ܜ/˜_�a��\���d�b���%Yo��Qb�q7�Ia䨰Ƅ/N��t6*y���}%8��S�<M][[��&�<�/�Yr.���t4,��uS�>%d�~x����ji��@��������{���՛t�&�C�Ŝ#j��m��h����;�~����'�^\�ݲ&���o��-2C��2�I�Yg�hn����]D��@T�Mp1>��}��#��OĩW%���e*޹���]m�+���T&v@�^0/���]ﲬ��ut�[hN<H㇉��Сd�>�%�՛��i#�_<+ /����Y����B�n�[������}���sz=\�W:ϓy5�$�%��U8���%��Ť������U���k�(��j�ݿ��E���Z���HU�j`�����:|# =5.x��B��.��Sy����l�z��H`�#��b=��x��"DQ��#�Z��s���������8y���[<4>R>��VF0�<Q ws���M�ο��;��k�~���7M�7��T���kΫ���w<����:2�E䧼�h������p����Hź#9��`�vO��P��+�i����p?b��(�`�Em���n(Ky���\�u��ݬ����a� pD�	�՚��'���K��� �}%��r٩:s��e�9��*��9y٣C`<$����*)`n���6i��c��gc�:���_Ȏ��JP%6����[o̗��z����'Z�<(�P���Up��U-�h,�t2�[�~��!�7�Oq��M
���#�@��N�k@}��9�X���
���k�y8�AJ�ʙ՟��óю8���\�}���L]>a{l��^��n����d����Fz`/��ma9��4�?6��A�X�f�B�y�B)��WU,�E����P��6q��|�~_�f�����m�Z��A�Py$�����8˯,*}� :��Yk=J��ҍ��g�����56?׮+�P�����	�~�AȄ��@$]`	���P������-����{"��?�G�i�����Y��ʉ��>JxW[�c�#z�+R�]Ft��\�ͯj��|ZU+ːoO��'*b��}�3������5d�����+���^
�d6cTܪ�8ּ
(,`�		럯� F@Ԫ�,H��hmE���ߺ)#��a+�ǭ�\KZ急�l�����ߏ<��l�M��tՋv��ti�d�(J5��g����t��oy�2��[���^Nh�n��w�>��{�i��+�rDժj��q���j�7t��7�b��-�c�ڧ~
dWV[�_/���sa�����y�ގ� )Q{��*k��q�H�n]s��-R���-��D�x_4�����%��o�t�NS�������`o���;��U �>z,I�J*?�Y�G�W�i�zኺk����Xp�*_C�����b�����	���*��K7"7��f{F��^bI��UI� ��\��S�׍A!�ԉ�!� #GD`�5}�w�L׬ڣ�sy3��� =��o���a���,Io��[� �҉�_A�������T�#�'���z����Aav����SVlM�z��� ^yϿ5��D�V��D�I}?��K����oDu�=ءd����r$�\� 59�(߶T*J��fO��W.�
J��.t҅���У$�1��_����<n��~EC�4��FQ�W=�pzz��j̺>��nK�U!��%��Y�Ω��8�%���˚;l�\�T�>U��H
uÇ���#���É�^?~�y[Ki�WA��Pw�i����f�t C����lF�x�ߞ���h�O�՝���Uo��u�V(Rܡ���C���ŭXq�]�;w�����z��ߝ�g2������k��J�׈r�|{�"��쏞��o��/S�Ѿ�䛊��X���U����A�Po��Y���5H��2%V��3z�B$�l)�����I��;����k��j5�iS�Ǵ�.�ji�j9��▰W�o�:Yk�W:֥n�:X��H;�B�ۈEz���E��&�k5}ҕ"�H<#;��(a�����ޖ�&�D8�6G��9;|_�f�k�_��kS7@$�T k�Hv���t�`�8��w�]�:7쮁a�[����J����\m��r'O�w.�k�Ȩ�P�xՅ�ޫ�����Cwl�~�� m$x�����BHf�e�����:րi��qO����Oz����њq喾�=}���R���5r��#�8�^��e֪��S�Y`�1=��	yeeZZ�9ƹqM�4u��[0�K|�����(��[�<]�(���I�M�G���ѿS�����^�【�g����Ɗ3�Q���]��ߦ7�7��g��l�D-�-��1� t.Z',��2��Պf���/a��ǰ���N9�"4P-��3j�l�v��﷗�j�5�:дE@�Q�?4P_Rx<�>v�����BƸ��L�c�)=x4�$��H�[#����
�g�l���)� �/��{x�Ң;�-Io��q���ז{��v��f�g���1�[��	,�b�@�y����p�E�GR�uV��z|v�ldg�����w�6��P�u��Ϲ�����Zk����ǐ5i��q�=j�^/p��	i>_
���a'�ka��߮aM�?��>�+��d��R��`鮪��6g�;������Xp���|HCwU����c��Lq�ٯ�O�ܛ�6����Չ�T�Ld�YMn��Wޘ�q��r����_��%���<���"hwp��Q�(��BO�_̌}��makh���QTU�c��*T�<������&����LS�KmP<C���=..G���ݮI��L��acC��a�L��f�e�H��XoO[����Ewi����a��~�y �R^��.��b3^��u��@=���_��߆�@��3G�x�)C�d�;<�67�`�����ef[I��6_�X�8��?̖��/���v���.���i�FV�1�0���H�p#D���'xP$�e~s� Yش^���ϻ��_�:����]�1���D�+dx��]����rU3����A%}`��F�u�ju]2P�1�V�ߩX�4�@����������ҝtg�c�,+��N��A�JQ�Z�*�["���u���JUe�;�-#e��-����O����ڭ[H�I81 �,>}nEX#	D�����g��ae���o��Cr*�i�U�~`:���Ӑ1K��hRn�Ms���/�/v�8��,V_t۾"�f���Q�C5Eee�'K�q�h~��7aR�}[�E��#(SUA����5��;����I��UQ�qX1����y�I9�1����[���-~�{�!���7{G�`�1r�^��eD��Ɨf���e�}�J���ʍ�~ͬ�Y�G�o�:-���Ս��6u�lB����3��\1�*sЕ[�-*�����[����_w9��q�{V��^]�xrgC���?p/I�4�Y�����'�,Ci\S�>�%�~���+8q���F���#��#}��so��NH��9O[pD�ƭb㔛��El�(Q�ߜ��f_�)ů-̃3�UȪ916�k�\w@55�/ŪX%�/�L�a�tU.gzx��R7�dɞ',xzl�m_�I��s;���b���U|�[d[�'�6������*8i�:��%�~?�)0l��c�Kog�E5�3i���":�ٴ�d�"�m�ڄ�<ԍc���I�ros��j(6��$���z�����1wl�~��a�j��%l� j�y�m>؏�*2�'�[��~&i��h��y�@��Sӝ~�h���>�W�<�����M[(0�g5�=���6���BX��(ٷ���	�^�o�����I��6I��B϶���T�������vg���,+�,f�����U��y�`Iu��5���c	9�	�nݴ���(��q��M���x�ϙ�u����>`B� ����mUa���_-_xr&��)��eD�S��[&>
����|[��^0Ll�Kh��u�!��k���f玜���(3�q'o!F��Ʒ�'�c��_�t�UK)̙����C����|�»W(�B��u3��V >�	�8d�{	.�U�,Tj���y~��g4�~DJ��'�aȵd�E�N`*v]&ᔙ9�,��U͔g���2'��8�|C�gR׶������ LY2��v��X�N@@Pm9G�y9D�nL�+	S+�T{0.�E�~ ����2ôy=����D^'V`����.C)р���Yy�ƴ��H�T�H��-:=�nɌ�n]a/�X$B'~K��d��@N�cϪP�_���z����#�߁C,�XϷ����zneIFb�1����7�����}#��I ��i�'�*��U��!a���u��f������ij��mhZ���7��yI��dx�&."t$�H�H�� Բ�9�m�7�,�k�TL
]!��)�F:R
Y�2�9�B�/�����+�u���Aqyy_$�:t�#��_�+���ő��r�LUm������L�	��p����Svpȟ=�SH!b�GD*�[�|#���ض/����\Xx淳Cw�ϿYƃ��u߳�����W\tp�))�5�>���;m�-�W��6�zC���y�_����0����N�Vs�>c����AFH�!��9��Cy�x�������ۢ�WT׋��@�Z���h�vaF�W�?Zo�ݮ~�Yj��.��8���"7]c_�k��V�=!�>!�o@<j�9�آ�1F#���c�x�����8�f�8�ư7�GQ�G����� ��Tr��q����x/F�8t��Vy���*��k�;Nz����w�p��\bfcM�Sko�U��n�V7����J�jVv�pt�?�)ָD���n�\�o\/-���:+j�N-��J5��w)�:��L�W�-���I�,:��k�e�Qi��c�6�K`
�΅�b/g����UA���Qwy����C�d�^i��~-L�t�nX�H�T>��3~p�.�_b�mŸ@"d��п�Nwx$���5�����ǃQIP�������=�of{f���@a��RR���b��c#�\� � Qj�X�	Lt��o�LI��!�N�ZTy�]�s#�'zpQ��'����Ᏹ�[v������[�ܟ����?T��l5Z���'|��Ϯ��ȴGH<�߫W�E&&�L��ftv�i��*�F`:QC?�X��i�Iۯ���J� [jZ��y����VUw��� l�r���8�c��͆6�<�8"tы������̋�:���ҒB��쾔��1��쯟�|#~_�O�����8zGB��~u ���,��N�<oH��fk�|j�3��a{��ß|xu2�� �U��.���[�
���J�8�~�|�C?c����z],&:��_���?Egyi�շ�HS�c�QclW��y���4��Ђ�O�s�Ǐ�_�ҫ � ����`��	]�#�+�*�h��Oc�V-������ m1���5��ZӦ�<,��m`��r}t4�/<.�W��õBN���T��T�����d���:���F�蟧�'OHl1*QH����\h�Oa��U�����Bv&6���Q���q���(�2���@}���Ϩ��w�ͫ���x�끫��:��8Z��������Iw�/A鍺���,��X�L-�!J7A�t��p����1�1���E!ť��,�a�M����h�� aJcJB�Ll:u���5���Z���@̖�9�A�Z��Vq6>\�ff�v8St%]A��}X�k��78$�2�Q`*H� �n#&X�̹����O:��&���,��Qeyb(��ě��N�ھy'w��Fd�J�HOYy���_]���`O__�7�7���?�ؔcV��~'���6]$Wգ/+1#���Y���N�YII6�bΎT��������caa�����T�j�|VU���{��>��e��5�ڧ��}6�##uV 41{�0abW��������� �rE�()ޱ���1��{�����T�������v둈����@���rE�#�m��Λ�pm�qsjb�p����̡�`gb@P�DA� ���*k��E���vo�	=���Z_������"4m����Y�:&��i��|�m�%}�*�a�$�;��_1��ly����)���5Asȣ���臒�(	��e=��D��'@{@���N��m�A�O�]g2��[�T�m�`'�Ev^۶o�D�M��l<��Mf�ps+\��T�u��ؖ팊�rlD�^�;�"H�:�#ۈI�3F��)���rJ@�O+Z{D�������O;|��y������/zM(��֯�0��$(V�7}��h�ЫW̦���D���>���̪��Z7qW���H�Z�(ԁ�MN���㡡�X3K70�݇��������
�t͇���r-Dy�'FH�1��Șa;�[F
��ó�{5�xM/�"��:��a�tv��r�]�-
�#�q-#|��
��F�Β�\���*j7�=r�G�$!E��C�i��Lp�Ӡ�	h�[s�+ ���֢Lh�8Q��A���(G���Ä�G��R��,$;����3v|V{#_Y0�t;�-ꟃj�=��V������Տ�>��(��$1����!M��2r���i��MC>���\�Ș�<}R�-)�˶�P_�Z��	&�^,n���>��H7�I�p����:�j�Ս��������%�;�H
�̱GCJ�\M����1�����YQr!�߽MyY|�{��)�0���� ������C̱-'�JH��B�"׷e�v�FPL����(}�:%A�R"�_n���5T7���	�{�J�VH`��ǎ�`�.YNg�Hlo�j�)�b��5��w����@�w���S( ��kA�Ί�Ts����x��8�P��v찵l�� ����gO�I_ǈg�:(�Y �[���������`lO��<.3��76��9D�5���Y�����V=���_�|��n+v�.���Ș�~)U����g�5o�J}�"%ƻ�z%#��?Q�D�6���8 �U߇l���(��_H_�sW4��vfr �bE����2��Y�0:�=j|�R:�'sPs������nL����"�G6%�_U���@	!��3�M.-�;|?�����.�w+?I��N�*|�j:�q�0�2}W6�>�x��@vGvf~Rh��Q�����,1��`!b,[ws�R�W���w_vW4�r8��'���|��HUZ?�q��G8���������C|$"Bh�g�˓�Ƨ�eN_.�<�Ľ�%�#�t�^���]�c!fh�B��-d�~g�|�m�!� F����jϖ�"���~���Q
��[F��l��}����;��ng�ʐ��x!�6��s��(���@@�{dz�F�D�Xp8�CU�F��kd4_����9����U�ݓ���U٬�>���ɏf���k��o���%`����/�!���G�b�p�m�+#���{����!�8I��-ɤ�=�&sL2$5&*;��2�rdf9@��s
��Lo"P~W�J99�Q%�x:�s�O^��_ڳ���9|9��D����_��<�6�9D�u}�����*��	��vMpH�ϵ��J�b��m���7H��9�
���|��;eF�.��=c-�z�=�~\��a�E=��5�6p�,�ujz��X9dEl@�	֪mE�bj(ƶn��d��T��Lw?���	�j��/�A��@�[s������8|��?�K=�0��!+P�c�#�?Q���7�}�G��e|&_�\.k�ި'�Q41�tnmi�%�X�׺ :>�~g:ml�/;C��mD1M�`��O7��l����
f�^(q�2�~=��8�-3�;��d}V\П����t��Y)~ƿ;�4��~Mm����d��Ζ ������($2�w��{s��XMt���\������$pV�d��?d��0�n�+��������h~��dw�L�\j���2��6k�����J^Ȣ�g���Am����9���ȁ0C ��5�AYmA��Ω��ʎ����6�\3�� ��b���%�.���\�mG�R��)ύ ����S���j��zY�����jY�:����Wh�K�j��H�fw�í�>�3��.�¢�ĩ ��lJ�F��P(�h�cP��`R���"��(Ivh]�N�vs�D�9�6�8׽�t��e��(1�M��
-`2��*�kNSh;���(�#E��nm��`1�p�ЏͫW(�`Hv�6��:? �HT[� ��e��b��)��i[���4q��-6B��)�˖�j�+PZ^�����2C�-���̘���=�>���Ft�����k�6�`d��sb׬�Aa/�Z�2�K����oKO�\�al��f���	���2�9�8�bЄ��v�1����I�� �W^ߥL2~Mۋ��}�GgI���bI♖��-3�n����n�gffd�[[r�gH-�>.o��uR㻙Xm̆n�籓+��V�:�I\��^�Իo-S����>I}�� �N�z�|����?�QZ���ME�]Z�o>�8�T�AF8R�d_ɜ]X����Ĕ�(~#B�P�5�l�`���\B$�sx��M@���_�ְ�w�S��Yg0U!����*������3���w8	��66�a�~�y�"AH���O�kPz��#u�a��3:{��/�=��}���hQ�u�P����yQ� O�;��p�n���n�L�'oi#{�o�ĭ��`�m'���MD�
纟P �{��MKӞA��6܌�0�_�d����4�~'E��j�����?��:�%C͊��ј�1��߶�*:���N��ɀ��nͣm뙨���9�I�	��8��$8��}^��u����@��,F���M��HĬ�`Ez�D�s���W|;E���+3(�bN@ �%N/tB��L�W֍��U��}����ַP�w��0��$�c�GW��n"(��AĬ��㸰>M:��Y"'��>���Fn�"��e��>�X�?�P̓�����J�V�����Y�\A�'�˝���N��/�1
:���\Є�~�����B��sZ퇿��<_�e�i	
�WT�{I�9�>��,�l��p��yB�>6����{)L��T��$�2��q�ֱ�;'�l�;��u3��e��5<�øl?�[_���
��v!�h��ѡ�^RU��a.fT�r��L��w>/�q`��DL8v�Kx��/
���� ��|����r�߄�)΢[��4p�ɥ�{|���%)��?j��~�]��K�^ƕP;�r�5t��3[WT� ���-���b���łd�ρV`k���K�L\ǿ9� Uk�Jɘ�"����w�_�r��Z���_��"���}�����A�w_@A�n�c/^5J��5��(�(����������Cu�w8"wx=�-��ۜ�ؑ��T;B��_8��a��&�Y؈�6c��UGM�/|��M�\��<��a"ɒ TcÝ݆As���l$��]_:���)�R.&$e7�V��O�-I#�������?�9OΫy��BV_g���$O;
�k��|Ujr�)"�OY����T� �3>�v_��Jky�^w�ܯ�d���t244|��Jv(7����X�/n��ao���%�
�/=�U`�&a� ��EN���Z3�L�����V�f�I�RM_�{����ĕ2��\�g{%In<K�[�T����u�w��ԍj�ܫ��f�k�b̯��s�'d�]ɔ~��zb����9� �JI!1�5{d�Ϋ;��L�Xq6779������g<e��8�8�-��|��UX��٬�i7��w��n��j�}|�~�\��MD�n����K2�>�2��^h�/��o���U���:�� �a���ѿM����	�-{���Q�;��Sm��	�,�2570��5�t4�Z����e�$��Y%��(~Ta�U��l�Y�t-�+$���&�8����:h!���^����R��^�֝��ļ����[2�[��z-x�ˎ���3����
��ZΌ.���I�lT(���?�-�a4{� "�_:�C�Hrn����:�����cƎLgv�~�21G��(�"�Mt�ԋ�TI�ʑkK������໎R)Pga�9�?K���n1��Qb�Q����p̯e/W�r�oq�Mrd0b�:P4�6�6Y�y;mdd��u����@�⋮;�M�׋���Y�EI ����wz�� ��̂��b��759���%���+�%0E���y+;�Lb�_�h�:�'n�YԐ3����8��l�ػ��i����,M�Y��ʼu	U�[����޴ �z��˱�qw �O��$˘%1��U�=Z���KyIs\���a�AT���q�K�U����O�����4E�@�GԆ�W7Y�Z�v�~�E��ь(�t ���\-v�h������?��oOX�� 2}d$+��	&^��S�
z���W%��TI6�ݹ�Ʈ��B��]4{��ۚ�������M_�u38��Q����^�X�NJ��_ĝǪrCm�����Xꠧ}'���
�����MnN����5�@�к�S.�1�`H��*B�����q�V��PR�p��NY�"Y�����%���p�"pG�ر�"����,o�$��|vz�?/��b�����S���-Be�4�}��C�l0�^\�O�˝�|(~:�<{�8�w��E�SQWJ��i��e����#�F����e�vg8S{H�L���垹�y�o[��גn���>X��_e�m�ǉ�E��+�e8�,�w�e���D����9�N�%���M�
�Xg��tG\&�����:���S���ZwJ��`V5������`���(O	|�SV>�n�Fuj����l�t+���gt���;#O���6���I)�Q��*=L��7Yt�L���������E���y%��?�;o�9!�N����ּMvL^�S����pӪ��7&XMD�G�0��#����7�J$����}5�^O+�V��R&�b���m,��\+�����(gV�<ɗ�q�O�h~[�?2���z�/t1�)��AeX�U=��q"7v�b�L��ܱk����}6ӷ�Ӧ�dP�s�C���J�%�xv�_��i_R��Պ�x� 4��������9O�rz�?YLa��F������힧[1=(wӇ̹�[��q�Xn�_���)���gq�E��,<�����zP[x�_���(~��#u�����K���?,��������o���鵓��rp;���di�6�uߖ�,��i��'z�_G!J�&Z�&� yO�c �-��C����O�����z���@�jd`0��f�'���&ЕK��L� �M!-�
Ǻ8x��б�lW�ۦ|���$}����`8>�Vv[/������o�a�)�j��ʐk�p��ݷ���UYYu٬�mi�s�!�i
I����NŒ3m�fn8����Lj�r���?�0��=�����0G�����v`&΅�.�~���g�"�n��M�`����WY�.\�I�ę�p�� e��v���վ�/iLQ_M����d�������b��%��U��oD���(�e�1�����oL���9��f�\�FV�`�pJa8�[�R��-��������!|"K]��*''��݈�R�a��STQiN|������p.���]q5�|�¶bv�Gn}�t��������z�f^����ǰ3�.K�H�g-���M
�'*e�*I�̃�����X����Ј*�(1�7~̲�*�0��;}H4fe�z��+۞`u�������z��2�d�b���}��b�;�Y�Ԑ��������vr6��%Ec�j�ülb�vGC����Ǫ�~G����ᇫ��m�i4�H�����&D�)w���e
�!"�H�Kϲ��%p�8��A��Wv�C	GC�w;�b��r'�h���h;�DزÎb)��Oϼ���:��K��<�������;m:�,A_�I�9���J"���}!�I�i��\c�a��G�eM`׹\��F�J<�4�c�O<����`B)g���.m�T)��� U��L����R(����a=���H��"��`�}`t�`a`�)<�F�}A��b��Q�dU�̳v�e��;urXڢ��9�ja�[���i냀�f�ՊLK �T�.EH��0�_��mg��M��Os����G`[�щ�%���@�A2�y�����M	zD�Ik?3$��vK�X�+ևx�J�o�,4�M�Al�y˙>�᧛M�t��T<E�C��tV�yl�gx�/4��(�� Dc�`"o������x�]�$n��Y�'\��ci�w).�,Q������m�4����H���UZ�1�gZS�'�L\�w��H:</���� �=�_h�R��ZJ�$���e�tM�y�b���{�"���k�M�@�_�t��,�S��oרC0��J;��H*��6���A�UW�<>��Xl��U��t�_ʐ������/�&��U��x4�Jo���L�OҀLl�E8u�	]y��v��"����O��Ih!h���R������!=ɫ���.T�����=K�
����E�!p�>��aY
��V͡����1�P����4?��� i�UB�lZ��8l<Y��Qt?!�^�<1���	}/b��r���M2�m*�k���F�X����-0j+d1"�ܴ���F"�k�;,�b��'�dZ��f�V��0T�Q�MD��JA#�#�&������m�wg�ղ7�8G�z������n��� &-Pd�^$+�c���q�W����1z���ҭ�Q/��.�?�`� B�G-��:���D7�*Y���1��RJ��V����ooS���?��$���o@�F���;����˽����������"�G6�w�p��Vվ�Z���HT��¯Y��iY0�%PBŁ��J��E�Fh�Y�T��D�����9��ߺ�n�z-�J��P��`�5��*I�i�<����A ���������eN=�%I��'��n�vi��Oլ�7�/M"l,��˶�5U��cʌi �ϗ�������K��ԇnQ�oB�LD�Cc(�%���i�'��L�A
���a=A�^A�z%W	�{\b����-��)�F��튫�y�y�ؤ�3�W
_�ϐ�˧e��3����K~}{�̗��F�6�Dr)z]�ێ���>�@`�V����I��E�
����[�/��Q��Nhq>s���c@L���[��e�WM��&�K5�,��5�8:f����L�Ze��D1H�Đ�VS��.oYh���m7a"츭;����-��2ޓ�Q ���hׯEgT�O4=�){C<���a	8/�$XTm������R��{��oU*=�w�~��-|��E�p/�1�%dE�~j�}�"X����@L���Z֒��$�)�����w�hT^��.a��:޾+�|3�\}E��J{zߕbnYe�����%����u�d�zY���n7>�a��M��u9،bs��������qe_�ؗ�6ܝ{�bc�X��y���,Q��5����~�*{j��+.�y:P�R�~�����4%�Xc*c���[�?�Fݛd��g�!]"���*
�y^�yDab��?&2ꆁ@ ~���6Y��%SŔ���Zj�j먗:��^k�LX���ΌFd&��(���"ȑ�&4�N�V//wn�X�6��"����p�2җ泽t2�F��D�-�N�R`y�h��C���&��B��J��\�p�a
Г�qJ']"�@Q?#Fܞ�y!ń9�#�ȣ�ܯr�g�`"���2b�6e�N�}eK��sU��*�HC�{\[`JN~�S�[����wR�2�e�I7�&���N�ֻr4�9�|~5��pꕼ���Ld��e����e=�X>ۤ�e�D�~�ڒש�3�>u�Y�iA�x���Ț��Pņ!�f������>��+�-�<-���~�C!�3ud�zLM-E�&��&m,a&�?~���ǭ2�K���sjx�P�Ƭ4�7l_�5#ܽ��}����`�xI@�7$1N=21w'���ik8�a?:��o��)t-s�M��D�F�x��Y�9U�ґ�c�G��*�]n���f����N=܀=�ݡׯut;B��*�:|4a�r�Jv���m�z��d���}M�)A|V��%�ޏ�.dD��(�$G{��C�0�����@c�ckfCm���j�,�q�ؕ��ODW������{�xyʱ��r�t�mVC�Y[[�>�["�����e�rDI�Lx>h�f)b$�
�䄸��P�P	H�Д춵-��JC�@���H��~C�Q�K�2��Y�N�� $�����t$NC�b��i������\����s���N����!4��\����]��K�b��C���;jK�9��e�0aYz٫�/b\
2�D����ܦ�V�	T5J{�d�����"�L{J� E��&�(��m
�I��H��ؑ��_K��5_,s7/���M�*i���-M��n��p�(�F��0f�sM��^���W`	���ܵ(��!f���\̜y}��Y���������.�M���H�y��Z��r���P�3^������×�c���|�U!$��DԄ�]C�����k�Q�T ![��܃H06����5m�v�?��?��4:��{ro''CĨ���_
� !�@�!h���D�*�b=��}���:���v�?��Aod����1�*���p�t�W��6��W�B}���]�Ug�#�@�X$�n{�B����'�����k��Q��L>hkJ��Ǜ]��eљ�.���?�ޗ�ds�:���,�V��|�cǻ@�0ٖjT��&�L��ɆQ5[������ F	8�:޲��~�"Ĳ�HEnFu7��%&�I� L�@�(M:��S����W#��A�h�W�b���M�$D��sM�["[i6f{�I�ZkLo���H}��`^�Ĳ<�#�M�h�b:Ҷ�WH+c湕@�L�Dn�K�m�٥�����|(����	=A�Ġؿ��_�k���DX��`�p��9��[S1�7�Ǳ�:֛�^�.�|Tu��센v	d���~��� �|�+�_|h0ڹM\t�!��Fex"����5HO�(�~;1`��M¢�A8��L\�y�����>)���yg�3Te�Cu���nЅ����ں{n���#�Թ��q��Î��h�=�>Ky�X&�h�W����cIb�ƻ�J� ��"���`8��m�(i.0A(�@j��������vͺ/�+8�0�$���a�M���3Qڪ��a��t�/1�i];W�iVy�jS�&����E1��*�NU�2����.�����|�E��,%$�6����X�^�G@L��sU����ep>�T��+ڊ��/�O����!f�J�Q�g��c�W�UVp��s�N�ׁ�|�(}��`q�����C,^�د�<ܫy��?�t}��7W㟲~^֢���{������>�8����DLR�*�ΟTs|���,{�w�Ͷ�TZ��]��@���q���F�!��h��^/��߽��k�c�$����[GfNS%��,��_���b�Zj�т�4�$�Q�����j��>��?��}͈�lDk��)����|~���0�uob:���.�������[���K��� l:���v=��mۃlN��2Z�k�>����d�v:��c��GU�t��j��]c��	�-7B�M7����?C���pl"�yK��QkM��jO�F�G� �'1b�=�I�8A(a	��O��to����yxZ��5n�o�h�����d��)P��+���|mu?<�Q]XJ��#��b��$�V!U%1k��	�ݻ��lL�`�3?�,ME=>>B����;�#��.����U?qG���c��/��������������Z.kr�*!��$WE�X�[��ۉ���qm�oa��n��[���']�I�AYϻTй��WR_�*	Whuw[�#`;�`:��Ѹ�'p��Lu�9����;&�
�x���F݈�����J����$9��]�$����Z�A^n�il�0~��0s�G5�i�ʻ�y�ϯw�k8�F &��[��n<��M9�s���cQ��(\��0-ڣ.o�9q��(7mh��,0,�!�KաM%�0�-���$���j�Xv�܋S֪��w�z]VQw�9�ʧ�U�p��O�U<]٘WR�w�4ef�'���4Zpo���J�?,c�]�gX��{��>��}#��T��7���
�LV B��%0V��?�j3!>�D���a�k_c�eHs?v�g�O�&��7�$z)�B;��T�������~����I��k��J�Iݎn ��xa���c`F������m+�A��|%\v�d��5F+R���w<���t�"���\�{>@]Җ�!p�\ť�
#oC@��f���3p��B��L�L��d��i'�l�J����ٝ�d�X��G��H��$PMr�69��,1`���Q  ��������oO��9�p��8z$�^l�:�}*K*��{�߷��?��6��ǿ2��:�~56�D�8t��[�N�b���a�2�9@��
��H�@4V�T���7����^�W$�̢t�&�����_�
1\���1��3�xt�Q?�D�W���r���p&(FO..&��9�z)�!>��0F�}uɺ?�?�o*E_�{���1;ܫq��cG,��,���R��`�XII9���a[���-泤eL�K$)$Yl�v�&�PR���*7G��W��F%`{��whr6T��q�0��T������e�+/�~M�D�Ғ�ko�eTb(�RM�ț䟿N��F�]2WK�d��]��3`l_{E�r	y�C�;L�p�����m��FT� -!�7�"�n�_��ַ�h�E^ΨX/|������2��������Q"豞��%:
�)��S�Q9����<�~�*Z���M�	6�=��_B�����͝�ۉ�4�/�Ҭ3WR������7�@��VE��?@��ܖKq��5Y�t�:�<	��h�F�0���&��?��XG���GT~��w���Y����w�?�~z��l�_M����ۏ{�O��^lbVBt_�;a����/�B]~�HG�>�	w7`"���ϭ:��[���j׭�+���׫���紋����3�4�������<���*�,`��_j�z�6m�u�,�q����
x���P�+m��r���<���*M`:���f��D���e!]/>h\���I��/vO��Y�������BvK)؎��Y�΂�C��M�]jgf^����W+:fM.Ic����p�a�_�[��8�}��  ��j#����7� I�[�*I����L"⣣#�#fU&��^dMB���L�*>�L��L��ZX)��N��|hjĎ����E�4?�C��.TO���ȘCm�-F�0Ϋ�)��]�C�6y<g>ĠPϷ�{l�MW��㠶2��w�$�Ƥ_�+�88��V4�V#Z�2��TʢT��U꒤6��a��7�8�� ���ˉ_5�$�!:=Zv�_w�T]KΉ���_	Ձ�hj�k	X��K.z�T<���;Ey��Ϭ�귍/o�ȡV��0���^���\V�f�krg�b��t���aR�����D��ڡf�.z����@���j*d�Y�h�@1QnBvs���HO�����s�+F~�Јj`����8�L?����@Щ +����#��+�dP�x���i��B[��IB��8�{���纞"�/G�ɵo��K>�1�i���P8�N����eͷ|�T���'�Ef�f�֎��|�7A ��7�����t�$���x�"U�:�#�������~��μ����&���}Q��g��;��*���$�VVP�aݝ��xz��<w>��ﶌ��Y���,����b�jCz���+���+B�q�tNU� ��z����]Ǧ�6��`F��d;��������xٗs���}�*i��W󥹸N���Fd2�f�D�F�B(��O{w/���{�!�vb��k �[�zW8�7��?b���u=,?�D=�8�V�K��l�K��}�] 9P�PIZ�8{h�y%F����^�UcZ��E�����瀚���i<�|܋3k�h��C͙>8Ѓ���PZh>�B:iu{�g�% ӈ�#�I�4�_}�����3���8��ҵ��ǫ(��E>a7Kd��N��i>��cX�r���}X�(Os�\��{���lH�zA�	;Z��L�šE_＝�Ma�;����n�ʦvx��o�űD�
w�i�Ǟ`ԁ�vw����}�JЁ�P�ջ�S�$����:��S��̪�����[ ����5���{qkq)�Pܡ�kJpww)Z�%-��ݝ�,����{�o�f�@&���=g�yvՇ��ً�ӡ�A>:.��\i-ч�������6�~�>�|#��B�u�{���e��u��~a[�������X�Kpmwi�P@�<�_=5]����T���%�Z%�h'a��+Sk{,�t�>��z21�q��5]D���B�/&v����g�D�|U7\R,�S������|���';��
�R"�{8 �z��4���z�~j��B�^�-ϊ�f����r�g+� :�NL鱸�G��h�q)ܳ���k,��m�C󂧺������mҏ�P�`Ņ�m @-�q�T;@k��P��B����u�O� ��/�#���%@ɻ:ߖ]+Y�b @��£�
Tc��Ƹ%́�q�r7�h?����e�:�dP�7ֵ�u���{��Ġ����:��OҤO�$}d���-GF��]�u���R@�W�����wZ��PB�3F�m�?$&��^�"=��* ��?��!�ġ� /�,T����:���&���:Ǜ���]� {Lç���@_�a���P[&�쨳IQ!iȸ��?=!��ݪ�eJ�n4����?J 'YY����_<Yxb�bvSu3��MW!�:�]�W��X�[VP�E=\��f\.(n�o�+iMdy��F����X(�a+ÑU_x˔oR�f2�EAj�%�<UH�Ǔ_!o��$;�����Zi~0����'� p��%0�X�'-2jo�_�&M~4�#ʢK�o���L҇#y׻�Kx1u-Ͻ��I��1�^n��mt���6�solQ^!���WS_+n$���T���|%6�)'�f�:b.!�q�2�ٰ/;>;��Z3S�~��3a���M�b�����xLV���#%���ZD\O6mmm�+;=�N͞�*�L�e��K�oc�a�Q&�]���n�����N�L#|����p��beh���)�7I봅��g�;^��QB�K�a=N��}�}c��n����!5[�>YMw$�@T)�~M��Ǔ��t{W%��&5<o\V�;?Op��˱lFC_^V����bk���)�o�Yi��������a�ҭ[���6�y]��VL@d~��4'�h��\���4 ˮ������f��k��*� (rI���ș�H[?4�%�k�.b�q��9@�,�$$Db�Ͷ����S���c���?���x�F�B�4hs��[��b��c��fA<lZe�]D�s� N%*����\��a���3��-2�O&x����F�bj��XbA�{�ի������G�c�}�O��(�J�F*��=�������^�q��毋����:j4�m�߼�/=����w�/1�w�
��7�J�`[��b�8݊���\v<pW1G�\�E��o�`�v�eA_����L[�h�8{�W�p��?�pt���d���@�3�'@a
�5���<��	1d6.F�&ԨMYt|��ס�5y��6��<�Kͣ������+mF��&$֖s�~�?Tl�u�͘ޅ�U��dj�ߨQ��v�T�{վ��;�`J[�;!3"nB@� ����E��f��U��G�AA!�j/�Ȍ�f�5-�g�n�"}Cң��7-�R�/?(��/UfgcUt��,V��}���?h��~y�����&�
�qC�2�4�9�~t&5.߹1�q�%ϨLY]�����$��p!�wc��Ǉ��+���U#pA���Ô{�2g�0(?U=����ވ��4x�[�t��<�s����v�,حLH�s<��vv���;�GM1�晭��	���#�0H_�Lj�ޖ}T��`S[�	�\���~�6���_8������R��	Q��f�Z��Q�/d��1����7�}�-�\/K���$
x�T�=���i��ϧ;�Y�y�e��򰆽f�W
M�q��;�_V?�'���q|S�F=9����X򾇺ެ�Pzi]����:)��~�_3�#�q�fX�5����� �U�k�����*�N͂�d�H�#����H���K��&�I�����+��W9N�W�
��ڻ$m��6
T�����t_�K�V;m˔��3OV�?�#�y��-	җ�c�-q>���8%[�5����հ5�񦕷���Ŧ�@���[�?0�呴T	���)�d[�E����NE��Yz9�_k(���m�^�*�@$�҃����s*K�ʁ��³M+K�Ll�R8�3�W�~��}�X�G��k|C��mAq��5���@)4�[L��U&�z��#F��aJ=ת�L��병O	:�[�8]�m��Ǹ��f;����ϪY�nN����ݵ������-)�H���������-;,2�\�w1�YJGG'7B�,g�[�_�{�D��YT�#���<飂��H�Wu�N������z�`kRO^(�`g�#��6� ��\o�]�ջ-
�k(Ǹ��=�-1H���\G~��*����+C�{�W3m
��#�\N��C��t�[�U�1<)$3�f����\��y%Ve�絫�N�H���OW�J�6��izf�x��V;o�/� ����|nl�7_+^׬��n����)�ՃW��8򥏂�ҍiE0��`#	�غ�^k��a7���	{��=n"�����nK/m0����k�^�!q��[7�)J�& /F����TF�ղ��p#n1_�Ga���h�2̃]�b�\)ac�m�Śh�Z����H�@���G�beת:��Շ�@U�)X�x�YUF*����Eh��B밶=���=�(�N�E�������L-!Td
c�5V͞Yg�3��@�|Ar����o�7����uy�����R(��^$1��K����~����˥�:R��EUv�ǉ!3Z�����9}��7�>�Z�FR��s��s�C)#���~�m闆{]Eq;�A1���z�;n�Q���b2���A�PV+���/�͏N.�Ə�o4�OJ0Q{�W�	��/6��]�5�C�t����,V�2�x88�1B��0}��Y���z���P;������Kp�w�D�_v0g<���})��Gv`�YvXT�HL����u�#��$'"؊K���C������=� s��?�;U��Vّ�|���m�����{y�~<�k�S��b�*��f��-`
Y!\�gq!������F���BTID��Q\3j�;���Ⲫ>���߆0�7X풞[=�7ܴ��!�zRsF����_өw�V|��Y����Zʂ��D��Vg�N�yHM�g�ʡ�#޺czԪ���*tg��'�_)�pQ\C=��K� ;�zъB��j`D��R�^D:E7r�R-q��K�}a��ՋA��q��vV`�<3��ǩ ۷��I��G�����b�����q�17�]��a�p���qlVW��/ED�x�ڴC�p�sn���2���`85��g�p�6ᴏ4; ��[��C.�w�v�
��Y�QtQD�T6���@�2��Cy�@�e��$JGn���)~�ἕ�=���p㸭�Iq����M1��E��CGۄ����M�g���蝡\ ��5"�}i<�R�9��[�nHĂH}���1���{���FiYe��a�M�Nf�CꎓC#&b��z�&ܡ��šZ�'|I��6����L\�Yd>L@|v���x+��xN��Ɩ��}�kOW�h��d�> �׿�ϸ<�4��8�=�'�n�|���	$`/��z*v��m���#��O.��a�E$$R�v(X�#i~tz��Z_�8pF�I�e��D�N�#G��{9�Nת�\s�&߄S�<��r�R�����}�`Z<�nò�2]���#��|>԰;Z�哮�T�R!~ʭ�'��x�Yԧ?2Ɋ��8^o`(�,hz����ƾ��w�NsF���,�7q៖cS�Y{���� :qoٟ�4<���8�D>Б�U�Q�����H��:g^R������"����)�3�r�wԙ�k�/��0�����0̮���g#팱�-�I�#�A��E-�C��xp�F|z�r�IBv�t� n'-���pc��&knYӊ-���)�4)�
7KM ��,nE�]�|���@(2�&��hH��p��x�O,��;�v3�}���|�e�G����Yr��?��n�}�br���C&b����\�����\H�	Uz���ӿa{5X�T�1�玮<��N!��\�ђ���P�;d`��G�J�Kj{�c6N=��C��`�,g�����B����[�B�f]�ն1�̑�z���˶&2��Q��!K�������⛿$�\�0������8��Ń����P{���I<��|R�"��R�� �^�>��
��qgnT��a������[Q���l>�6�� }��u{�.Ζ��m76����kvJ�;(�QWzg8� �""�F=���云���^ZQ~"K�/��	���d@���
�QGX_^e�`#1�BL5��_�ho��M��d6k�z�J�	&��N�o��eƭ���$���i�'�t캊,�D[�� �V�:*�T)J��%�uR����sP��j��-d\���t涞 �2;ӏ�������9�����u�Vv�^� ��}��R��Ŷ�����"�|��g�;V�9�ȧ?�+�N�r(agL�ǘ�A�+cO�\�R�h�����6Em�������c�K ��Γ�7�LKY(E��z�9�%�]~��G��j�w۫X���k嵺xc\\U���ى�����z��P�c��)b2�N�Z�zN�-u2��A�m�|���Mn�݈[��1����r� ������$���MFOꒄI���U��+NS�,0��N�ER�s<��4�5���G�)__�E�	C�>4(��e�!(�_�O�7�DG��$��>���|$4.�q�=�^�w�Wl��j�$���	�9�?xUk)�8�t���0Z��BwN����'�P�GOuc#vvۅB�M2���I���D�1����%qv�-$�&��ӝ�9�?�I�N{n�U��3T���ǈ?�&>^�d�En&�Ϗ�c�Fd	#k���덴Y�w.��A_m5C?�%@8U(ϐ�c%%:���ٰr<���9{�ЪSF���)6���<C�PΫ59�3��w�b�f",8�	�k�ǉ_�
#k�CaӤ�c�&�GP�{C%����������ڔ���쉚�ĦgR
�̽���h����P�7��a�,X��/f��'w(,�Q�_�
B�	����v���MY�j䘙�_�``��N$�Ig�2m�ǖ�@�B�)��|z%K}��70�?���H����9P^��zI��І#����{�#v���vE+���R�8z��sxff,\�dco��z9򧐷k7�&������Z�N�JWK���?�y����4���8�HC琚FԫD|3el����d`Ѫ��1���tw������R�����l��*�s��]L��� �'c�� ��y|M�%��B�Zߢ,w��%'�à\��߶%}�O*7H�J^_~� �@�x�^eɗB�	j ���A������{�{yn��L,N�X����F�{M�%$�k%\��kx��9��<[�>��5�8OW�,��k�cyܥ�տ�*i�����w�۷Ǟ���pO��G��DR6ז�~�����Jl����5t�"h�����=g�1�Ỳ��$�.�����WYMm��]�n{��_�ǅR��?��,Q_GbL��JO����]�+n���V]�L��r_����b�ŕ<f� ,!�dǏ<t'uV���ڡo1�ߕ8��ё���L����Żk'^�*����m�߾*D�c�3�
x1y8L�M��MH �E�=�l)Q�ż�Q��R�b�vL��(Y�d����7�T#֒:�h����9�8�[.*98ir,am
��4U)r�)1`�"HL�u���[k�K���%���w����o������Ff���,���ʻ��{�Pu*�d/��g_�n��@ه[�;��,�gC��K��"��Y�U�vu9F�ʵ�~t�4/��K�B!z�_i5/T�(�������U�G���(<[hÙ|�fw����Fh<ϿGv�]u�����Q3F���cЊ�������P~j4w�:�;`k1� �	��'�WY������(��C��n��f��t+�3����J�0��(,��C�rSe���s��.NV�/�/tU�>�P����禱�~ݱ�"�� Z��s�;�۰�f�|s�]����"�i=�J��5��@+�h���%�Z���ۦ:��}hPА��w��K%rj��,��2�(vjLzό�޶Z�lv_1�}�g���Yf����yߔ�6�Wt���!y��0*p�DV��w<��-�;�C�y��!�=;��4�䭞���&j�g�smޗ�r�zA���ףծ�BV��y��}�+r�l�9�ס����&2	2��*�;J7|ОJ�^�题�)�Ņ�����f�75�D�S��J��#��i\��8<o��0vO�b��D��a95d*Mj���Q8���/	ur2pm���o���;����bZq�K�Oʕ2�v
�;�}z��;y��@D#����z('����s�|��`��IR��z�k�m*��lTb����c^�?���K5�G����Q#��M���k�,�Ctt�0����K_�vTX��y-~�n uT��(Oȓ%Cn���{`�w�|HU�O�>�>�������l�uޑ���R�!ڤ�
�p[�*̋a�y��0���I**q	����ݪ�B��>]��J�Y&�\?̯��8x��ޫ���jH�Jcǳ���S��w���\t�%��Xv���	ؤ�Zk���h�� ��n��B�y-�l��G�R��fUH.�+���J:,�=�2A3��Q�y�Dag��;�a#	f��B�kn9�[L�fܝHڮ��6�Rn\����=����^]N��ON�z�	(���R�֚�x��>���m�� j��р�_:�����|ܹw�zTw��`d��٥�[�[�}p��bo�r�Ţ
A�� �_����+�{%��K�%I�>��z�'��>��H��L��vİ��O܀Y�]�� �]���d�~���A��uEԹI5�8o
ư�d3���@���X7̡F��!�s��3��#��[�h��p@����O$�"�zK�Y$�N&�A�%�[@�Pl*����1j�*V��ݿ�ݘ�b;�����;O�[�]�h�J�k������7�AT�:4b�uX%���<�,:�r����_���u��Ц.���+�ѳ��lq�T/��=����ߌ�꬚y�rȲ^�+�@�kUm;1;�?��4�
�G=�/Ub���i�I\�7��� �mx�
�O>Li}�A7Y�֕���V�z��x��.��$1i@J��#�S#�!�Ϳ�J�=����̹iJ҉e$�SI��_Bޒ����Wc�M��-Y�������?� [N�.Eu��B���}����3�[vl�7�ߞ���q��/��foVJ��q�|Up/�'�& ��nO�����{���2RF������\g���C�uB�����M�3���>3�|/��O�A˃��������B�>!������l��YA/f6�{�3t�k}P�}��x�n�G�/Șo�~�%�@���叇#lw����]��|�'�]�ln����p6�����a�3���,���8-�t������!�"���@TQ����Ԩ���uL���9R\D
�(i�ǣ�ܟj���Co�5ҁ��!,��l��������:���m�$�����v�r�,��������V+�hu����5�a�WY��&=ۖ!\����3��`�f�jX�Ϳ��9��w��H�T0�'9��*u�JX�z�^�����<��eХ�٫�مg�A���&x�4K�A�Ӽ�I��N%ۿ/��ĆS� �i��l�9=��
��gT\$��,m�G>����Li�Ù���՜hL�O���V�E~l�1�}�� _�i�B!�/��M�Ԇ'
�4�3�x]��C�evڲgdY8/MኞNu���f;7��d�k,%Ql��	����ӐA��ܲ�ё��4
����p:jQ���\=߼�c�8�q�Z\��	�;v�f��؀=W*ms�"�Z~�s�Uםro��*���1aeC���X�� ��E���&��sl�o|.�D�ʌi�5���v0�7�ϻ,�����.^�XyG�i�g?Ix�]�5��R�\<�:��ԃ��Z!�
\"|a�6TB��>�u..����|�,bS��A%�Zc>~`�.�j!�p0En��_�j�����,�:�w�w}�M�S}�D"�8�g2�	f��0Mz�T�s����b ��䫅��'f�?��
ِ�O�S3�Gm7��W��ߩ�� �G�O���dn�2�́ATF�W��ZחwH6y@���L�FUp�$�?K�~W6p ����P\SM����v�՜x[:��L-��8�2PW[���D˼(3���S�:� �3�R�y�l�9����1�����l����Jw}�ne�mS��	b��0Ŝ��܀D�.��T��w��c�,R#ng�VI37=��Dzi�gtʦ�`��$(���D���Q����A��68��i��-���9*ĵ_�ݩ�	~.�D���<`��A<�Z�[ً����S�{g�&~�c�Me��w��Fv>� a��7�4@lIi\\ ���X�SV��Ͷ�zN٣���,�̄6@��=e<ZVW�YF:%�AT��9�i�(�g�z$Fa�*M�qP{�\�@�$�j#��ô�oN>��IO��sk~,T샴?P���Z��k`<S��Yo�G����b�S�Yئ6MZ+�0=7���J�GYĹ���]g�y�
X��Vվ�]�4��j����m�t3����01(��|�~��d> ş�0�dp�;�OU��17�ă_��`���(��~���kμ��Ac)E�y�x�.}G?s�:-SEQ�`�_������Vө��Z���te������̝=�͋���8�����]����W�u{�ƻV����G����%f����2l��}�#ΣVbv9�󵈋;.�l9���E������%9NگC,:T���7�d^�w���k�*ͺ�#�5�����>�oLd��c4�'�՟J��D��|�$��4����̌V���+�F�B�4��q{�o���g���5悃ˋǩA�	�Dq���aF����b-c�b��/ʿ�p��g<J�\őe�9�C,���Kf#�������׎��d�h���E���suIh�X��|�pUlqqr�@�Y�A5��ʡ���T��I��{b��lC�S��m���g���.�c
�J�\�85�f�����q�h�iz
����]���L�W��/ҽ�ĘUsjN3�	 �E�j��v��ǲ�ҩ�-z����|�11n1�g?22���T�?j0�&!���L�fF
��8:���F$Y��������t�����੠���C�ړ1J�?���7=���Ό�L���9�$�"J�}ת��QD���ʻ8X��+���n�TW�r���0����:Cݺ�������P6F�hr�DU}Ԏ��b��k�Y�Z�*۟�r/A����}�	��[���c-���
7p �%+�aE:Ψi�_�s�I�r-��
h|�=�B�r,WƏ]d:5�8�����w׾�y����7r�����:�\�-�0�)��$��K����j�����<�)�t��<����<��y�M��Z� ���$���?I:bĚ~����^����.[��'�sq��=#�o�r�V|UV�ڤl-k���G�V�_�f�D�q���j�+W�蠮z��l=!&��L��@�?Q?��C�9K�����s��L����Y����<�Ǩ�wF���\y�f�(M媂՚K�B��3@�(=K�Ҝ���S��w�R"���uY���Aa��8�8�����*�a�d@+q����%lR>�	��������� l@���3!�B.�]6�Ԯ��eI3R�p���ޒޭ���  �9�x\N�H��x=�)�Hn��o����lc��u45C,���&��~��cqXw�z�zQ7h%�
��w�@C�Xo����7�~�C)y���Zq�]0�k�	l���������zN���Z�''��4r�$�\V�C�6���'����t��N'?���Y�+���C�ٌy'@�(�`�]����n�����$+T�`/PG���c��u9ca�^[CCc�0^�σ��韽X#�>c$c�Ȑ.�r�{u��c���b���|�ujTqMmMnELe:�@��p����i(Ԑ�9-�t��>YG�IJ*y�� ����K��"�6�(���!�IJn$�o����|�e��o]��ܟU>Hh����#�o9����g����un�vs�	i���C�i]���d��]�r�,v��~`f������u����G��|���
?'��k�=��������)�bHTI�. _OC�6E����Z뫵���4���}�,P=b�e�=:b��y* ��8�n�Щ3���s����x����yl��4������7_I 	[�2�����:mv����o|rm�����w�
�������Lv�c����	J�o��w.�)�w�=�5���Kk� )B�}�g������3Dw����
_��D5�q�)X q��H�َ؎z�2a�Ҍ����?�'��Scm��
�i��`�V)���}�lfOc�&$�5��a?e�h��!L+��MĿ7J���׻��ݐ�G�L=��2b��_���8��(9e ��b���f��ׂC[��0�r������v�M�X?�t2$_�y�"� You����s�\4��\���榿��8�fe���"�(�W��<=������ml�io�zI�9E4�"�|�	{��M��Az��1}�1��5��mơl�jv>�}�K��#�q�N���])�6�����D�� ?�����������=���EG����]�VX�p���*#ti�C����ON�N�}�٪���t�؜�`m���:٤���1�N�LT��a݇�e��s�IO�>���aQ��pC�-�w݌��-VS[����~+x[R� P���lix�&ix֦ř�B%5�l������e��cG~����z	����w�+���R�?� &��@s;X�w�1���c�
:7k��t/Me��Y����{�t�RQ���4np#6��ȳj��QU��xޢʆ�[�oa�qE{���_�M�O�P.�u3i����'���}b{G����b��n���Q|91�^W���I�I�����ާ}Dë8�'Q�J���Rd%!!�$�t���+"�ݎ�&��f#c������LV�*C��9�X�O�9���3�!�w����l7�bGW��:�R���y`�)����Q�]��$?���5>
r�����M��TN/8��+�����N��-���l��a��X1p�e�^G2E�5���t��ިT翇�-dh�v�K]���A���{�iǚћ��ޜ�0��c���ۭ���^�~��9���W&sC�ӎ�X��j pl�k��� 4��AO/�i�&�y&@S���	��� �	8be-��w�'Lԃ���M�~���H߲W4r�l̍������:����{ai,݋-�m{#-D��V	=�2	�Bv���M�_����M[	sCA�T�D��a>��A��}}�yI>����γ�%���S҂�i��	�z	�X���ςM)N���G��>�g�=ۜ���^E�h�oj.8����>�2˒������E>.P�|Ssh']�}����1�u"8r�����ʬ4M�4痃lam�tV�;�[�9���6橡����<�9�0��{�lfe��;����<ԥ\�&a�/����8��Ⱦqg�'\1Ps��`��)Fl�0-��&��;�$АE;B��΅$B�TY���#L�hiM1v,w�v][�{ ���6�Ö�B6����BV�PʅK�ۼ��W�sBH�'|ָQ�u]?��e���P��o���MZM�c�Ӥ��W;��E�xg�WI����r������Ɋ��Q�Y���))N��M���	"YB4�hi=a���JJ����O*��~���t����z�)d;��X�s ap_�U�UwG9+8����2߰c4�opru��D5���E���"���	`��ky�"��<ݴ�&����+:����\��ؐ��g��)�X949�����ڼ�IF�mWw
����N?�4�M��v�b���t�N����_��֭��W(4�z-#@����}���Q�Pt[�%��zڃ�8%ϵ^f�h����&��|:	[v�G�F�}���XG&.lI�0�R\G�f�{�}2�_�߾}�Y�3b<$A�2�p��H8wXi�˄d�9���N�K�~,ϻ$�mw�Q���~h�ӣ���-���N
tƴ�_^��������?���^���U�y�r{2���=�a���r��qO8�|����� ���a����o�!����7�J���{ay�T���Š�||W����F����4r�2�)�{־����"姯��:+���!���~ E��-�-�7Yr�ʧ���F����%9�ϵ��Ɏl%�B�ٷVu�ƽ1]��T�$R�Ĉ��m;|�/o��>�4���T�	z�|��RXX(�#�i�ьF��t���B���"�k���`��۱��u!ҕƳ����FP,��?���ܫu���.���|��+eJӈ��&�A���v���,i>=�e������O���i�Em*�^�hMV!�%�4g>;�!�x�*s$�Fȓ��[ʁ�bq�K�������� �UQ~�a��\L�$����~лSM��)g�R�����y�H�BX
��3|%�!���x\P����(Y*Wr���#8�xУ�#GKvc,KvRH=�J����(���J7
/���v�'����M�p���Dyp�sI����V�gQT��H�¨���ԣ��y�[�/:�h����	o7ܾS
S׋��b-�t{fQJ�"��W]&%v=a�U�2�ý�e�,3)�C�i��A��]�0^6�M���*�]�E��������;ڽ6���]���r6v��{9���Xh@�>�5���Jb̕7 a���J?ͮ,�%ē{���Q%�x�!�x��?G��*����{�Y�^�ՖJ�XpBg��f���pa@�D��9��RB�KE�V/��D�!(tJ��nQ;��
s1 ����-�B��+��#�8�p��6�"F������aQ��7�#{i�R�G<�ixa��{T$Β��J��"��0쳔H���y�y-��E���!	f�?�9ԓ9�����3}���󯔍�G��P(����q,}�p�
I���9�n#�N�]TdO��_�z�v->z+�k̔�ofTl�da(�UƉ���Hwc6$T��g�R���t����T�����ow����ߦ�*,���\����{��!��r��p�^�,.
����R�bk��� @�WL���:��Ǹz�鐷�Q�:�����7&91~9l��v���Umm���M�~(�� I�V�-�#V��B��䥖<�'n� ����NA����m~�J�0B���p���`}zRUmq�M�s2~a��8rUT�r�/�c�T"���k�<�l�R�]���y=��23k�aYGo:ƾ�TT�s��Ė�Q�/H����iV3U�ᘘ�f���1nbbAo�A�� Gz������W[������#1�V�� �gٔu�e����I=����2fm��8
a5�4d�����6 mR)��_[�:4��<�qI:�o���Jlb��uk�k[��0�J��4%�����?@nM;u��x�%砩�M�p�.bu�q-GS�r��������D�g��i���f��^z5������3��O��\��yb���w_�;�Aٷ���ӓи��`T��A��}���G�$�&���u;ݿ:1Z��2�`�?$+��C�f�_�H��4�'�)��"2�b� 3��`:y��R���;p�Se��q~L��%qۆ���w�&L5�1'J��n�u?z��]RTV���7K��]z�Fg�IoyQM��'*���?����Rȏs��n��U:�>�x���*Y��ъr.��2��g/�Ύ"�Hl��e�Zp{��@!_��sP['kI���q"~�c�꽥;fLV���4Q	�S�.E�wq_՗��߀�R��qY���8z{p����kc�#��ԋ8�lF�d��Ǫ}�FW7�O��m����-$����7��U���I9(@=K�����܀�&�0n�����s��t޹'J�A`U���l$[��<^:��)2Ǐ���~�A,A遁��I��p⩈"��4[��F���g3M]>���H����sf��6.�%z0�`���y�'��"E�B|��� �����@���{�/�@59!u��_��)�C�y.y���zY�xO|e�����P��+��	E������Q��C���%ũGtU, 0w[^^^dd�?��Ӷ/�)�l/#L�".)iF��@�vۗ}Ƈ-M"U��p6��x�g�;���̻ھW���o�^�� ���e�T�8V���I<����vjy��,��~�e��ߤ�	��a	��6c�u~r�v��>��j���$Sm[��D�<�h:�hnwf�l����+u���k3q����a۝�r�E�8�� " ���+z#��y��}t��drP`���^ ��|���p�ij���a(����~
�s�f]$Zf»��R�a?Gbe�m������d9�mb�7:�`	1{�
���ge?�q��T�en�;6"����H��A�ڹ�E�a��O��6�6%-�Z�q���m�ʼ�����5h�8
�C!���6}�~~/�_�=^	�πږGo���cWBs��g�}x㚥bGw�p�{�kG�ϰ{����#%��&xiCG�QZR�o<�4p�z�߷�fPDs4}����\��p�}V���!�2��q&!������c�51a�{�^<��\P~)�;Z�\��T�;�7"��J$�����A'�uԚ���w��+������ ��T���Z�o��6k���V�m��a�.���Oe��*Gv(��m�;�NZ B{f�IL�M5
�K+���_CP��GYM/���Y���5�A�p��9�2���,C˕];H����sa��V;+��č5y�T�R2D<��9����Rֈ۳G{l�in�?��YYY`�J�(P�S<¾��������PFgE������p紉3���;gu%o�F��B� ѡ3�<�ٴ�f��iPم��]�#]���뱈.N��7L��uR�����?QH�͑g��faW0>��$M5N�����P��AQ�`��+��ΰ���s� ��]�}
������>�fFs+̮3��]�p&navz����|r��h��.��\����

�i��BLNګ�z�Zgf	ܰ��è�mѬ��6��&���rs{J�h�kT�9`��<3F��Y3��2����!��V`�;�T����2x��L��Q���f���ڴ�чn�!RN��w(K���`ܞ�%.�,�e���]�Ȥ֟i關q�_6��@��_���X�2���N��;�+f�S~Ȳ�E����g��؜<��sǐ�8�� �Q���i�Ii��	���)�U�4��(����-Va�7�yG���W����ĎS���<��Z�����j.��m<ߥX��O���d���.z0���չ��[���^~6��z	���Gm�s���V����6
.���Vd�@y�,\���g� 2�t�$�12��J��o�O_�7�4��\η�f!�6!�����c�6�u��^�Lgy�I3+(�	��P����-�Q��L
>�96�1K뼱AöEw2��L�\���t��A`��8�T0��PK�I������:�_bđ>�`�O�Wq�=Bhi�C����;i֨�"Lp�@Fn�q�P:��Z�����Uܬv���bw1�<��[�4��pFRLp�qd�G�y��ж�*��zH�ٺIn̚y3Q���i�֛�<ՏZ����p瀕�|j�B���1�z���8.��:n�Ȣ]߂yUX��ñ������l�u�[��61�j)����;�ST=����	;���w##sϬ,n.�/!���D3S�Ӎ�v��������$�4	�
��+bNG��D����+Z��a&�#�?2�.j�9��
5K���fA)�m��մ��b����O^�a�̈Ƨ�)����Ւ���أ\�͊�ݠ���L�}V/����R�����46�]i����%�;z ��(o��a�&\�И���hљPJ&�w^*<ĸ}�BRKKK!�����$���֗^7XY�rN���wY����Bحu�7 �!�w٠�t�K��.-Q���H3B�N�Qc�[��AD�0|�� ��F"�z-��£YL�5eE�É:�y8!|}iڻ����L�s�z�c�:Z���eAg擟v�޷u�����O_�v�}M)������w(P�X� ����
�X!�J��Z,�]��~���f��2�d��=��wם���`snڹ	�;�t�M���|G�pN�T<��U&QLY�Qn�2�9[�_v ���upበtC.���*��u����Ȗ̯X�B6��������V��\<v(�?|0�ܖ�r?emr�:����1��AR��8��ܩ���OVPo�Qg��~29��2�\!�l��	Pe�"�hn��у�ќ{q��稡;i�,�[�Y������+�� ���O����6z����Ӷ6�{�nٿ��K�gu�ӂ�?Q'~�N��3�"3�m'���o�t��(�b�!������ܑh�����^��5�6"���E-u�E�,c����+���P��3�f�����m��W+�$���M9�ݭ2.��T 5��>-V���|;=P/�l���(TG�Q3
�nl���E�6�Im�&H�!~��{�Dl���&~����(Gh�5���i�i��Lz�����%)W��q�k�C{��1mITkwjz���Ժ���̧�D�m�FmT���!g�6sMC!�DD��>�-��Ww8!�leVG�fLX�o��D%���+�C�o��p�LBJj|�ZX�AY����us���o�����צ�Ǯ`����_}E�����CGr촹.ς	���<��i
�kU1���x���1�����95y��@��7UF���N7g3 *w���C-crlX�گ�2��n������j�+Wz������qf����8����a���$$s�I;0��;ȶ�Cm	�+>��[�{���`o`�C�J��G�=?�+fd�[�T/Х��sݘ��ZʣV�f�5�*`&������ԴC6���p�A��2�hE�)l��@���3ؘ�ׄ�Y�~�_�_����U����M�Zsek���&w���:�/��N���x�bf>�Oʹ��^�+���?d�]p��=γ���)��-�ǫY��=�5��gf�Xҗ��Jzo���b�t�~=����I��]_%��!d�� �{�i.dF�%��E:w��;=I	�8�ngh���_��D��:#�k���@n�ū��;W�Z��΋)��3�Zm��[.�3^p��۾י|��~�ɣ�hQ��u��8�h��><��&�r:��{ؘ����JL��_�R�9�蟇��Os�"ȈOk#"Z�"�����	Z�H��]�N��#ve�Է���j1�-�.��6V����>(g�.��#�׀�$�Yi\j.��:	��Ϲ�[y�Q4�[���*9�{�(�Z�B3S&���H��b`B]U H��t�mL���B��Xt�T��'��UҒ7\0�5Gzb_	�dud���ך#��6i��	jQ��=�?��������R זOOG�������������l�����c�@���v�+��U���,�m:i�y���q)�#A���1��hɞ�w�Z�z���f��~u	D�m=���N'h��-ى��a����h�����=�P/Y�z�-+�T;Wv��)�g��,��]��
�#S���6h:B��zKwK�9��YGc��|�;��:&���9������!M��{́޽ő��c{${r�3ߧY$ۓ��sV[P�K��Sݖf�W=��Ô���6{V���m���O�*U��Z[r���e��%�Lzyd���r"W���.$8F��q�ٟ����K�wY�ҙ.O���x ��)��V[�/�>��wF�S�?ASV�*<�,�6���ӝ�^�9�;M�Kľvf����H������Iݹj�o��[�~�5l���u������u��mݛb���_���kFIU<�r1b�a�<`��4�����|��j�<U�VB�J8Ҽ�3�dH�U��h1�4F�zӥ���0��B I��!�h��@��6�H5Ԙ����->�*���,]����h_�u:�bu��f��}Tx�oJZ�&J'�{���ӱ��������2y���?�N���ԋV׭���#�Fj�@U���]�+a��\V���0��IɌ��$�ѳ>��@��
Nz�Nׄ��MY]�3%�ߴ�i·hA�fFFK�,�Dd���K7do1��?B�@�Ԏ��}Tx�<����`����f˟�dq!!���!7���\�X��q����3-��m��hA�Z~B�IaR�fR"ҋ2/��T?��)+�b�|����k�>��T;r���lv�B��/���`�����gk��
>��lg<e�Cr��D�V��5��E=��H;��Æ�ME,�%Ӯ�K�@�rmC,S��M��T��U���L���S�N'��㭗��&H?ܸbF�.עqz����nd�t����X�]˭.v���H ��
`1[��t-X��,p�R����K��mc�����h�(�����qZ�������_�0�@����t���rt>�LNL�f���Y����"�i�=��8怴��
�������A�Ԏ|�m�˦}���_� �X�Z���Pf����֦zi�qL=��6�<Bf�	#H��߸?(�����3VC#��~����W�S�4c�_���r��"l7c� w� �)���B��6]��B�O4bzi �4�^V��;90�~^nkb���2R�~%��b��r)��I	ڌ�os�J���M���G��d�/�T��RR�b$���
���e'�爼~��(��)&@��H��"�R�t3E.(��$�-^�&�f�����b׸��9��S�����OE�;�7��������dP��G^Wb��;>>lP]�U'	A�q����߰*�3,o7�C�ۗ��26�$�%��k�9I���?�a�2v�)}������}�������땀N���bG�}�
���`�A9���.D0)[� ���~)�X�/�&Y�s ?�~��+�X����$�)";*�#���lW��7�`�y�:i��U^I9,�S��<�ɒ�p�/^�Xb��'��ns|]jO�0&�$ ��eۖݻ��4���D:��� ����u�u���B�؏����\��^��%#Sdb��Zo#0�G"��k0>�Ƿ�,w��0���s��c����fסdpc�/"����\9�6_T	E���q��3�gU(k����"ϮV���YJZ���2sT�C�|��[�����x���xց�� A�!�y�����9��LFԚ$Kp6.�ޡ$����*y�)R�znIێ��;��ib��v�~�9^t���{�Os3��D�*�$��)#�T`���sF$.�#Z�zW�H����8	=ذ�)�_ �K�?�n���l���\s��r�.c)H��Rﲧa���^��2ig���'��f�ң����e'�;P�їd����v�_���Wv��+���6
�S��&�Q������?�4:P�ΑIEl�	����>X��վ������=��Y�4A/��63����3�*9��C���\�� D �#8f$����
��޵w��\�ztG�)�e ���f�M�P<]*���:���8���m��̊�o��O����1�K��O�q-��i��#U��S����p!���_�Ut�/����̍�"h��!������}p��}�b�Z��'���d)��@��n<3
�~̟�3�ʲ�j}��Uo:�[6�����l��6�O����vB���H!�w�5��s�΃@���.��!t��ￃ<;0��l՝*Wt�S7u|�1�:l.�́axd#�ɢ�&�c�{��?����7�6`V��㚑�����o��8V��q6�W?`��eWd���P���꛺Q�Oħ�����q�0�� T�k�8��{xMk`�@3H������C��ͷ�}���
��-"����CJX����R��X��n����?��mo�b��8��#k+ip~~����}��K�a�QE�s>!�<A��*�_�F�{S��N�9�x��ÿ��s�4��rp/ԙ	ˎ����Zj+�i�Z�����ڒbJb��\&ݜ���X:��agG�E=ݗ���z��f<��~�I���mc~�"��������ZIh��%�w�zp�_�>t��K�����A��۪��T7���ʹ@�������cF�nݥ��d�^%�I�K�l^�|��D��d�U�BZ��:�|�[w�A���Y"�q�H�5Kr�����t2���c���pQ�2_��n�턘7#ݶruu(��v�ǉ����o_P����%��D���:n�8�p_2(k*��w\�I��_E��A' �矛D�:y����+b9��[�gLFG�U�4S���!�n��M���A�SY�����KǚO?���ki`���s���Xg�@C�������8��Up)E�ӵrhp�J9A�4�����_t��6�M+{'{����o���&Ã����6;�X���5��I
�c����ik/�ȓXdY��I����8���Cz����� ~�Ҽ�Q�N6��j(�D�~ن�4��Ґ7_O�/��{��ap��\-v�=4ۚ4��Z%�}�`Jw�����\�W�s~��S�frٌ=��Zn��q��.���6���b���QRn�?�p��>�0n�����bj�q~�
S��^1���l=��D`s�����&x7�%ν.�
���4y|N~!��4�� ��M��QeoQ�p~�{Alk���	�MX 1��v��`���H>�G������yԅA��zgpu�b!��b��22Ys�.q,LH	��@��QG�0E�Pt^�ӵ�k�=DN�,��T���恑���T�z7�~�}F"EP!.�O2��TƕHW7k����1-�c���~W�A��N]�;w<A3�	$�)�
 H����#�1��������bR���~33�4C7)��}[��_.. ,�D�^@� n������'�<�u�������߮^�$7U�Ys���ϐ��3�[���=�i6=������l�F��)BPWZ���~)�����?l��%�4�|�V�I o�9ߢV���b�
��i��3J5�^���KZy����HV@����-n��3��q�p�±����7g�CW�ޔ5J�Dg?�o�7ۤ�_����.(�����Oګ��K�a@F�+b�tI��L�z�G'��i#4�xkύ�E�R�ã�N5y]VG��J�N��S�_ ���a���7a�*΋3C��,J�ښR,�s�y�]@0��o��_�G��Tp�:���3����׾�&���[�wr�T�: ���-��S��_c�1�ҷ�o�<h����+�9�Q�r�PP�B�9���S&�ﻚ�&cr�-��O@K遬��j9O�=[?�j��	���q���3�eTgk�Ii�kl7��hg�q)~�y4�����i7�HS$4&_�C}�����F�w�*Vș9�e��{Z��V�������^g�%��i�&�Ǣ\��s�E����������%'�gsJ�5�/��z������5&aIQ1���>�5UP_݈Wj���o������r�	��t~������Ҽ���c^��b.�GU)�$�͛Sa�r7(�K�n[���'s�o�_�w�F�L�`������h���V%�!���y��?�I"�\,���{T��Rz9�V��o�-��q��t=��&��jm��k���&�H�<۷Mt�lA�q`����y���p����\�z���3����\������l���w�Ŕ{�RtmBV�ƾ���k�ə���:P�2�A�~J:j}_��d�;��������>�'�A �h�bss�q	�~�2k���2���]��3W[�n��<��z/���0�d1a���|h�]ck�o���y��-�K��`������&�J0�
�5!T#�)��9y��N��ɭC�dHs𻥩'�GL�Jc�����ip��cB�\(��#q#�mi��J!�qԻ�hW������U�0C��o�N�����y�o��O4�},ú>�d�Ȃ���z�yQ��L�<9��oK]>j9o"�rm����EJ�O�ޝ11����oe�����`u�OaBY��us���văl^�1a,
�<h��k���y|yDA~���%�ON��n:�ݵ+��mܨ��|fȃ�K�s���f�֘N�MY��%]$!W�?,BÜ���z+�feMm=��)z���?W�%<X߭�����%���gCC��;�wT�ؾl.0��P��k+<�l�PY����P� ��Z�G�7I�<�[�:�`�t���5c�}�4c?U������2���sD���㕪�[�QC}ݨ�3�G^R{��ͫ���r�֗�X?2���[�#8��M�뉞ku�k�wܑT�Ft�]��vmJ>~�J
v��^�<Y�IԄև�̪�H���ɟ��ƫt<6�����5ײe����3A0PW�F�Ҝ��2�^Dq)Tt����eI�X�(#g@<�m���QR11m[�N>�7�BJ��n�"E��T<m��c���S�Qb9`����O��LM�I��I�A���0�Q�����i�/��k{��2j������6X�Et)�kW|a�Ý�������{�ڔ2B����#���N�8Bv�n (�i�_�����Q2ޟgq��HB����պ��'dD��U���'c䃙�a�=��򺅘sª�2ƌ�M��h��Q�s�Q���-��:#���sE�����q��O%.�Y֧~l��1�0�#=���WD�{�v�::�m�>:*�sIm�&%�!��-�%��YN�!�t�����H�mWTeqr4[�K�Rq���WL�=x�VV�6	t4����n
��[l��Fv8z�Q�?���5�M_�=���%�Wr��҆k����#�l�(�Y	.�ӷ��1`!���b�H/��e�m��/%��֧>���L��E?�W�,ζ��7�BS]�4L8�Xtٚ�,,�T6�q>`�w�n�HB�����ș�/]��[��w=�-�~N��ri�#o��q�]�e���E>��(�<���^��c|��k��w!ۿ��;T��s:i���5i�l�/���ɺ��u,�xu-����<M�2�z�ɏ�%��Y��7�P%�>�ӑ��B[U��9�����`V�3s�$s�o���w#�$䣐�,�׻6��Y'\!� ϊO�-���y>��w�U���G�D��[]�_RK
�)�ӥf�f�FP�,�?���6��x,�܈ <��&4�E�k7��jx�.k�@�&��#����ՙ<&M-��w�cK�>�3Y����`w�6C>}�a����ugv�.`����P��w}�)�˃O�Bv�tͬ��������_�ɺ'����A�:��o�y��NeE���T݀�S5X��ƻ����iƾfu~�@�����<u������2IKK��_���{mB{�6��x���~��k�
�� ��5�.<r;=��&��:Y��9��I�x����CnR+E�m�61���������%��\�v�������U1s� P���8U�[��q������~/�������Njdo�g��8<��SB�r���{��@[���� ����?���j�X�i��z�kt�_������
���teC�#[�7S���1��O�|�S&x1jm�c�yZ������Q��B�3 G�OA;�����X�$�hJ����T� �z�V&��9���Q8&��1�:P�p���Z�<v��t>�7��]ko�'�RjBi�u<�E����l���
٦B�Ts
���^=�=jM��v�����;zbd+�lJ]����s~�I��~.V�k��+�Ԛ�l7�\3����.c�<�9���0x���qŜ�����x:/�r+���%y�.���ￕ&�R�ؒrr��,,�QѨںڒZ|���U���c<�ؚ���З8�^�e�[��p�Ѷ���5fE�e�����卜N!3�t!vQ�`pW �֏����S�,��Ʌ%������h�KK�_h�R1�ejVo�<O���t߹\/yX�M���loE[�s����R:�n2�5����
�Ey*�.3=��y��Yjj��diT�[��"pQ��3���6�z��T^�RG�E&��d��N�V���j�è�Jo���bs� 1�7~��7�ـ�69N2��n}�ʠP�H$/�ī���ɽ�h9<P��n|���ooK�V���	Yuݹ�V�o��LE� e0n�7�18�k�*Gp�t��PA>?\y���m�9�Fl㑗�C)���q��"2t��Xb���i�=|ﶶə�P��#I�I*81������N�����}��F29�t�W �bb6�vr�>o��> /�j����!݇���]�].�HBw?{�.�^����0�?�9������Zym\�ڳ�0A��+�hȠk�����j���M<�[l�i� �G�<ې� ��_	���xT5��H�X������0؅)��}I%�yGKK��T���/�R��,)f��1�e�r|f���L�IC.~I�$k��O�����rG�����$D-���B�h(�Dml������R�=X�eqab=���[z���n���}��pX�+~��x��������j'/D�q��R��7f��M��)���G��f�g�s�ޅ���=۷}��G�	}_~��`��BZ����t��,?v�ɷ1`BR�.Nsg�˘r� )����~����3}��_տ�vj�E��Vw�и�^�z��FI��:�0zO�,�z"u���hn$�ĿQ ��cQ�+a[[������}�[J����H������р�c���{�ِy�3�����L����`٢���I��)�ZѶ-z��o����^����ң��·
��Dc�e�TD��j�Q-��H-�؏��j����Qo@u���'W��D�k��Pj�R԰�������a����(�C��Ad��w���j��xQH�U��RDj��*@�\J�tn�}2fD���WXI���+�>^K8��9Ҙ�5̫bb�@dK�%���A��I{��!�h��8��ډd|�dۉ�%����$H�nԵ6Y���m:k�:r������ى`��s~�Dy�W*2�Y��U?"C�B����+m!Q��nnn���b�w�e��Eߛ��[���ܽ���	D|9=$6���~�������+OG{3a6�9 �ؿ�s���<�:���1yvs۠�䁈a1�4�����a0Tb+�D��	·� ģ���}U�#����éA���r؄�O´Ԥ\]y^:�v��r�py_k3IK&��E���:V"߁f:�%���z�LD�Uj&M���6�>���f�k��nsU�Ƭ��Y�� y�@�#������%֣*��6�vB�����N�֚�+��������9��� �F�-P�� �@O�0��ӓ��Cqa��H�A�ȄM�]�E�RO��[>��k�R���f�Z5<��p��B4T��IH<`Pe��{G �vDX�jwEA~��{�ܑ�J_u�;���0X2�>��X��D(^A^(�ݩ��闫FF���Y�M��x��?�~��	łY�kD"���y钥Jl��\���)B
LG2��)��'0^��j�x�G8P��Ҧ}28v����1�{A����IFJ�T���@BBZ۹�^���4���� ���p"ŵ� -��T����!����~�>|47UI,�m	�C����|���$� G�m���>��;��XF��S*�������&�У��� ������]���!�?����EoVC<w�<Z��5���ns/��г�����*+��{TM���K�+�z&�����'h�l���:����&���_u�1;���2����Q�}2�@C5@瞴���k쨨���),�C��:�~qqaz2��;��� ԙ546Z�}%��m����mhj2�.Q�m��5���@��c�0R�+$�W�� 2ۏ��oн ���`�\��|9�BOW�t�m�ԭ�EG|�jʔ
�X�M+�� ����f���^�ڬ�e��W���L�+��XR��zH�h�=�'5c�{9�����A��[���E{
9�"8�a�/���.�̨�*�؏f���H��,,���=:)�:��KR�̩+��]7�SVs�5ɬ�����W���;�Oe�#M���W�-��k���BLPo9��{Y'Xq��8K�;�-��pZ[O��8�^�����-�|����	ψ���H�~�ֿ�ϙ_���!�r�{�6 eˁ�0`�I�к!������թl�h��������3�5���+�����s�������Q7Sm/U}y��t�Q��UPh��[b}�u�����w[e✝wTj�"��Gߢ--K�9^K�V{O{�C�>/C%���v&A��.�R�$ta�a.��Xr���
j�Z"����(�j�������k���i��֥*Z[[[/G��X��CD	�~u(��s},��*a͚��G$L�7��Ԃ[�l>;g(`��bw����֔����y,r`����1���\����y���<�ix��M����+��nŮ��d����Y��+����ى!�h>�Ǽ.���@�]��g|NN�K��"�UTa�6�AhE��
#�hDe #K��}G�t5d�}���R��[�Q݁����G�1c(a$l�9�ts1/�����l�[��||w^�'����p���p((�]��,x, �99�hk"}�U'@����t��&(�E���ϖ��88��uk2.Կ��:,baa��:���� R]����"�����Q���n:� �t"ZՉt�'C2ЇP��ֶ�8�G!��R��lmp[O��� ������o݃i�A��:{�6��cҤ������P���nӐ|۽��Rot; �*�@I��Ҥ��!ߓ�j4�o5vKQYd�M��,W��ӓD]E�7���}�-�����#b.��g�4�).�M��:�FB�D���±�Q������6��ѳ`q�QPJ'�~~J�{�=��3�b"�=nLs���<8.i)�DO�9� ݎ
er�]>��[�,�B��#��o�[.w��;�����$�ߟ�f��E5�a�G�-�m���)��~����}?�|IWz$j={�_VZ��Z9����N��5o>���@��]&��6q�%$�;��vt�uIc���d��0��cg�x�#�|����mh���z�bd�Uo�F&����,�LČ�P�`k5���SmG���ҟ՝Phjz:��d�/���0����t$�����KY{049��_aޒ�'�'�xOw4��Ki������`����r iU�&�+G1W����U����� �+�e�܋���cQ	��Hb���.wG8�?�­5D.[�b�B���s��Ė�Ի����W�W��@퀖zk��N٠�o_(��g�(��g�{�3��A�6,��8V�8DA�\
��G���]<�]����	�p�\A�f��~������^����;��@��Zw@,Byhd����nt]	�IrugN��tS`C�x��gY��2,cbz�u�����ܳ�yKI�:x8�vg��V���'79�B(6�XI^upu�Ĩ Гk���>X`Bp��C�2�Á���K��5�����D]2�RM��u�J��<�1�f�aw�� �S���kg�'`_�nu&��e)�/�U���GH�iao�!-�&��_��)���h�q#��BgCl�	��
��@r<zy���Ef{L����ME�Ҹq�K�,�䞣w��]F^E�(�U�b�𤋮���Í`��`�����|��������&Я��0c��2��3����}*n���K���[��x��WРұ_4O@#��ӊz��S^�5 P�j��CD3=�;Cz���*�xߪVM4P���np�Bq��O�u��)/�)OT�f|�@�R���-Jv=�v#d�pW�� � %?/�VA�u�.����&�$�`��#D3�P��t��㊄��B�1�����́�K����y����/AaYș8;�<��[C���{|�uύ���x����l��r./��H.2�$M^���}�Ŝj��ٶ}�IYv�E:k7ϳ?⒱�)�id�~�������/���lm��`
z������q�} ��8���u�Y�o,}"4AU��*��Yn��,6��^ɩY"�^D�3�Q7W߄.���9.J��Fs6~��:j����UV���V���[+��ot��m:�W��M��<�E띉�b/�I�S;#�J�� ��\�B�<'�A�ir��Na�����煉l�K���ިפ`Ѓ�U%BvE���`,�8n�W��#
߻�RO��)��H���y���ђ]Z�t����n-��w��)2��W?��A��'����^�Df�����vh���P��K��λf`wЉ0ܵ�
�=Rts��2a�r�g6�ϓ5AB���6��N�	b��B����r�n����/7NMvH�@&}�lL_���(�
�v�-��2���L���]5̿bDV�]�_Q��с^Ŗ%X�	91J,I����Ә��_Ϳ,�X��*�![P鉒�t<���gy���|��Y�s���(a2jh���9( ������M]4A��B��s GuǗe$�~��ٟ����#�.��c�$Q�O��"��:e��ۍ��;�M'���+�+�wگ�yZ���&�|��X8�_䉼~��ް�v��xTn�3�[9hq6�̇��r���� '��X��I�L���W�!�SDJ?ck�	mS��\�r�[�z���(���eu����AFLr���k���[X=�q�0ø�c��H^�v3=^��<hĘ"*A����Y��_4��%y�)���L�*�q�m��}�n�+\�F�����Յ�|Y�k�(��n"�Q�Au'E�)�$ "w[W%�8u�����Xf������LIG�WM�/�#'Q�ۊ��)D�� ��\|�7�T�߬����r���L��>�,y�m�Bs���Z�L>k~l���oL݆�6�@�9�~���Bd�gu�q�l�c:���3�j�m�c�ms�QLKo�����'��&鹫��O��"�u��W7�ޒ
�3!��U����`P����$(�ԉx�򡨵
�mvN��:��͸;��~�~��@��W`���t��W
��.���E� �
&��G�������:���vG��u�U��P!Q�ޤ1M)!(��@���Ӱi�>Z����D|�_�Uݵ1�2���і5�&����]�}�+>�.ح9���:��N+�Ԍ����x����p���ʐE�7������P|�8;�\�=���0����	���Y�������3P��VÞN�k�N��K���F�W!zЈ��:8`U>^����|��9913�e���~t��%���R��J�|�] �u�P��ر{�������� �����C�in}mG��������y���/R�2�_��>},+���Q_�#������N���j���h�[LbI;����݃2�u�4Jo�nsʜϭ���ytk��q��g����7p�xU�,k�%'����R�%(^nJKy�	4�1}Y|HZ)WM����n����@.]Q�"2��Դ����=:�LI
�����^!z�~R�̟"V|���U�.grwv��8,X����?����ִN���[���$ʒ�H�yR׽�`53�����5�p�ӓ|7�s��z�m�����i��p�`�g�U�|Q��0�8�@�c'�F�o5����pWӑ?'��]hO�Tg�����1Ϯ?���0��޴~7�h|q[s����m'�p9�l|������k6fV�3����h�A�T�&)���`�	��f�ۣ��$�IcL����:0ȷ[e�Ź����0A� l٘;W���n� F���]Ȋ+�����<��v��Xw�R�J��SB��	R�s@K�]��'�~�T�H���]�Ϣv�d-C�.��j����j��k���}�_��Ү`G� dac!:��XTB�?�ţ�Uh3��9N�5D��=&��/������-}<�5�Zc<��9�*)a�v�_gQ�쁩�ǁ�#���icJ����$�"o~�����~=��̡����!<`cv`�z��?��"�X_U61^:��w/5�:��y��֊���tл�z��朊#oo�ɖ��86�\��0���V��C�wF޵С�D������yk52���:�����*��1	bB�S"h����zI�P[iO�����E�D���/(a���w��Ƭ�g��tl�Ӎ����Y���ϑzH:W��6T\}	"�Y_PR�����)�g{����AtA���U[W׼?ՖHScW������xU�.�	�<o���
I�ֈ��**��t�~-��8ώ�
���� ��Wf�c��n�4=��"���*XF�u����[�$����~��\j��!j���TLd���(��R2���΂�~��ɉX	�t1[_'�^(�P�M�Dރn�)܁�{�Cz���`�$Cm-��TW\�8�z�16��!�Ђ��Qv앸��"�W��,nn˝�A	��OClՌ6���XȺ�=4�q��x�i��ZΈ���:-���(H|}�*K��l�a؄��1�((�-e�~�7���%�	�:����@�Tc���8h�7���E�lXz�
���r�Y�8f��+1��n�O�$2D��~� �|�/��p��K�CJ21_�1����rs��^q
��Pj;����j`�_��닉�E�G�i%
hd�uƐ�	��H��蹜����-���Ⱦ���Ͻ�jW/�}��oNܙ3�N�7�ĥ�$o�,o>\>E2���[�Aq�0$3��Ǒ��1WZt�I̋�3K��|�>6]>��=���Cw��&^���ZT��?�H��Y"����S����]�7Jns�+��C�-�6A�'��FF��%�f�ݏÐ��P����W;T%���B4�:���Eo�'�_�?�.还��~����r�1(���ɻ?='�����dm�;���U�lY[�����m�?	1��G6~��*z��o�[�}���pq376��1Ŗ�ª����"��!M
X�E~D���Z�e)�y//j��/ו�i�U��ݲ�jH�Ռn����P8��M��ʪ����'�כ1��*1���A��=�4ڦ2���j�F�}02�7_g���u�����ii>(�rO���0�)ҽ����9�&k�fub�ڠ�8H���ᜅ�,���Аt���5����A�JNx4�J����)��r���Y1]���va���Fp��A�<	))ࠪy�A�6JG����w� ����rl�MlUVxx|�)]_p�?�U���!}���W�]~R���@�7a>�T;_zQ�Y�2��.�?�_��������Ø��z�&q/p��M�Z�h���tTP&0`�q�n�9�.|���� �:P�$�N9n:>���`v��0�W��B��Q�[Z�y�
k��y!Wf}u���8�馉s�
� } 1��ݽ=)y�c���"����EL�Z|�,XP.7~�Gy�q�gu9s���u���7#����H�-^�O�������s8�o��$��!f5��qyh,��a���W0�+��M��R���I���K���T��ddrKKb6���CE"i-�]B�0�4�B�/4�{,�E�P(��O�X�Y���Gya�	�U�nK�c��ۇ���,���I��ek��Զ���+�E�'�$$�G�����|��8���7�W���9�,�hi�䷥qh�HnӪWgs�>6,�ik��[d�,�cHNC�rG��z4�DTa���OX�S_(
j+��"=<]UD3K6��{�ַ�?ؘ���Uڃ<$b�2|�-"�6;��,�KW}#��C$�Ϋ[�0F���q��P���-'�{�)�NA�yE&ވ�V�b
��)���6��R�6t�<Utii�����Z�t�!�O��{��ق�����&c"����Z.t_8������aV7�GS�(��,fTo@<�l�Qz���K�����:�f�S�ӛ��jE����հ��1�㎈
�|� {�m2��,Q��4�H�0���xi��+�f��1cϣ,�GU�uڼ��� -�F�;<�I���7���v��Q�/�Tک堫٦î��#�q� CA,1�~�B����%�a�>����؍ ����'yT�[A��"p=���ewW�r+�I�6TR�
)Z'+���b�����K��q�8�
K,8�t�V�A>�wz:J��	�82�r��q��m_#hҙOA�����;��k�d��F�[8���
��޶����>)x� 3�]��ǿ���>�>�S	v������LN�П9�aV�	����:�̃`�%FW����4AGG����aO6��r�	$aџ��}۷h��NR:˵Qk+T������ފ�u����c�T�Z��Qt�0ij�l�w2vv�e�WėY¹�)��H������i� �3s����Hc��f9>�#
���A��/�L2�C���q,L�);�c̉����@GC;�E�����j,�����M7eU������6��}�m>�z�r ٛ��[�E1�a&<�?��:*�����S:��S�.I��隡�SD�AA��ia�!��!���{���5���ଳ�����s,���·�ArA�7A�?ҏ��k��F�X��T����'d�Þ��n����]]</SLL��Ŭ�$��o�&����i���[Wv�"�Q�d=K�
 ���/݂�1�ۼ:|[ǥ��W�v2u����u9Y��u���w=�vࡪ�W?^EU���'Yk-��\]��sw�Z�x�|�@�����;{Z':R��~?$?�JKKN����P�@u�޼+���k7b���#�h���OMV��g���}�viݧQ���@1Gl�0���-��ڮ���L�&;	_��p�nl?Y��-�]��/Fŗ�������s��OKio�U�;��Z}8�k�gn�ך~���DZ�h���j��*EHb

�u4I�c�&��׳�lmK]��gA|�+��BGG�ւ=r�9�GE������3;4E�f�ŕ��ۿ����1�ϑ��$����������_
!��&���Fh�Pq�R)�l0���Z�u�⽞pu��x 	UaN�ñ�WN�$rZN�:V��y �p�!�ig!�0���G��*���Δ�јe�ϞKp�͇/I�d�c;��	bEU��R{�C�kB5�Zx�Z:��ӌ��v�������-��.�V�B����"�u��9>a�zZl��{:�-��F��Ġ==���.������]�YI�?�����Djk�>'�@/��ʂ	v��/�����X��U
���;��I�0Zt6�}��w-�dq0���m���/�ϛ}ha�4sE�Eg���V_.$�4٦��_��*1[�=�o�Q��>���c��P.W����yj�2�NVv���b���Y�W�/"E<���L��&4p�w���|�L�Th=��!��C<�@ ?��4I)�i�r@�Ԋm�}��{��� ��f1 �d�$D�~����H�?&���,�$����Í�d4ùJ� #��-��E�?JNK�Wd�s�G!��ݫY�[ſ�Ԛ�����fP�LS�D|�}M/r*�Z�uw���v��X�ť�njW�Ly�Z̨����¸���紲4�ӑ�"�vg��|��e���L���Svb�߆W���WP��oT+��0rj�*kj��!����[�����A0�i��N�Z����;�^[��Gi�N��&雗�~�T�ߧ$�>\cz~l�lזy5_��w���	w��9��.S�x�$4�~E�Qa
�r>��h�4��܅�K�*^b��d�?8��Tֶ����d>���8�&��3�>��2W��vvj�Xp�!>ٌ-�oO���'���a%���10��AW��$ؓ[ �,����%��J7[t���c�YAi��f
+(�*��xr���6&C'�)nw�}^�������k�$��_2$�=�%U�������1�;�1h��˪G�O!fy�-Tn?�c�&�&��c����6��r��)_�hSK�s����Aw�䃣_�xS���x�˵B��k6�3wyRHn�^��p����^�����u�'��5�K3����+��;k:S�;?nV�X�fB�����S��90�Ԓw�@17�t���^�fg�{D�n40'����WVjv�BFh(:#���$�A�:��ظpwC'2cu��̚沉����&q>�`�JAj¤��F
������ �9�	n�$v��g"m��=+ޏm�+s�������+��OE�W�j��0g�WQz,*��b�ϕN��
�ʰI�
w���G����gffĭ�h��^�9%#��)���J�=�f�N��6C��d���?�����E�;̐+�� ���4�8	��3�C8Ҳ;����F|���3[(ޟ\������g������c��^���.����\�=��[�rov���(�����Au)��6�d�Z��N)� 7MCl��� S0%�Ve,���:�Y��sa��3��L���{&��ߌ��{v 1q��ʼ�fܴ�]A��4>ԉB��r������	�	��Α��>�k�6��f�&���^��:���V�_��Yd���h�v��N�~�6�da+�j��.o�����E��+v���k��Si�8�r�К�P#�������r���+�Y�g_���[���Q;ntJ�g�)?�gǵ�Y�.v��c}�C|��ɕ /Z$�Ci��lz@A!c�����{՞ns�r%T1��״��pW36��<�g\IҼ3u���t̃�t�����L]ڰQ2�ݘe!v�\s`k)���(9l�Z6Y��(?ں����iZ�����Z�7�Gd�}�ж���JM{�y�'�D���"��=�\��f�`[k����{��W�Y�<U�D�~�������z6,����n3��� A�[؅<7�+�ܕ��=[�
��<�ʥ���y�*���i�Eȗ�zng���g�#l�pz�2�1:Q�$aX'Κp�k���=±�΢ҍj���U�P�� +?,w�!�ɋZ_�����N�����	�.���n�W����4�����2���>��\����=Wx��FQѹ��hv� �<�6+I�a'U���,��g�sav"���{F\��b?�*��{����[�GY�e��pw�����1���n��N�տj�-jƂ�:���-1�1E�G	�ÁQ���e����ʆ�w/�-��0�q���V���:wa��g�|����y����-̰r���t���`؅FXy�3�����sЧ��[�;��X��Hk\�c��>�<=ۭ-uA�1�I�J�x5�a!U���՛{^�Y�e�3I=�w*��.��i�?λ�Af/QY�7�%3~���yv5I�[W\G�$s����4�~�RWUH��0�
WCZ����G�������̆[Ƨ���	�[i�-n�GxD�n�*��<u�H�5�\�;�\	�{�z�O-6Em��j8��i��ꍍ��7Ű���͐�����E".�Ń�:TdCqdy�����9�2,����'_uǿ�TT�H.����_�+����}��Ӭ��_B�յ��4"Ʋ���"gB],1���x�'����)� ��u���)͹�Dϓ�5Ӭ\]�KO����%�YM[�3�	��)G��:J���p��L:��%�c���Q5"�9w<�R7A����xn٢����"��+Ո���5f���@�8B(b�2���p����6�o4���\���@̪��/���<����f���w&����a+}�h�ڔ�m_r�I��t�%��3hG�d�Z��u�p�˩�2��#��ۻK K�>�qK;�D��&�i#$�E����V߭�'��*��*�"-���h��t�A$�pC>eU����p��Ap*�{)����2W���*q���3ޟF7[?�O	�C]\j��t=��6����ͫ�����X^k*Ə���,��\'c���B��M|��ZJ���`as���'\�nwvb�F��/<e��A:��cU@�2��=/�g�x��~2��8�ֱ:a}J8��g�$��)�����m��,V
��2}�'���b��@=��om}Z��έF��F156�[-'�������}2h\��?١�O�00���g7���!�5����u��b��)�+�$C��c������ȓ�� �ZD�
�#�g����Fr/��u���(T�:����s�p�[����ëa,����E�q�7�$0j�p��H����
�Ȼ��OZ/�v�*W�^��5�[�B���	�6���"z��cR�1��XB������j��l�<�� k�/l|�t#��W�͎�,nV�y*�
4�Xlۢ�$��U�m��}MC����_\Ot��������>��g�`���b����_ʋ�\�ܸ�ǯ?��Hx�Ny?dڞ��Wu�|�Pc%��F��;f��.E��ty'�Ɔ����|D�M:�㔗�_�e����$�I��+���,���̾s�p���e�k�$:|LT�C�K�)��������o��.�| �flՄ�29o7��Il�����s�Ћ�d���zM��R���?k9�'ö͘�$����M�5i����[�����'�?�@}��m�w���K�lbkŹ�w�l.�'�A�W�?�S���>�?�2���0^<���%E:O�뭁'�Q\%�%��j���x"�R{�a��w)��l�.�3=ny_��H��	\�Sz�����7��Ч˳��\���,��Tm��f,���V��M2g�p2[�'�������
�N���Ob�/��C�/����k�3����>xŖ�3���(����e�����6�3{4J�/��h�iDy_��ʈ���W5��9�X���D��7��2_��h��@;�hh�9�*	`E��@�X�|�H֣��+M���1n0��͹�H�|�E(1���v�����n~��D�m��Ʊ�4�;�y�>Kt1N�n����=+��Ý�e%Ohбw�vk�Ѐ7�b�b�(�򂶵RYScH�Ϯ��	Q�p��#�zV|ZVܼ�;Z�`�+*�F�ɩ|�%Xd��;L�����ӵ(�! �vM}X���\��X��yJ�����u8���6-_��x��s���4�D����[��1'����hc��%�ធ���&�3d�sx�1�W̧�) Q~F�V���m�7����ϕ�_�d���_���z3N����v����q�s�-�V���d���g�+jڋ"ĕ���=h%� ��B�A����G��������HG��v�5yq�-7���B��r���9�I����)j�l&����	ξ�P/���C΁�sXP��ŖI��E��9��2�%'��`v7H_V�{ǅ�w�L�*�Ɣ�>�t�<K��g�uq��*nr8"}�~�{+\es12��T�I�8�����8���qI�Ut��#+�5�y�wv��k��0�O.�n���V��l�//.e�r�������r�$�Ɨ{�!��h��.{�G���r��?�]ޣ��9[�Ns�[�_����);�:,��j�4��T��~twy��ΐ?�a�r�t|t*��{<ud ���t���]�n����E Ua�_1	�C)ف�b��]�Y���n��XMw{��å��\��J�~����$S��eEf���9�S�ɗ�M���/�>�I^)#gI���=)p�]DRyV���sW�ĩ�q�IasZ���u.�Z��a��X���Ј���c|�b�O��K7*性��e�Ҿ,k�0䚥�|A�Ҙˍ�}�KU�t��m���C�KЭ)I�'�5W�}�s���9 ���=���[!`�7fA	����*�`l2��T-~<F�_Fh0���%#)�Ά�Å16v��w�������D�Ify�C~�1�JxR��I$T��	���<3zv�G��������ox,��{pPna����5p�υ���ur���AXK^ل4V8@��79�B�X�&^���_PV�ۥ�9;��&�Kc�'������S��Y��\����jc�*I0+3V��g�j��K�g��]8!B�E�	p�7�m��<Ί~zlɾ�5-�d	����O�YvM�>�f����靆�Ew��[ޭvܲ�-WbouZޕ�q���%� nWҬѽWW�������,I��w�Kw 9��=��[��2'�xbdϑ�������* ��� ����������U�c��IeKO�|BN <�4���q����L\��T����2�~����^8�q�.RV[�<���]`!E=� �N�_�$�[���,������	<���ht/`'���e������R[�1�-��o�"*�N�k��+���ٓp�D��M��ɕ�#�g����vY�VW�D�����Y���M�B�$��W����>w�a�(���T/@`���B�84gزeTΑ�K-��.ǃ=
��c�pT���vt\1���5�g]�������G\�� �}7(7���̅	�n���"�9��/��ik�/&!`Ӻ,���,v�����8ƍ�q�>C�'��Z��P�����J	�zG�?ˁ"�Ν�#��9-�-��R+�a.G�}3��2u8��9�b�_	[�p�8�H��-�[�C^���nX3+��9Q�O�o1G=w�J��[�F i����~���PB����8��F5�V~�:�b�t��Y���e��*+������Љ�Y���=^����`V�O	��+��X���
+�]$l�d�������� �� ���Ȝw;�pI�u�7U7�Hw��{�?�Q�ʬ[���/ex�����q�� W�vؽ��&<z�o���ۚv�[=�K]�]�@���Eӽ�_^�<��>T<w\b�@6HÍ/�I�V�F���KGW��6~�����hi�*	\��u���uM���Ž�;��4_�Km�XMz|�)[�[nN{���O���i+�/z^"a��~d��L���#ٺ�iC�}o�<�-�W�N��;8�}U�ÅS�����7�3(1�z#� -�����p$W��.�����H�AK��Mn�`��bO�4�1��ٿ�5������d������p�4s���Ɖ5��c��X{�Fi�cc{�:�B�{�fc���[ �p�,ꅘ�G��L�W��	~k7��|ςڿ�5~��~i��D��������Q��2q���mA�Y�Wl���ӳ]}���(�)���z���_W�p�IbJ���U���U�}q�U0/�n �K��O�/�e������zl6�n`	N �iE�03�@r.�Pd�+�b��í������e�5}�ajby��z��!�t|u�	0�+\�ѧ�~u��eV��i�3��ox��(=��V�o��Vצv�f�㯱Ʊ1���6qS���k�h�� �+\nmq�r3���/�d`������[���ڱ���B$���~��k�Bx��
Z��źZu�W3�r���σ�m?��Pj�=[;۝nv]{>[e����f;I��V��4b2g�U�`M���&�ľ[Dk�����d$�M-������A �\�����ѷe��证j$���^��gU�&� !�&���Dk�@��}D��ٞ�UبF��!�Ƨ����m��	�sL[��H��I��W��Y�����*EA�X*5�a��{��u�;aϋ3�|ˮ�&|��r��HD
�k�fp1M����4�,W泛��&)�Z��;nEn�,�­����	̺�I�6&S��	�gA�D+5������rL�mv��5�|Y�_{\��A�s���^�gG��h��}P�]�W8���Ջ�5�*��-��'���.��Z���s �S����Stt7�;A$#��&�u�G���[��}HT���(�!L�e/Z����H�_��{���%ԇ5N���W�IyI��)Z���O��J�b��>��������R�K������\Hn���z���G�}E�ihf	��	ש��="�p�Bu��B��]�pX]�y8v�/�A�@����X'�M^:Z�r��*f�T5�@f4��!�y����d(�LĢ`��a�k��b�+��%�+Q\DfT�e>.{?͂�
0ک��J���x����8�ؚ��3*cć[c��?�A*)�����a�������6���y�A����zE<i��U70!��I���!4�Hw��4��ݣ�;���;AGN�ֶ��M�ogg���X%955����g�(�x���0��q��冱8X�z��f��{r�>_��Ķ�1��y�m�`a�9��lH�8D[ϓ/mh{>�$�����ً���Lq^��ǒ�t��:��.�3�d�Ę?�K�YU����ԄҮ��'K�'�����-�5�D�}
�t�pC�'M�0@�"ڟ�U@\$~EĬυ��&W�b�����Zwor�_����a.{,�z���zmXJ��,��x�˂��cr{,�()��I����}��'���[
r�OCK?Re�~���w�N��-s�X�&�8z�h�~Gơt}x?�v�wYg=�z�u�"2���%;}D��l���~2[Re�`߷�RjWjk�8�FiP�+N��5i8P���]]t<%��z�&�3�P�]�4����׋=H�֘�hW�E�c�p�/��ċ��˼��%�+;��Rlۢ��CD6�T4�2XE��o����t'��bg�h�Xl����<��J:���o�S�CI�όJ�+=V�.���Bw�b�I,O�gr���,끫ID`۟��@)�걟͹��1�[��k�u�ہq��|u��|���A�A��W�L��T<��ٟY$�B�7�ᔔwDVzuYxqx�A���dalln ���d	�'����^�-j���޺ݤL��{Pb@n\��6�Q��+e*TI�Ӓ�H/�_)����Z��p�O�����?����܈�V���b7ĵtcW�Y��6�9�Oh�2=h�u�F�a,���I�K�cZ�c5����s�I����XD�5�bHٟK���	Q�b��PA�%lXY�tg��c�S~}� ES ���#Wd	S�if�ķ����gY��I��\�
}2S�R,������P"���F�(3����m=���"���ʋ����Vg�~�{�����j��ô��?����h�"%�������Ę#TqK3�K�C��B���q�so����p����v��,��Ĭ����?+hBK����>�Y(=V��MB0��g[��r�Z�P���8�L{��|�+�'��;�98���ߣ]�3 :,��7����2��*�ڍT�	F$.J��mJ5���gJ��zpaU�zs՜��\� w��M�֥���Y���kL%]Ms�?{/t�7�Z4�K%)/��,!��|B��~�y��p�)�F+%�6z�r$��y�X�ȫ�osd��"�l���7f�V+N<&����q�q>!������*��8���1-`Kx��y�&�{�)|�g�J��-Ye�[Q�L��;K��.=�����G��$�3������
�hV��n��-������+ss��-m�o�a4����v&F<ݘ��vۍ�ia{�U)��g�	,�>D��f�
e��gPdVSp6��_���K�� �����Jf���7��� ��6N:�Pe{j�
�/�B�>��p���~�KZw4''��R%����\)�W4'~���Z�.�}���E@�_����a�=��A�k�>c[�4-n��S�؋X���{�x���a��4��"�7g8
�L��ؐ M��B[��VB��#�^��b�5�s7\�U�c��B5gDh�\2l�V��<�U�p��7��� _����*����-�m�Fs31R��5?�:`_��.Г6!#�@������u��P��xNω��$�ʸ(�E
��г���eɓ!C�"q��z�V��q���A�F�����	����?��ݒZrx3fV�s� ����5R y�@�������x,�&����Q����	5���#�~�9Ot��2��_��ܘ&��_�YG���"}�'�k������_� ���19oOv��YX4/�98
�B��g���b5fϾ���:~��9r �qB����'1�]H��b�����XLL.�9.Ķ��g:z�����L��R�}������7��4~�h�Qi���[:+�#;l
�|��q�������2}���W�c*�~Fd��5X����N�#�B,��W���~��/�����P�.��<׊�a��;XeM��6��� ���XlW0 Ӫ6��U :5����gV#h4G�!R���lc$`aʾ ���ί�u?���K%Y'$���>S �	נ䳺`ᣞڎ�`-�w;�A��v ����F@H��f?='��׆�^�sꏕF ��p�e��N��]����lWИ6Yʤ��
�@<*��ῐ���޵O:�~WR!i�1Uv��WG������ŉ�z$�n����Bj����o����!����ڔ?\�ߴ�] c�2��O�P_䌏{����ϟ]��0���W�7�����I���څ*����!�!c]���7zhl�j���	��R�A*��~m���^*�a�+��>�ja(���X��NX>�N�xb��aA�`t�.bsz�:�"����^{��;vZM_1�Ç�$�vL�� )!�yc5}��W:��c�JM�k�����VV���27�t��,[I l�sr���q3�Ek�f\���Y�?�@"�2�T$�Hbig��=���.�L9�}@-LLe�DZ��^�#��O������Ո�w��v��2� �~�:B�-3�^���!�ԕ-���`3��C�N��"tAg�A�EVY�B��ҝy2~���\�K��㱗,�0{�}���iʻ���;���2b1���G�ҿ�ʹ�8�?H�r�GM��g���	�lP�  ��/�/z��2e�^��3�$gj�K�8-�N��2.����ђ�! �(��y��&ǞN�{��7�ק>���ݍњ��[�æ]|�_�tA�����A#]Ɛ[*w=,:^~H�G�A�gr����a*�űG�mZ�g~\��^��\�H,��4~e�w���rqȺ�Ե�ޱ��R�F�`��ɦ��-`�㭅����3�t��|��}B-t���G�I7p��
Vm9V��iaI��?� ͋���g��_5�����cn�1u?�����ňk��E���q���;@�e<S�_��O�Hh�U�ڔy:m�@/V�ߖ]�O����RD탣n$�J�Ԉ�u�J�YW	���=��6��Q��̈���e���\��=P��[c19���*��z҂� �:�m�ҧ�v, ���*�2�q]@:�va�F�K
��E|V��~-��F��i�ࡪ�x0R��ߊD�Ws�`�F�'T��|���������9�r��_�T�~����q,Q,r9G�����w��I>�G6���K�wGD2X].��ĳY����Xۜ���f�z��K��������!(?|S��x����oTR�"��~�,�߆�Y�{_�l��07��CQ֜�ќ3v[n8⫆d)W��1�m~n��;�������X�]@��8���m�{���x
!�|Z7zHsQe����o�14勃T�����F+Xح�v��>����Ԥ�"���c�i\�-�����y���ZIM�
�������_�UEG��	���Dڥc����3W��F Q�)nS�G�/���e"��m�tj�c`ﾮ-�~��%1�m
��o���r25�'y��9�~�S��\�$�KE� Rlc|��{S�Ŏ1�lًjĤ��X�ъ���N���1�]J8C����G)�=����ym���Q�0+��lϧ�+����9�Ɂ"Z=Y��8QpLR%����p����6�|��s��Y�������kr��L�Lrr+G߰��߽CB�2�W�/����_?����o����^�I0L)Zcuw�X|�?U����x�0j!-ꤐ��BOc����\~8��h)����~�_��&h;�b2�F^">�^&�,3XW�����,�+ݳ���ʺJ)�'����e�{z����C����P���t/K���Q��������~�:��
U寪��^E��c��4�l�P�;Xgs�����ְ�\�&?/�t��I`�t;>f���s4�cz3Br%wЬ������QV2c�$T�$�����NםCKM��x��ȫ�Mޫn����Rm���n�<�:X�@���/�L���r���Dkd\�hT�FB�p����"s�6 Z����}3Y��R��j�<Qـ�������ρxڨy�W�C�>+�E(l�\-��"�D"��k�Ir/�+E��}�	"3��M_�7P�ݔ1�	��	&Cz�߾$P��^�62z���xȵ��/D ͧo�d}�d�4�uyV>z&v�%3��:!��t�l͔ä���Td�sR)G�l[W���bF]:��O���Ў�L� 0Q��2�6ti���D �q�ُ.�������(�����Ŷ�XZ�L��aX�z�|AV㩲�4w�q�@��ƭ�l��¥}'��~��i���D'���A֟�i>��l��<��U��[��cK� �,�1؉;O��r���+�����0!�lOƇ���F�R���d�k�T?���jIEK���OC�a8�H�
6S���]�b(x[-Hx���Zl9�������D��t����-����ZjQ5͏�U�zjuOUr\i��1�H����U��/	��	u��ʿ��݅#��f{�J��dY����J ~qËuFT�.f4#K����C<t|,�� ������7� �h|��7|�q5>��%~��IX��j��e3��6#��0��+�2�`)��i���l��i���GL�Z��cV7�~.�!k\�B�X�4�����S�4����
D]�"Zfm������zڲ�4s?��L��9R*��=\+�{o�͍��NԈp���Á����4�rk:@�/�m�1+�8@Z�J���%:]��m��u%ݹ:�f�J���P,�g��w�����?��/8��
$��/�ВC*s�vI}ޯr��m)���J��w�a�e}.��=�?���(ܗL�4�� VZ���y�+oLH �76� y�jqzv6�?�e�y���"��ӂ4��ܭ��uɛeR�����ʅ�c�}T#{پ���'� Ӟ���H�)�T�}��B8��)�e�B�5�v��/�U48ca�6�ue����l��_N����F�n9d�t�K \�-8�:��lܤ��!c�G���p#�Un9���&�A
����j=�������� ���9�F�$����g�б)�}�]���(��7�m�^�p3ت����:�Q����3��Ǭ�r	8̒�J��dpfSV�ҲJv����/f�3^Y�rq2� 9�)��εÁj��ͨF�X�D�xg�x�^Ѣ!*5P���&��f�8A��JSȟc���h��y�*v~E+y�o�Nz�����z����QVg*�7��]�Ku��
��	giii�k��iv��7_"d�9Kq�+��Q<Ԟ�}]
Y'm`�S�X�llLj?&��lq!�%ߡv�F�ū��7�6����66��p�z�Wd�⺸�_�c�2F�61���C�����\��ѯ1pCg���q��]Lx�b�׊��y�RDR/qa��NI��]H# PV^k�7���Bb��,���t�����2Q�|}��Q�����5&���$j��R��4�x�h���.�^�"ۙ����DJ�?K��&>������7�,ٓ�h\Q9��"��b�&�i���|���)��<*esL?b��t�����M��t7�س�D]R"%^$�����u$[泐1w9���YcJJJZ��X�.��n���C�S*
J���᫩��I�u�U�����Wڢ;�����DX/�Fk�rat��n�g�z/��{�~�t�*>��NFf�"�.�����B�\�jZ�1l�#냳oT�_t��ĥ��j?� �vM^_���`�u�	E�H��n���u�i�=���X�0��E��9k�}���i�h�*?�3�#������s�L��x�N��U�<�>C(��U�eV�e3X�[a��O�b�Ⱥ��l��}h�q���l�����D��W�S
T���GվsS��]��+Qn��/�<�p�5�Y=�g
E��sM� ���vm�h0�)Zs�t\N��5�@��K_���kV��_�w{����X�}ץc���7V��cV�b7��2?���,����Wc(��*6�j��^5���C���6`�[����=`� |�	��z�D�}c�6�����ٖTLt�����]��<��Cm�Ƚ��ݟ�,��RL��b�doTc�C�i� J����b�(G(_-�p)���͑t#A�ߓ�W���s�Ϲ5�6�޺�E�����dm|{��E�U�.+��&4�3�\ �f�	����Ⱥ"O�P�%�:D��,u_����E��e�|��2Y�
]G)�7#�H�+�>k�= B�-�����gU��շ�BFm��kױ!`af�wsy�����9�poL(��K2��lݪ�c��M� I���؛Sꥇ���$��
�}��q��움]�b5�,Vd��O��)||%###^$w��;*v��cT=�(�4>P��hP�P�m[��h��Jv�>g����[��tq�Zi&���c�W-�iR���
�$ҽÖ��]�b�
�
�,������5(>OMAD��-�ck��qt�Z<��f��������.��O��By��8�A"�6�:)�?��w�>���wz��z�O������~"�d�J�u.��������'թ�n��谏`�qJw3���_�A��I�>�~�mBCH�ɽYEP�,Tr���]ѐI��>��7�ma��%�����<�d�z�_!lT��Sseh��͒��,l�h66>q�$V�f[�� o�nGm/qQ������]�tw�����
?�V�<��� ɕ����@/c^�q������P��t���z�k6W��9�?�oovC�CGϐ�Y�7�(�z�hL�W�h��&qy���=����=����>�6�,��_?Md���#Z!�S!����5�Nf˟�G��q�Ad�x�
>|�>���@/��o��/v��6��I��^��m�-��ԈVm�	q;Sn�o�e���K���d���4�X�~��#���)���]��#� �ˎ�8�Rko�9�W	�b���i�\cΓ����KY��~�N�D���c3��H���41k��y��P��NZ�r���!��m&×N�2��J����Dm����B�m)1�o/����3�^[��Ϩ�?$��?w��m̕@j��΂s�f��{k�U��n�M��y٪��X^�F,��'̸�0E�AW�~[�˱�LdM}�����5b�O6z �AJ7�V<nVS��5���K���������n���w��M~�|�o�˳&u������ժFX�@v*� �|δ2��Pwl@��X��y}�j�(�_F����+�$�
)���P��E���� �)د	^f��(d�zp���a"sJZ�;H@������%q� ^��~T�̴k��)�t+�uI��5A����smΨx=�Rl�(D�� :�1jU䡴��0I�
ko���Zu�<"�L%?xV9�z���7��B;�܋�P'I��جZ�����UZC�uEͨr�����Χ6���mkc���^A���c���6�sRo�=��mE^�HT�4\���͠@�G�?�ޢ���oV3p�����L�&dKK��aI��P��R���Y\d�Y+�W��D��LF��hy�`� {W����wq��1�%@sp`��黛�2��[��UwSpu2�s��.��/�9�,)yy��S�m���W���/��.�SZ)%��~P,�[G����d�5���!�ߍ����?�V+�_^�i'��y��Y�6��?�ߥJ �+�� �3�Yorp�!Ⴢb`��4纾�e�*/%K�kҏվ���ZӽY���O"�"o�F�9��B
�;��_Wԛ-�)�?���$RZ�.�n�4򷌌�,'w��B�E�/���/�B8��bͨO��H����$���(#>oln��Xw7�2�A�{�){�����5�2���gCnN��K������ ��� �3��h�u�*�Bdy̟�1�&����8[2"���`�稦����|b�f�²�ⶤj��i��j�ÙN��_:<f)��|PPЁ��L?i�׻�w�Dg(��fި�Y�?xT&��*x����fi��2�^?�
u�����0�_A�F]�q8��#E(lg)�����v��Ry��M�g���Ǔ��c���H���UPQ�B�u��0��ݎ ������dV)��;eQ^�S)|�g���[&Fk��u��us�ß��8O��b��D�]޽sx���o�Ҙ���j���2��/�-�ٿ����s$<�H����i�!����Ki�\ 
��}i�Ł%�@���Ë$�ۯ�����O7��L��*zw�O����ס��'q4D���$1ā����S�uj��s9F���Q?�g����+��}=Z�[MA*��WN$��0�Bm8�ex��P���W��ۖ^.0����<���X��g�Մ{SƆ�n�Z)�=a�c���Y������R���lh۠�:���[�ڃ�C*�i�!a�Fłr]�A%���R��oVX��x��/�>Y#/��~0�4�H_C���7�:����ٝ�$d!��..ˑ؛䁥��=<{��]��׫a��-�����>�o6s�5ro㬟�G��T�R���*K��G
J�h�;1Đ������"l���9�V������F�B�� Z-vG^������yI���7�GZ�Mx�7;���q
��I�+�`�P,L��J�4f(�?���b&���;.3���Ѯ��W��@φ����pg'�!}��m��ߍf`ApЕR\[X���mӝ���̈́_�n��@*���j�T��DK�!wk[�3:`���Jʮe�N${�p{dmg�q!�q��m�șo�!0J(�vx)3���4������[��l
.顨6���.1!�7I�V��R��8�9�_��M_jjͷ��?��3����{oѓH-z���#A���E�DD���^G�ޢ������{}g�������>g���>{��hM}�nY�0酜�� ��Q��������eK����6��G���	���K
���Q��#���Ir�'�7��?+��`C��c*�}���ԟxz� v4g�KE�&���k��q���UW��q�{���_�ld���w�%2�p�S�>��{X�xA:Mڛ���2V\�]�ꖕ�{0	<1y��o�yz������	Q���6F��r}����u�8Ib���b��م�����9�Y��0_>�鿪��*h}��lh��
v՝���{�a�حƃ�J��8lsL� �A�W�H�8�LM(�F���$�����J�`MQhN*�����ɉkso��RS_/��9ѹ+w���5�����K񼽪�C���_��_��[�P�e'�e�餳�f�����LD{�\o������Ǉ����V3��Z�H�o�>��ײQ!ڶA)<` �ŏ��ɶ��e.�����ן���D���IvK֋��p�ɑ�x)A�/�Zin���m�'ci2����S<��ñ���z��MS>�#q���#ҝEz�p��[���y�r�`�"/dL�8�N���,����n/�t�ղc�/K��zP�����o%��:��x�j�%؍� �V�̠a"��;��K]T7�Aᦱ�;b������P������dY'-L�w�@[:&�����&%��+�V�fZ�'�?�J�z��ٳrM��[���){�Lju|/����K�3\���Nd����R��|�1
��a"�z׀�J ��Ճs"K`m�2���G}���_�䴡ɔX7�*����������������h\����qR �)�/�p�|;r�o��tص�e�ӱɃ����֛�}S���JFi����w�����<?M���-�X�H&]�b棉�.��͐�>���Z.�)�VU�z�N����$�MA��bykC�!���@xN!��E���f�9���4�҂z�rJK����1������;H�e|��&�/�E�ȏ��:��ೳO�<i��ߨ����ӣ<::z]C�C�TPP�<ۥ/.)Y�9;;yw{u�,�E�,���J���#x9R�UY�R�&A�����&<{Ϧ��~G�4�:��J(��ۡi]����0�_Z������|�_��;W�6-���x,�8�8�T����w١׫m915�o2��5o(��F!'%�˼4�A��9�h�q�3^��)횭pt�턲�ؘ�D�����ls��QNlu���!��$D ��k������ ���6ʒ...����[��=N--�Q*3y�� ^���Da!���(ZR�y~͉z�?\@(~���^�fg'��{/TBb�	+�B�*Vf�p?4�ef`�w� ����n�g�ms��g=J�sx|�GDJ����ʿ�ޚ��-���8���%3[�ɯ종�����{$%$F����y���x����y�I��B5�_y/�F����`pBb������~O��^�/t��+�u�10D��奲��i�����^	�9�3$����hu8XW��S��j��X_s6E󇗻w�F�G���kdX���"'N&7�(�׸�n#�$>s�� ,;���|;@c
'٢����`s8s-��gr�3���^N�Bܾ���~L����k�:Ȼ�k�:C�*�Tɩ�6M�}�<ݍ�	�9����11�h���6�|��SMъ3.RM,�$,8rd�F]��6:@`q�b�����n)�*�8�6<�+Y�7u�7u��я�U���g}䎈�.Dsd�O7e��/ ��3����4��mz�m����߸�^������{ ��Zh�|K�u(ޗ˔�J�� E�$)�(��ǵ�Pg���ǿ4�����n��NHBW�=,��k�����Q��T~g����r5Vr#uKR��3?"N�ʶ+j�氧ɨ1*!>���x*>U��jgdW�}�����J�r}�,ٚaV#"j�{Je>{~<;1�jA��H�b.�<Uf�Fn`b�(���\);��2���6��K^K+�y�De4ۏ;V�|���8���9F�4���ϣ�	ƧD�>�*}��S+]3����~mu���ĕP��\�����󾤤���­NmzBB*���F�b�݁�ZZZ��E�s���?�v�B�b����7����yF�B��T����D�M^�	t)
�t�E�.
˰��+"nϾb�2����`�7��K�;S�!X�}����0\���u�{aZg�{tɸi���]�x�}c�wXi�����@c��ø�'C��*󋺃/ͺ�����5x{�	`�H�<id���7�pm���KeTB6
�#֡�6��;l�b���[��H�Jy����&��.���š��''W���> ��k���#~�q.�=̬�U�Q���[m�9��=��'~Y���[��k��D��*�^д�qՊ����e��
Z�3xun�2]i��������S�X��|�w�_��o	��a\�DX�X�%$�n��M�*M��.�ɷ��V���ř�ô.L"�F�	i����x�Z�1���V�m��떇�~r�
O�-I��!&��w�^��={g��=�������#��f���QVW~iB[�;����V-�kg�:靿UL%���AV<�P�_����rs[�a��G)�~����V ��mp�Lq
��ފ��v����N�w��K�t����U.���u~�wH����dSq����,5[=W�hM	�[�������mO � �Q_R�_�@�gs�w]��ԃf#�sw����J������f/15<�?�.&�uc}y�.�� ��NqI~��0�P�c����ٞ��2�S�G� h�AD̊�N�;`������mvC�$������g�˔����|L���D8w������;��b�diGH�N����*�\��K,ܴo:H�ј�^;3���6h��K�g
�C?��u�֨`cUz�jH/��W�oV��+q�A��*�s�tp�TQL#j2�D���̺VfD�B��k�<������W
 ~W�����.1I�T|���F<z�yMb���	�y~ն�C'��뫊�����s/���S����IB�]0�;[8q<��q�FGE��-� �ڽ��
�HL3酩aS]�Y�WߟvA~�6[QZ0�-EO�ƍ��s�c�T�"����s�uT�����)<��'BXm��6����f83.�	�Em`�j�h6�3�c�˭�����_F��/�z���vgy#�	˳ù�_�{�B��/����Y.ꤟe=�	28�=��貓��`�T� ��~��&JT˨`3H�}u�;��η��Q�E��@�zv>�4

S�NK~��Ws`�b���1��ҹ;(���#г�8�$�|�e�0y����&�*�|�'��G4�q��:�Vi=����I.7���/�qŶ	ևZib&����OV<A<w��)t��Y��[_���FD���yH8x}�4BDR�S";P�"n��;���G��X�!��(�:�3͕�(��o���&O'4`O� �;�^s8����uv$l�:�Ď��D�gy�v�����"رԅ�Y�W�i�`���1�����B��|�͟��|��FU�kjz'�^c]T����w�\���?�:�||����k\e
��}�(����T��뇽c�7V�վxϣUU�m�L�x���`Lpv���U_q 7�6b��W�����_<��	)��[�u�����п�-�������{1O��A^�����O�Ž=u��#��?��Q�Q��R�x&ɄZ:��+�Lsh��L�\Z�'��7���Ik|�U���)ڣ�ذ���f��$�^��i21g��Z'�#��������׀���>W�s�7km�A��ѡ�8R�O�D�o7�bv>bk&=A�|I��"�<�m �u&0�랡�o��nu����:�f�KZ��xEX���{��
Q��a�m����C�-�t;�e=EV��B��/Q�ᔐ��8^��g��Sşp^�މ��t�����R�bO�t�ssv��!	{�Z'Y����06jc�q;��.��Aeo����w�d��k���.�:�[�Cm�3�Q	}����-m2ch�n��߶��%�\��?F&~��L>|\�����f��[����3�+"�����(Z��_��Ŏ�	�=M1b�\�/^�(�u����R�2�YvnK�|+�g�T��n�B$��x��H&g����h% h`��D��ﶷNN,�"���`?-��N�b���y-�t�.,��s��}��H`�%����&��ٮ�3��?e�_��͒B< �}7�����; �g&qN	�b�G0��=m	��Y�������q֨�~ei�7bIE9k���'k�F�������P➳���Ew��HD��j&Kxx� ��2ݚ�8�/{��5#A�߰�y+]���y���I��3�}��/�l��F�� �$D�O~���W���J��%�&�?H��Ox���I7��,��+NɿJ� �#Kd�����D�����*j����d��rE��A��	�Z/�}��H0Z#P��3,>��7��DK����_r��,���9�d�L�p��X]_�J�i�ãP<�q\��s�~��S�m)\��Yij:�}rIPyDр�f�����S����{�2�S�$�NZ�Qڡg@@�"/�Ct]�d��t�V5�Gڜ)�i��Հ� Zw��n�z�����q*=3.P-��\���`��W=���,o}�`�6���������"*�_s'�t�2"�y:4�b6r�ik��Ͱ��S!�Ѐ��	�ah屵���Q�cQ���4���]G���!��	�\�%�Q���p�O�J��?/�'�-S�vuay9�*��6<҇�n���!	�d�������9w�&�wJO|Y�$�bw�a�(�y��H-�����|bp7s����@����*X���R{������Y~y6>zĚ Vǳ����F������Y�ɿ� =�(���Qg\�m��Q!+�xDb5v���x��^ ��J��&���j �jqK�fSƿ��yC3(�؁8�Jz6�̕et�_s;���"�7!�uT��C�!6�~�{1��j�H1�����[��;`탬7t?~�>�z8�aq�{u�7� �o�����Õ�f!T�Q��_�R$�<�*�u�z�W����/�N���)��z������Y��&���M��X��3�P�">��0e]�+���00�����M������6/ND�����B%��h��I�d��`��µw�C����s9��X5�B�Z����~7���?����6.`����_��"�1���n�6~�����\�Ĩ�&$�?�U�M����Nj��CAf)�%��r�z{��0��%��ׄt�2���I3.,,EJe56�P��At-��F��4�&gg<����Ʒ���²�EΧ�I��<� �(h�	��$k�sB�)�=$~#���0���7�9�/�q,+�c9��ʹ�U�.��/��E�S��0�P4wa���n��mFU�m�b�>9n�ց���ި�@a�����(�P�X�l9��JQ�B�2WJ&�������L�H�>�ϐ��]F-�9�{�ɾVR�?:>�w���s� ���r!�|:�aS����d��s�rR���S��I�Q_�L�yc�)M��i��n�6f#iqȘ��ܙ�bO_���2�����ȟy�8��V������s��fۤ^�|��Q_����*3�
۳��8���6#�Gl�Q��t�����ŧʋ�:�:�@\(��RS_�s�%+S0�+Z�B-�Z-�d�b���\#eggg%�o�[O�ߖ��&�LG��$A�G����P䯞mb���23GJ�*K�ﶟ2�l7���	qq7r�Q�[��mMz�~ �?�J���W[�"�X1rL��6%㰔V�n�����c3�=!V�����t�(��.�T�P����uض,�D��6�a,H2� �������vG7t�ƒ�M���ݙ���ȨH�5�v	ʝ0���zT7D�a�K��L�SpGQ>�D�eJ������ ��(�p��1e�9�>��b�N�N�z�N������I!�3c�/zb�<������V��VPٞ2�������b�����5�k����@d_<���N��^GlƿvHRB���#E�Nr��:E	�$�ϟsw�iDO�kp�A�L��±�'W敮����֘�=��;���jHNN-�d���D.�j<e`B�8��ۡ<g����>�/���V�a�q�
��}����FF��O���A�^T��{��Xg�'��#Z�}+��|E�m7�ݧVkE(�YG�2S���'7�SC�.S��j%��^�u�[��<��;MJ��A��rr["�Q�u&	 ��G�;��|�;'���s��Ѥ�E��D�����Y��؏�w��O��o����g�G�֢m�D����W(x=���o�e�JӊǙ�������A+}_s�4G�ʁ��D��OH�JɋBŐ����M�x3{��*��}ʇ�b]36�Y�D�C稼OTm�-\]u�
9J1ҞK�����=��l�����ޟk��O��G�}b21�#d��Ɵ�R����KO�o
������Q�m-�����M9/��l�|:P��ނ��݃?<��q�VB�RPT|��>���~۟u <�"����ayE�n��2�G�~�7U�^b��p�s����xr�E�sw8	�����?��ԉ���_F1�����T^ؙNT����^���:�j�p�l*A��o���;pK��("�ݍ�w��i?x3��F4brfU���0�1�ƈ�o�ؒ�� �*Ҭ�b*��Rp�03{�k0={z���%WA󆳺��톂��L�����Ǭ�h�i�Cj�H�M�fǩ��$�t�l�lϐ��ypu�=��d$�ӱ������5�x��Z�4���8���4���AZ��dlޯ�%���Վ%{��&R?��U��o���x�B�)�@(8~T��
����'+}�P��� �AVzZ(�,���_�A!Yx*A��]��d%̹SvOP�[��A�x��k�O�)���@�pLL���LS�u���W�6��im���������G��C &��9���YE}/]�o.$BAj4E�y�Q	�6�2U7-�a�sk�2R��P��fIYV���EW ����wzQЛ�����6����i�䯏��&�D��֩'d��
ˣ�F�P�#W�Zɦ���'Ϗ��y��rG�@0^"RR�XN]ug;����-�.:E��'x6��Bg���{P	����V�y���=���]�k�~�i���Aibrk'��1:n&ߧ��YS�):ByYg�҇�?[=l�A��"�5���!0k
�{�����o��H�[qiq������ɷɩBڃ!������.�.���R�u�X���
�:�f�ĢQl
�� ��Q:��\��[	H�Z�����}	��趤|�P<!�/R+$G�czT�j�>JIύ�B����@�dI�.�ܦ�&���xkC1rw߽]-���]�4Aġ܊��|Yv�0����y֩NX��b*�`��<�x��	��>~�ɧB����$,*�r�܉����ú��ۗ8��O�ASL��s����Z}1k�F���t�ǿw�~KD��t���,nU�[-�c�Iԕ���G�|w7��I�+J���i#�&��5JH�5s��?4���nJQt��uqq����9�T��Nf��C��Ӳ?r/D>�V-�E�Ț%��d�N�3�C�� A��~��yFp�A��9��>f�,kEC.^xA����S�ݩ�&�0�i{�r\�x���ZX���) ��Y�!<�1=	A�s������^)f��u�Y2�K�p��Z�bl�������gB-�sr����!Q{Я^��ޫ?�P�L�'�[;�v��1>P�ѣl��л��Q�αv`���&���7؉���˱�{¶L=�r���zG�ϟ??�?W78��7�<�$����	�gY�\�qss�]ិW�Z��C�E앒��������F�ɣ/����,أ�G��t�Q� ��9i
V���\����C1��A^�k�$s�	QN���,n�Aq"ߖOEc� �k�1w'�@�
ӓ��d� �x�A<��mu=Z��ˈ�A�����:uvO��B��hZ?�:ԝ����m�Bg��;�}̄ǒ�Y{p�S�W6��:���N����4�ߢ>[���QbX�45�KXOZr;M���.U(.VT��K.�z�/t�0�`�@mO$����i�P]Z%��YM����6vQ�te�[e��)!�j+��O��gE��uII��]�/f�=]���9%!&�@9�Z�\͉>��*J!J�za����m(]�r���2B(yG?��c���6V^H��GBˤ(��yp����J���h�/��K�
Ry�!�5�Pv�tb>�R�O�YP��+�qm�,�!��Q�ns��/��I�:��K�n����;�O��~��7�̞m�B,A��"�}GPIU����8�@x^�o!�M�2���2r&&���('���Ŷ��R��'$t2��n����Q�8�i5��B9�)�i��@��(���+7���h�y\JHNOO�@�iT���9�`�\�\�/jӡo("��~�����k��2�����;�o��^?��8�A1�� �hv���w�vr��L��أr��_Rf)Tfv��"����]aP|������@ ��>���y�6��q�5E����[J��z0����o�z��H�/k�cG�P*�cN�p���ÏF�2{�0���5*����z���x��8!�O����xpᅻ&���3...J ϲ���>O�16xB8F�lO{��;$���o�#f�����ΨSk���.��Oz,R����������n�u�;�y����(3�-,@�bY�؏陙{ �:iF_�
��kQ&�E �X�ޛ�n�3�<�IR��"f�i�^���}�V��_��e�(�ZJ�	}Fʕ(�ѥ]�q���A�Z
���˸��QZ'Պ����7*�����l
. #�CAx���H���}�`W]�G�����O�
���ԝK����ҹ&��� �NO�'^�}��x4Y�n�B�syP����ҌVηF�=�q��ۛ�ڦ8�ߛ����l��_tL�F�L2��_n�����5?��`������4C��E-��y���l�껐u@�zt�r�O�b��F�i���Y� �����F�3-7{Z�����\	f���U��pv�_|,
�y�g�<�B~O���q����uH%x���\�Ȧ���*�ל�ڐ��Lby��U������k >%'o4"onz`�n5[;_�n^�0�L�uyyt�8���ߛ�����=IpR�j�K�(�ʮ������!25��R򍅩���h�>d����1i5R&�ht����7��7l�ZG�'�S���pjg,%h�8ǰ��6+	������ag����V�9;p�Y��Ly��,�����ݓ����,�Y�#�a`d<<ZS��	��P6�nL�e�e}L�>#�Û���p3G~G���Q�*6��+0�2(�D3�i����F�0�<k��<y�,�$� �X�呣�j�#�"���ޫ_j�T���K_�#p/6�ŻM �{n�݁{X#$����?�ﱏ^9:�Ⱥ+��r?��OD�ٟ������=��I��8dؖ�ާ?<7���>K]
�۝���z��7Ω�f�2�\{]��YK�c�� ��i���A¶y>L�ub�%�M�1VQnh��.Щ�DW������R��g&��-���>�z��5K$����qa���FIF�����j�_�<Jc��,�aN/���p���1��E��~O�a\3hO��D*��J�[��t6���>��L��V���p֚��Q���g��lR������X���]�m-����c�j�3���lw&x��nP����I���Ѫ�?�����_�u���k;�(%Y�����sbs�7r8Q���t ��P��B�զ���c<t���PҪ�ož�*,N����)����n��`�A�*���%)���3�)*KVr�E�h��W�\�=bz�h㽥��!HK��3���%��@)
1�u�wWz[E
X�L���8�&Ys#�1%uT���Z�˞��-G�5��|�5+�k�7�=#O�V�5«+_+�Szn����t�$WnG�<��Ep��V��D�;�T������7�3��U��J�C;ִ�/B��{@�����ܢ�vL���0�S���u�^�%}h@i�Tpy�S(
���$������
E�Ũ/��<- SR����f�qK)j/����/�T��Y���+*#�0��C��0e}ߴWs4u�(�s�&��B���Ɗ�єV;s��ot]l��(f�����z_m�-T�3]e���B�B�,�	7j�@��̀3**.����@��`d����� ����2.�Mǰ���>��6(�=�1Y�5!y:;�O>8�P~K������k��Q��@v����T��9���^%�z�-��4xY%��:� ��c<��ᑛ46��!c�;*�V���[��J���7>��ދ�ܿ��2w���h���u��7EGfS�IU�,���	u�t��?[8��<�b�zs���Z��p?~Y�jc#37/s�&ݘK�����ڴ"OZ<���C��q%�6x§s���5���{�
+��qI'�凞TVLD�'"b�nGF���g���\(�1X�Q�p�����,hS(���u�Л�P�*���[Z�hm}�CU@��-�^�Dڮ��ݓȋl��ǘreؤ"@���Y�r�������gi����.�(����}�G03����S��A���)t}�#��\��N}$����qd��5sz\[�����K	���Y�~�dU3b^G�� ���{?^]W�X�3���x����b@�;�k��J��&d@+F��$�#���&�C���� _�@�0u��8"P��ٷ�?���'�*�#`#��L&��	�ΪA6J�9� H�ğX��2���MYږvO$B�Y�'2�.C�;��Q:Uܣ���?pFm�d�h��ɗ��\���X�o�����p�!"��&Xwn�����&˹�Y%�0�`��)G9!X�h��C�[���_L�R�,�Гף��n}S'I��(�D�P�e�M[��]�e��:�5�����`R%D�cgVN�������Y{-pr��<�WC��sd?2�E���H�l�'���w�����c��:��^��fӺ1����y���p-9ߔd���D�z5�7�jQ&//V▩Ǧf��|U��9��Ƚ4`�ӗ�b����[o�S�������M����-s�[,WX����$��1\�!sz?��\�؅�Q�ϟw��"S���[
��u�9f��<g�8	��8r��r�ݖm�D����J�,b��%�+�v�8_Ё�}ű�ߓ���Н��Z�N��h�"*0:���ھ@�!�7�$;�:ǅ�H|c$�����r\����?��A���4N�E�&}nh�V7�>f���Z�̗L��� �C� 
�芧�FȪ�X�����c���'>���~��4~����M�X����#	p�c3õ���w���p%#Ƕ"7M�ьR������͐��x��j�]h}*��a4����l��P�}	�U/[����xS���12}��_�=��d��˧����1[�l.�5^+}�2�Q;�Ȅ��vl����:��׿�w�qϨ�z����ͪ�,�������;���X~K���T�R"l�_�OÓ�o�L���m_��9��b�v\�L�5�ҩ(� A�a���FU�{����\��O�N�=��p4&t�kK��N�%��Z!B��&VP�����tx��"�,��|���ʼ�m]�+��7�:�@�����C���u�oR��PvOZ����+� ��(��F���"U
� 8�)8/w� n��:lZ��	��VwJ�Mu��tY�mf�o���"�:I5]?�p-���H�E��g���eyK;S�w�x�SN�����^9���~���Go��A���b�����>zm����I0Y ���冿�H2%���M*�Ŏ���G����(�lOk���?`��"fu�8\�E��w?��t��c,�}w��A`�&1�&���\�~�G�r/����H�4!f t�4�H˒R��}@&q����ݎ�.�C�<f�ߕ])���(|1�	�1�$���8��2mq�s�}S��5F�J����V �U��m�����?��~oetmm������� �60��I�9'Z`\`����{κ"��{~���[��N�S��[ y����yI��U��!stK�����#)���Y�$��)�(.� ���%��*dF�\���2��'Ŧ��o�޿�0���!H-&��dڋ��Z]���`$J��_8��22�tiL�T|��_�_������ݥ��7�,n�o�Ϣ�� c�� ���ȸ�����'䖎�+Wq�A��}씰��?T�%^V�E���Vi8�w���ʠ${����]� �Tq-k��6{��1Kf(o���jOk�aaM��Hy͛m%���T�7�Ӻ�[pGa�����b�8G���}�o��XX�|�ú�+c�+�Bfy�>��N1��5O�,e<�%��hn��^7]�8z��x�2� [���x���T���oy.�K�|y4������Ϙ�.��]b-W�S� %]�do�g9V�{����N1�����Q2|e��3o������%� �7BXs	s~D�vy`��^���إ�Ҳ�e��ܘ3�{F�>���/��>=Yߜ%y����%=��Z �ƌ�=&����I�ܽ4����[����(��#'N3ÖK��ѣ���r��?�!���O��3�6̘2"�Cep��/�I	x�qvGv&�����K�犜��Z�� A�����^R析��t2�l��]�f�݇W���Y�{z���*�>YA�jΏ�~�V�o�lk5ӸO@�m�&���~k��g��/��f�SU�[aC=�~�o�'����k_��,�0UiҞv�o
�%e{�-b���W�k9E0��l7�9H���E�o��dR7�Z�@��9����w���(�&)�ft��P�����'���Fe�N�<i������1l��*D��MM��W�,�Nx33^d�4 ��[�6l[�l���ħdsqL��w~���f����'Wo��苆Z�N�&��,���$PH��^��ͻ�<���Ր���/#�R�0#����X�G9�ԫW�m�ug�4r0C�y[O��F4����4�9s�%�,����2Vh��I�t�����:�A���[_q�y����Gd:w?yG� >gA�d��v�Cw��! G�	<'U��:J�/Ѓ&)q�Ò�l|Y��mV6��T���~���yt��y������
	E�`└��Sb�FS-��T0g�M`���c�c��&���v�w.��,����b���̴�.�Ż<�_��S�`�?�C��k.A��Ϟ��
��B	��cIᘙ-��.��Zy	¹�f$����}�=��e��[����Ãe��÷UUU�����7���!242J��lq�hn�Ӻ���ly�`�9�?�a����y��筨�����"��b�����90�����J��[�7��������[1������y��@Rn�*��0�(|�z�/�i��LE�&�h_m�O�>:j�h6W�3=3}{Gǃ��Tn\�Sޤ����u����9����u�9|�|qd�|4�Z�!��z�[�=�y�kr�[���]ћT�?ۆ�����;��B���5��JI �d�
�=�7m�C&�!����＼�g>�揿�I$5Rb�/�y�����u���'o�!�n��q�|A�r��	o_�☲`n�880{[�'�o)+#��<��o�_�Ei	G;���n��}_i��q%x������ԃ��_v�x|y���G��K��Y�V$�f|�[��Q�u����v��ʔ�Ge����_�DCK���c��ż$���jlj�éc��H}���Я�׫����{����o=��yX��X(��{]\[]<F�w������SG����F*6�܋��[�~8CC/*QLW��m_aʥx�o�Bg!x����"?�����SR�H�oRgG������K����,�e��/*���;L����F����ˑ%���)K�<*���R�o�>��j��lo�V���Io��IYt�xp%f�ڴ '{#�%�"d��#JE-�5Jv܇\C�8y� ������D$�9y-��|J�����D�OG$E��n.�J���VzY��67mm5��6��SS;GG�&���]��.���1P� ����K%5�P�g���yg��QW'RS_o����R^Z�ty�1��Z�x�)�@��P������.��8A9 ����wB3�xg���A�|ځ �p��W���Ʊr��֮�Q�瞔�5�ߚ&�h9�!�E=P���vg�~_8]~�3�Ǽ23Q�y���n�!�ڧ1���y����$:&&�=C#�{���
�&�6�_G��>&l�M����{�p5=����v�j��z�[�g�&��Q�wr�(���aPe�����b�%܋!�T�KQO�0G�Ƥ�`���^v�Q��;G.C�c�y_��na��3<=g{�������TS=�444j�k"��PY�B�¬�p�����:��{�T9���p�o&-_?
�O��֖�I��k����o��˟��1?-H��1�ܷ�ߍ�2N����l��^��������%$V[DSK�d����|���"έI�9�?��Ӣ�iZ��W�E4�?+��'p3�y�[4�N�����»0J�j*����ɔ�O��{�z�I.T_Gcch�e�Z:7�v 5q�MGs#Ύ��DWـ�_eA5�z�7�f����Wv�%�8�(
�ׂ���t#�v4|}��(?(p���XA�-���>8]��ޜ�����>kY|M��m�<m��#m$���4�{�,^Y�̔��eE�sg��p�ͯ���{�����V#�sI7��7,�S'���Lہ΋��4��_e+/���H��_]�t�9�K�<g?+%|��\����Ua`1<ʯ
p0��9ğ�y�;��ʩO�*tǛ<88辣�8��;X�L4v��z��n��q�~v�K»i�C���$Zv�RS��P{rޏ]Yڿ[_D������'���[H�D��Q���G}���es����=z����676��2�fAߞ~�;�����!11ۼ��{�G������ȑ������:G�h㤠�!C�N6��W�^d|��֎���r{�//�܁555��ՁD��0�
���P��H
G��pi�pm��m�Rs�-��#QQ�bi��0�g������v���}�⠼�L��Y�-)�́��X�:N��ꣾe���*@�Q�'	�t)y:m�Zdü	m;�J)�b��U��g�jȪ��*��)W���-���?ƅ�� #Ejs�gz��j�����6�2��.���|�����G�B�p3�˭7�|��������//-$��`�"�u��|�)�n�,�]ˍ���G�PG�9�,��X;&���|݌�<ވ���2����ν��0L�R�2OW#& �ss���j`oَ��/��e��_:[��.��i%�z����������-��n����{\�ܭx��˸�G�ߪ�5�T���gf�����#c�Zh��z��S��keg׏v�U���]1%����>0W�ӗ�s���`5�j�*9�Ih)��^�[��|RdZG@���	��j��ׇ`���5&g~��^��[��u��X+��6�.D`�j�NlM4��6����H�O��P4�I0�+�a�.)TX�{22E���ھ�8��,sNJoI�,�W�|�w>� o}�X��i�Wo�+|i��H��k��5����!�<?�0��ͧr0 �d�e�06��	w:0@EM5�������|:p<��〮2�09������4 �[��B��P��V�ǝ���@��]�紿��|fKۓ%E���J�|oFH^35P ��=�iqC�H�G����ސ�VJ�;�l
v�8?(	��k^��<���s�,U;���8����S����HZ�?k'I<��檅��~OzoN���
��%I��3h�qO]:|ll�B2��H�����fpa#��w�y���"9)��&�4%+,��x�t�lxU�ҹi�8���	җ#��C��Ȣ���]n`z(��?�mo�	ò�£*�	�P�+!DVU̓�����'a�$�±����"�bn�L���y����_�.�u�e��ޓyΆԅC�_��M)$��h���u^�!.��!0qM���LF�0�� �TS�)�z�sű5�Y�D�{�����F�k'�i�X���_��xć 6��rź/2�#m��쮞�a�!!}ǡ��M��ݪ�-��TH��Z��;�P+؈_���䶋�8Q��#�8QQ��ُ΁?a	b5�_��e	H6.��?u�ם#�Sp:n��u
�yo�ݻ����*8��E)HP������)�-����+�q��"��ri�����M&�ZC}vQһ��e�?�����S�Y�w�O|������?BN�O�Q��¹�$]Jٵ�f�/˥�����9��+s֕g���G�u�C���J([ȦP���EHFF8;��l���PvI%�y�93�Ȏㆽ��-�������p���y������~�^�.0�7��N7�t�TE����8��?�Yp��ޝ����~�IL��'���wg�ݛ/�Th܃邟�"}<��N��Ê_�M�b�H��\��m$Dw&N�>���t!�7Bk��G�]s�zo����DQw��D;tO�+�5$T�A��/�ۏw;���
�{n�k�.���!<b�m�584� �c9�) '�l���
K�����<*�k{<㩙c&X7@[N�8%w�5n���vi0���:�����C���oF��I�S�3=��{�+j�=��OD����t90���qp+m�X~��lA"���:�y��ݙ�!�sF��_*u{8��gu�*]W� aY�7|V�u�"�S7��CL���^�Q�O�>���,�~�'ާ��dgm�3�+�fVV�}.���O�);YӉ'ȿɀ3�;�wr�md	�̷cy$6���(��~oj�&���Ϙ8���|��.)kOK�m]�$KH2�Һ�nv.���i#���%��fb����srU$�i�R3o��~!��7���P�K�y�d��U�:zs���~���/R��v���:�X�A2�B�ٹ 2]">6��ٌ&bd|+W%�Jbbbq�˳ Kl@�T�{
�%ꅆ�Ʒ�P���_��`�*b�[?���(EQ1qm��[���R*�a-�~���<[&3qa�q�9H��m������s���;V �N��fu=��=o��3��%����1�ئh��LȊ�VB�b��I5�:�${(�*�{�ݫ��N$θ�q��+S�@���n�㌑Q�������j�/Z@��|.1,���.����-�y�F�3�H�����������mCE����dM�yܴ��7���Z�]�D<?��M��Z����e�JN�u��>6��(�ǻ��6ҊJ���Uq�g��oS���bb$��Q�]Vv��^OZJ*�7KB^bb8��}�e�3����ܣˑg^���SԤ39{��ki�o�_9B�B��8^>�j3淍2n�{����N��������m�Ý��t ���>�QB����_׆���SWpo^x�d�5fl� �"����#�̞_zd���&�;�Ւ�j@^ �9���ύ׀Y���"����򮠠�$������YV���W+�R����_��TUk>{�K�3z�U0�`�ڧ��6�f~�a�˾A$�W)��\T=������U���'�jc'L���]7V�A���}� ��%ր����`!V�h[���_�dq���Fɜ���z�r'��B�R�4�>�
��W3�1p#?�\W���rX��8h���P&�?��^K�����~�K?�7h|����D�nd�8��?e�cOR0#��2�����k�B�+�G{�uc���CJJI��	������������Z��>x�e�Qڕ��g�SOa��X6J���;����K,�9<���ҍ�߈b�x�������'(��ƷŁD���������T�mD��>){[�L����������w��{��&�F�/��R�;ż�iu�k�&����߉%;�w�siǮ�^�}Y��޹�}K+\��T2J ��IsU0ݴ9}v���e�fO����T��3+��Q=��X�0�2��5.� 6��Y�ҸM��q+� 7�*o�T���<Q�+�;e����`��?u��?L0�v�ػI��b�zy�dqu��C�%�.��>�/	=~'�T�6x[ǐKB�KU��Sv����[�q)�nzo����K|��m�8����R�`�̔��:` 1��I� V>�P�ȥ���:�| �d���Q1Z�2�u�2T�,99�,�-��l`��t*�"���t��~r���V��D���?Y2�:�^3��q��aQ]�I�Uy�?�F�{q���wl-�_s>:��V�_u����ڗ�0-�gϤ�u\&�(q87���R�H�rv~dd�?D�WJ�D�I~��΂�O� h�>�T�$uU�6�x�	/���� G-U��$�R~��z����<e����򹌆�
Z�'�n7�b5޿x�ٰS�@@��&m(AH�r [�{�� �3�9E!����B�E�_�1�wޑ���Β+r�8��`}tR7��͐v���`�o��Ԁ��t���G����tRi�8�#�(����t��ژ�J��')��.���:�
qzwy!q9z?o��C���O��'������D9�������>�����r�����T��Df�G:���s鹒ᱺ̱�Ci.���=H����xT^4�����,s..���-�k[%7�Vs��џ��L��ߕ�� �������t����6��HN��T��$�V�v�]o�ǡEX�#�R�]/0��GKMET�CV8�^�)|���|X��^�����xA��~G֣D�&� �.p��t	_�f؂��WVA�^���Є+�K�ܖU�i;^ի�1QSS_��P���#^��
e�_�jh�W0������l�z�`�h,+N'QV���V���';�n0����l
��~�f��V�#+r��3i�g��m�_�?L(��T�`�]t�j|/K�����z����r�Y���eF��f�l�gJ(����6�;;'gs��[�W;	4.�[7D�6�|���X����8zI�AȐ^���qo�N#���ys�ٞ�MT�퓿�x�C�xi@��ôz޽����ф��Q�X�Yէ�<J����F�?�����*�����j��W����Qɏj@O�p�
�	�\}1f��Q8�Q�r��ǩ���דy�)o�C�-�3�u��A�U��ؑRWO�e����č_�>��M�Pz�-w���ޕR��N�Z����Q�^�x�Xkֵ�|�]ҭ���,;/(y�+��������,������(�N��6�6�_��ɏY�eNI{���ֹ�+�(��y"l*l�"W5���$�fy�s��[��m�}��xA�����x¼��唶l��k�׹?;���+T����N>5��%���)O�l��g;F��5�x�u����[݋F�ͺ�	�T
�D˲m��uu_�wn&�QG�˅Gu�\�q���b���M���j'1��܁�YK��ҩ��'a�^��^G3.����������r��������A���2���eWq3F�/j@�V�����!�Q�^�����9	XA���QO?�-����X��bZ���U-��r�?.��{�=]f�)���sn^��k۫EGr&���M��<6l�4��kW)3+���ڇ��4�r�6��b��}� �;lY�yݻ���<�^T��^TkVҝG9:!bVL�?��V�-��K��v�`�ԍ��ŉ7)��}6i�J�@>�]5��c4�ː5���tw%fx�JD ��0BXb�N����V�I5tka���'ğ��\C�RG��ϡ�G��0�����/�[b��K����	'��\�R�����������D�,q��l�7o<C�3:+�X����2=�`�-��Gu��|��Pvx��t��(���x�]������⧟¾�4�J��|2��Y�o���T�#��/cK�?qy�s{�mA~�i���q�i{�;I�t�ƀGAn���>nE�����仩�o?��xM14�R�*ȽI�K��|V?U:.��O��8��3?k�}9�X�r�ܡ��K�t�?[�h�U>�~�bp�i�Q܇z�rq���n_��:B�G�M� ��=�B�&�b��f��.����QCp�G�Rr����@UC`�䶖�k)�KwJ3&sa�X3�]_z�y/$��7m�R��2�jd�)h���Ae��(~q̐=�w���|����پ� 0���a!��I���O�,t�j��SQsHTO�����E����|#g��1|=��������?UԱF�6,�x��|V��5�oWď�+�N{C�O ��"""��3��G�vI,\zO<�\��~N����+6����_����N�R*Gm&ښTJxtp�0�����������ALej��4��\��N�Vo���鄚�r\��fC�--�~�ao!m�u�m���JK[��� ���q���iJ�,���?�3<`rtr@⣗�C~[ZZJ ��W�V����&�u卦8���!���Z��@~L�[�]�;b�s4���n��ė0b��������NU�_r�8�+1����Q��\�5��X�kUp2���"�m�{b>�V"������p4k�?t��B�P��+դ�Dt�4n��`���(�Л��Q*Ȧ��ײ�A	\��p�@�������W�<���w�4���ͽ֌Pb�G��������S@$����k�垺K�u��[}Ɲ�i�&�u�3?������'����(��
�z~BOAZK�[)�"J��[xL��I���s�,i ������������T�����<U�ҋ��Ї��V����dϐ*r��&4;;�junD����Ld8\�jPB���v�A�+���u"|hA��gE������7Aao1�>Z��!�+>����L�f/)K�=v�!�AJ��O���,�W�p�T����`SV�b�R
�_>l�f�{��'?5M� i�����_�Ik��+�B9:����3�1���<�$8\�������=X�ͯ�����P�-�m�W-�D�6��@�g�<���𖯺c����?G�,��?%���V�"{Ž6̺#rQ��yq����(S�Χpé_bO4g����*OlC"8c��Q���!�j��;��1E��*��\h���[5B����L
�{���e��а�I���˾�*j���(:O�7�,��I*�{*�R �d����͏r��R�nk�e����4����	��QX�=�E{U��7��j��.��'����@/ؙ�K�Լk�"E��Z��
�;�G"w0�}1�0h�:V:!�a���c�_�&����cep�8��՛���2kh�[]___�T�a�Q�N��bl� ���h���i�q�о�m�:1��d��k�����[/2ֿ�`\���+�A��A(�M~�
D��j������
.��O��e�����Ԋ.8w��睇�!Q`�g/���ppe�G6����F[��6������m�6�Q��Pg�:��o==T$s��ML��.g�½!�7�:�	�M+x訾'oUxk�N���I�".�/O'm	ǣ��m��=�
_�]Ѫ�{o1�+H�~�V�Yո�[��z�:8��
���:�-�}[���+M�s�ᣛ��i*G�˓�;��Z�%w�����Y�-3'��~8 ���J��0\��ڞ�E�&� �KNu�8b"�����ٻj����eK�"��yߑ��;4�{�w�?�v�����684�F�q�9�e_v(<&��>�B����IY̛!p5<,��,˳i�=�#��o|{4 ��ZAu�jbw��N��$�����^�����G�T��h{�1	���I�UXt���G3:�Zj�[[���ђQ�cM^_�QTZ���TT�����j룇&-ˎ����{��U�ؕ-;����m�d�7��W��F�.��UA��.��͑�� ��D\ϾƠ�[:5=���  �Α��`e��w� ��C�o?zI�P��M�r�[��D��˦�۳�$��8w���Y���n@_h�rXIԓ�έ;ƃ��w26c�Ėdܤ������Q�+��Ӫ���_�D���-o��>� ���t������&.��``?��-�h�Zb��s-CԀ$�X:\��P'�\����#�|����D��)��zz�SU���j� ��`��t��i_���LF����8�G����߯q�s�;r�^yNP�ӸR� ���q��z�����mm<c��,_�Q����c�F{����y_>(�s�<����l̎'j����TҸ���&#>�a�I���C��^��~����r:S����[ uL��~A`F��		�z��7���U�Ŧg��7K��PP�����f��H�q�j��I@m
{�1���ۍ1���X���&�q�϶�$1��j���L�
������J���Ι��by0B[n��&��>�,�E"�>�4ݙ�6GCwg�tXϲ
�)=xÙ �X�e�Vt�����1�Kךm@��:�xVv.ޛ�#����������D�v�W[6� ?pj�%�v6.��žVdzS^s{�8�𫨷)�ŀ��);����Vt{ښe��e�W��T_1�,�D�Iɳ]ץ<�}�z�����1;��¦�T^u�C���w����J(|_n;���B����F�n�j����đC<�>)���G�u�W&#�2qlT��:
�ꁷ��\ݦu �kB��ҋ���q���mQf'��ٔ�'�5`�/�3��Հ�1����kx>'�����5���;0v¹]|��<�/&U��}�۶��:���]�������0�A�������y]�_���,G�=����D���6�����d�A�55u��B���Ə�+����m>|�pitq��cؚ]���1���GH�y���ε5���<�=E-�;�|���\��yb&��N�����tS��:�ӡa^\ǫy���[�9@�#}7�¶')��:���1��&�\�}z(*&����Q��\ɾ���cd�s&I���\ӯ� ��w�����&1��^y��;Ys��v=ֈ�ҹJH���?������F}��]Ϟ=�c�%a�I��FvvN%x`����ҭ��1p>wSVO��{Uu=�u!�Սj���%������iP���_��bjZls�B��(.G0�.�zU-Yx����{"r����]�Vlv0VN��y4����d^D5V�8�&���hz��tѵ"�c�_��c��
<���\8�4�>��3b������%OU���kmi����.�?�r�d�&���@6V]gy���v��g��F�~��@����l���V"�)4��gt�qoHws�D�i�L{�TM���#:�ڼo�ρ��z	lJ�[_熽h��7SݩҗSE�Ӥ�wf����[��x~���v��9�P^�`}S�jZ�hD�i���JF�E�C^����٤�����h^����*K�q[e^+v��߷E�!V֋���߸?NW��f�G�W�7q��gg\�dK���9��W���v�u�^׆�~�2�^c���OW�M3�lM�m�(�
�P�V64��E|r8􊮘��!��E�΍_K)L���b	�Xn���f����?#U5�Q11�"iR&%r%��>�,�m�nF�ش=sI��y{P�������CR���{ͨߒ�1/���P������8�j�G�k.�� �2;�U8���;nw��z������'��1�aP�P���#����)�kn���$>��(�rk%�r�鋆(�>}��5וL�3wV���;{�/c`�֥����� A-�{�ޛ~���ٕ��	��8���������ɔ� �[�qq�������^�;�m@�K⧭xK	j7`��q�\w�r�q��)Ks�-�Z���a1ٝӜޤf;7i������\�M��ĩ̴�L����q9o���6�m�<i}��_pSS���b���Y��~�'e7=w���^)y�ߜT;��h���
R&�=�/�d���D���߁�%�g#����F�T�������V��k�m2D�%�fQ�_%���m:s]ù��K��)����zzzU[�?GG��#Nwu"�,G�{6�O�{�� T�j9|������y>�ϔO�&�!�o榇�7��E�(5 ��Yvw��@���I��;_58vb�]F^�l\F��2��Y���@��d[�{�'3��i�un���M׎�r(�֬�w2N�^U�=�n0ڦ&3-������1KGҟݹ�.��N��1���/�2c����=b�o�S.�|pa _U�����J���՛͵}��]S�g�|7ȏ��7���1�T�������m��ӯ_n^�����x����5����ޣ<~��7��칺ۿ�>��m��u�����ډ��7�1�d掫g<2`�KI.�U�y�z�T֫����`�?������;���ƪPBS���	.X���5��$��5G�fƭ,����@���0�i��h��T��ȕ�b�j���p{�2ngLy�1G q��	�^�P}�|f���J�:�j��qX������*R�Y�K	��r�[R�<>���"M��a�O\��Q/'/�R�����Kq'e�4>s ]D���-���3119�X�W��37��l�rX\⋀����ܞ�KߩJ�蕭4s&UHz�]AR"�/l�`ط������çR=.c�ymmm����i]c��M��珛�9��wq�=�p�%%�B��8�<��2O�� h��]�`.�<P^��,�ţ�W���H�ұϴ�l=�]�a{��S���sx!���IZ�7(����������#/CKf���K��-�k�~(��8{A�H|]Q>�:�RTCV���Xq�,O]511������̲�������.�Wn�	Q��v��G���h$�\F�h�=ijj�z`�|W]]=U�fz�>6���W�!\ⓣ�OAN���bf||jT79���-�C�d ������]7��Iu+����:�vX�"��>�B�����1�)�h�����|�ΝS@l��Ċ�G���i@�������mQ��Tju#��4x���P4�4�:�K=��0mV���u����M�z��?Hdk���l-�,��eKe1K��ҁ߫l�Z���� UD<�&lߍ`L��,u -Ҍq�Q����	�TaS��ȫJ��=�?�_�,��f�����a�dWkv�ڎ�A���ч t'n�9ȜR^i>z��(�Y!uԀ�n�$�`mr�J��gl����I�X��f �}��H¤|�p�����^\��g�K���!��k�/�\��L���Xb�_2 ���]ȨϽ�̴9���@}�w��M.133�;!6XX��C��Dk5L�!�ԯ3H.G.��l[2�/�2p5��D��U�VەURV.�,B���1����'O�e_����L���Z7ZG8��p[饐�����Z���t�lF���O/W��0S��v|!.S�1���E�!L�d��Ɏ�<Wh��kk�����w`;'���K�Ye`�?��D&f�e�	.��Q��@w�/1���,OE�W�JW�!�-g'O�<U?����;]f�K"��CH�uׅ��h}�=i��l����V��.�x�[8��۽��e�.�D������%��� ����}Z�-���2�4�B����|��j�`�Օߕ��g���>|h83�Q�2����ٰ��v���꧹��jr=��J0��R�l�������/--=���6y�|�JfVV����r����W�x��Ek!�����?EN>�ʞY�fe������}�V��d��7]�tؤ�G�N�ɠ�N�?���2�nI��ޣ>S�dd|=�pu�z�����5���}���O�uu�jjj:���,��vU��E�$����'������#�$�������x{jû|��o���f+�p��:���,5�����s�MA,"��w��_�}w�����d	�S��}�w.�=���l�H�Z&"�����d�~���}������%�:y�B���~0�y��(tL\�qZ^Y�x8"�E�!�~��,�(Y�o�cn:	u՗��Td�nmI,���57�����9{x���Q������EB����˟�����(8[�[��A�豱��|�)�� V�����AEN���,?���O ����=�8�&�4�ɞ~�:8���qΊ��cà��i��[���,xg.��x)n�����%�}ڵֵ<u�r�;�WJ��`��l�Z*��"�$�����3S�΂�#�F����̬ �־~\�JKf�k�w�����p��p=?Ԅ�#���O�Q�M)��h���#��"�=׈~�N�|������V��d�lg����*���ٿ�f�_�;�Lm���v���A<	�����uz(�M�W��$�T��o�o����#�55q{p�Ş�k���ZG�@%����!��,w� �
��� ��a]����H����)���T^{,2���������m6.����l���#�SZ�M��0?;������۽8�=i	��"ps;���g;:R�����!԰( �W緁�1��oTH����Q?�|V[�x�ؾ�C�;���CEM�GA���3G�>���CD���ڹ��ǚ��1�"�����U$���we0�+!�ّ��HnTG����O�\�u����]��;�����Ilf/���@T���_rAt*�d�X7u�8�P�1{�r"���҃|�+k��l��\���EMd1��C���������ײ�rt<:�TwZ��B΄�Uq�IڠL窈��(�t)�:/Z�j�pJ9��j��ׂ�¬������K��b5��VxE'#r����84�5���]�L��Q���4Il�p9󅊓Y��T9��w�����t�)�#m��;�;<&�L%|xH�����Cv&)I�mv�gjXa7]��1=��#�l�±o7� �sX��&M���C�ޑx��c��WY��5�ޏR�7m%id��
�!�_kVA�4׉��,��]�u�R�@{�I���x����8,lI~9z��^]qp�$�ͣ���78o�����d����g��Pj�
�K�D�}pg� ��X�"�lr�"_Ѣm�韴T#d��KA/fI�.�|6&Ue�r��%.�T�Ti s�C!���w��t�>�x� ^f��
XK����.'��ܢN��Ng����%��r��n��G����O�U�u��Ύ���e��|�JUg���gz�:����l@����ظx4�:�u��%yB�!.�R��J��T���
�%p�w���e  �i��(Պ�CS$������U�Wu(jn�oܨB�5����Г#�	+�k�������P��wo�(��)��d�jW�x�?�[�6���=cZ
!���F8}��H�=���TO�'$2�z���*����?�VA��@h�C���c@�{oRܝL�۲[�<L��[�譊��E �VL��Up͡� ���d�RS��*#�>@�o"8�t_��1���_�wxr{�@���GY-E�N`j9����N�|��_����Bk���A$t|�j���v���W"�2N��sﭏ��{l��|Drܛ7oznL6�~��:p݌�����A���^J=�;w����+*&�z��f܇���i�����QI�r=(�3�#}Mxؕ���$eh��(����fQ�,��%�ث.�Ш�,��=~�AW���B!�{Y��)k6_<Α��[�ML<�oʿ��ɓ<����	c��>k��m"�KLL�M9H�1��r��P��/X��?2��mq��_�/T0���������WS��i�Ke)_T�X�� o{�.�"�>�Uz�T�U��x��i������#|�N�<���w��{w���8���e�b��pA�.3[���h�����j�k�F14F	 �4;+�<�ya�cV|�%�$N�!Hq�լ>r1��#G�J@ȵﮡ�w��l"B%��^��W*��P�z1Dqt�>F�[����/pT�_���n]B^ N��1!�T	�1R5bbD~-�ލ��j���Ji�Ԟ���C��KX7��"��<�[$���XZ����z�����ݽ�x���vu}*����h,�u����+b���aϸH�i��A;�|R@AO����z��|��O.�ǀ���
��N���N*8�/�����ܔ��}�/�؏�y�n�E.[v�M:,�&���`k�m�k��K���T8�'W����62q�Բ���tB��]���^��>��I�(HT{i�aib����Kc'�Ͻ����j��c��i�<��A���ҷ���ڌ�_�``�_+̻�d.^�1n;� �m��q����TC�,�k&,"��u�������ǒ�`j�5L���[�$ p�^�,Q��
�b�{�F7:ÄVG�_�ɴe0����x���d.��]W�f�#�2��;���,�$.'����@g;�q-��cء��2yڕ���#KgR7�����&�)�%u/���(S�{Lv����l.��y"��T�o���8�x���MpPA29Q��M��>K�����'��u���O	�K@��
}�;~V.�*@>���G����u�'bY��zC��.϶"�(��+M���B{"w^��V�A���KR��)\�ŉ�w�s>��+�.�n|�nBE��'5ϸ�D���8d��a(��IC�|5@��:G���C��.�O䟬�	=1b�Z�0��' �B��s�wԧ�{�����"#����%���qe�q d_4���g��m ���׏��޲R	�)C1�1_��f���r:;;z����U��%>?��zL�bD��h���bMLLd[���3��;�P{���8��<}�����R� \��`���c2�:��?�4�"ʽ�Bt������u_�3���w��ܛ����xo�*��m�WI`�����ﾸ����W?��X�Y(Y���e@/��yo��S�����vޤ�� ���8�q2��-��=����t篡;ھ.G2��u�o�'�>qr.����k�	ۚ�e�ݵK�s�6yް����%�� }E��ؚ�se)Q��~Y��<ʟ/��/o����5^C?�����E��~sc\�=�dt���5��}-p[������(���]�d��A��<,���W}��xh��q�4��]�aF�y�<�|�"�́!�c?����1	�ac���MGfq$�7
D���-�,�W���jk_!Z�a��p��}�˓=;d��W3N�����9����v{Y!3ߢȸp(�:<��\�|�ߺ�"i�&?�zo����z�i3�WXޤ��U�:��-gj27	�s��
5N���ͺuX���ҲM��r-��
BRv��Vʉl,�6��&�����>�У+��̼?ނ&�`#>�؟���||���x�ΐK�U�6��ߨ���T��U�y�m����郘E�&b��3�����qi�e�������_�s�c�>5���>�x�G�i���|AҒ*ш�}�M���ܣ��YA�*�9z�h$��
6�QO��P�s�=xF;�)�ؽ��D�5�{��������P�ˠk��P�;RO��b��=��[���Y|@*+��?�AG��ׇ� '26b��S�znF������A��:MC�ȗ��2'���9���J�繋��1�.aKo�^;Gڋ���șF71ӑ&���'$���W���|�����h�7�coM(�p�[��H��W	=���i�g}�C��D�O�������v�'e���s�jTLw�ܴ�<+�G�E�1,�A^�=O�߂�^"�MV�?�7�&��.Ad \���/�$��Q�eD�s��&s�#8;�0!�V嗫b�e��p��Sz�ެ���)��L�ʋ���wz�=�T������U1�6w{y�]Z���d�n��D��g�r0{����?k�q��ۄW��Y~ N����О�Xu�n��i��	oIy��r�.����/�^<=~��+A�J�_�	�����{�G0�'����۴j\��3��6O�$����& ��Z�7p�,����1��2���9�Jq�7*[���� uѷ	s�R�|D����M�1O~t� ��<� M/�w�+�&=�!�ܽ�|5�7��J�a~�������\���<�p����m�,������fy�ٗ��$k�h���D�[����4��������$C<�UO����m@�u���u}t�<�e�����"�Z	7~xm/0S��c�@��&܍�B�<���%�.�p�?����"�A7�9��m�:ٹl����C���te�4hkA�����2�jw�����)�f�����ku����&�l0� d{�����se�wy(�����m6�v.��.��l3��v<FkN4==�>���� ��9셍���b��h�n��/���q--�|�r�D�â��z�D�q5�0c�d��/�<�K�*���ᴩ4�8�"���@XcA�<p�3C���0��3iqx�IsE�g�A�#�ר���(�i���S��������g���I�1��m��A�_�`�klJ�㦌K�l��70�Y�h1�X2���^ƬX]��=�5d$3j�0c���hӿ��ၽ=�"�C��C�h�h�	Ԭ:���嘣KKKe���g�O#l�.�����SR0 0��g�Я�l��LRg��(yˮcH����,F��i���Z�q��;d�b����<����n���s�ܡ&PP�8�F=��k��o��p2{��]�E]��	�����G7 (1��{i6���_:X�'��䙥�u/�#x`��z�߇o��W������~�;�Rjz|�ֲJR���((-YS�e� b�]�*��/�Ik�n��j8����^���14:Q룜�� ���Ǫ�N���������b,]�1,��#����yӊ5�}_���U���3�K��?S�j	���Ls:"�y�0 nk�E��܂��X�T� o���P�7��p�a�T�SN��N��=�>�Vf4|4a�����L���&��J�86��%�8�)�I���-���y���<��֤�i�0�Y��@��^����u���2��8�<��x��)�rD���e��.�`t���\�$ڏ��T[8�^������7�V3첽������ruNZ:����CM���[�[���cEi&h�"�wê����R�@��uh1�a���7��\p��묢�;&<����G[�W���9ý�u�����d|!]��i꺹r��YGiN��^.�������[,���|<�ɵ���e)��V>��u�v��_��W�GQ�3E���r�
���d9����m�N��n�z����z48v!�}Te�pB���D��=�z2{'P�*R0����B�.JݺAUa�3?�V��
������DP�[��^g��X:�ΰĢ�Mzu�/��ͳ�G߅Xb�V-�UC8Ƥ�#eoOSqkR�1˻��X�?������5���<4�l���v�4��b�'� tvnn��RȜ*�7;܇Q]��~� �b����䛰5;�
�����x~��l$t�T���$��5��坖uI���@'Q:����l�ʴv�_�ت�.0�f�j�@^�o�m�.$<}��%��y�Ȩi�T&!���-�J@սT�D���I
�FL�T7+��'�-ɽoU��F�樨G$ O))�=��~/$Z1hM`������D��P�����2����4���;p�[��{�g����A>1�=i��ۉ7�iFL9�C!���̞Yj�P�5e��L�F�������-���Pn�Nx�GL0���}��5L+mn����x|íb��;K�D2�Ġ�p������F_�Ah��'w_�����Z�T;�������,�8X�,�>p�iY���7n�i�/7??@�t�a*!�P!5�p�׼Bs��?��s�jNf�ϕ�� ��Ƈ�9��X�� L0�J�6�F�����rmu׉g~��"�7R(���nhDۑ/g���dH�@�)#H�;���k݉��_U(����n��'M]��a����]^��'_��R�M��#������]t}��aC�hzz c?
�_�wXH^�.�ዂ_�9��D.l�J@>�/�}ت�V�4L�U�=j3$��&T��,t�ѹ�o���[9֝.��/w�U;�v��s�b=8[�♜7��Q?V	��W�U�Y�ZP�x|��������������?��q�����>��Nc9q����sݜj����IU󳊆�D��	�]eQ6�,x��6fLc�j4�/i |>ln���D�aؒ�l�����J��1a�Tˀ�����Y�*Θ�ʾ��m�^Jhh���H�詈�d�j��O�����R��K��g"h���s;�i0}��u���>z�W�*�H�Ɲ'����h�s�o?����^��@*�%�E�{_��mddem}�&�o���4���YW_*�<iP�v�+���o�"Eg�)E���M����KY�=��?��R&�4"}d{�����7��V��c���(��K�������l2���d'g\* ���)mU�Z ~�����VA����;�Ʌ;3#��
�s��&�����\t� �q��Ș-PX�|���ѝ"��ՙ5�ض��ԟ��%N�뜞|� �u�x���D�d�����Go������	�������{�����5*bz8�eb���R"�0ziQu�����0�Q��b��H�͓�������.��k]u��ǝu�KW���]f~����Έa��tI�fq�'��/+����&����q�44�׳z' ��mUf����0W���!�z[
�H̙��.w��d\���#�>���JJO��xlO���Z\��cߞL𤐽{����W����f���(^ߚ�<��vH-/+���$��n���[�la{�o��{���%r�OY�?�v|�F�?I{�B�;~ ���[ѭ�q��&�4�o��YjF���g��S�r���Z�$��P�2�Շ8Xji��1IvĿ��67Q�t��ͻ6���͓D����V��ǭ;��E4�S.ww�i��?,�Xv�V�*0em���uu�'��}��*� E��!Y�N$X�#+:�=�F0D�K@r�I�Qr�#���pw|K@�Ge�����x�����(!��E�M�3D*#YWF��q�k${��ɾ�.�ȺHH��^��6���5��V����xxؗ�=�s��u��uYm��A�|jt����D~��ƛ����ƃ�\~�'�|JP5��6s�����7��Z�/ �d��]8���9!H����i�'����)ke���	N��y�_r�&�6�֭�mD��zд���=P���\�ᾱ���ǈ�P�ڥ'a��ͭ�`D�_�4#7g<�i��?`-��}a5��>�YO@7����<\���3lMm��`��S���*��IZ�6��8����W��ԉ�l?�	�^g�Ҫ�V�����H�ݙ��sÅZ𑉷1�S�
6���}<����O���R9����FJX;��L����bV��ٚ:�/xM�������M�|t"{���gb&S���te�Ѯ�P��������	B��,a%���<��)Hp@���~<���u�����NR$g���n :��4���bT햹�2�+5�'��~/�d��~��E��
ka�Z">�[����3z)��:ŪkgG�Q�-<�J^]ݽ0*��,��w�����q?b������}ݣ�[�nǾ݆i
j�J��+�%7ا�����Qv0�~~��+Z$j�p,����H�}�zs ���p��f�K����޽E���cF�{"���?�>�\�?C��5�X'�%Fl*���7>|�A�*��ھ�G���������O����Y�:N�i��;o�4�F;@IJ��򒪊	��s�
��	��z����y������״�e��h���f��FFc�N_���fV�~l�me'<���Q�qs�JE�༎x�[ )�1,����ZgbW;U^�1V�Q��H��8�S%�i*|�'�����eC�G�P�p�5�?��Tz��-:6L�UT�;	S�;�۱��)���=�D@�ږ�`���n�-����ȁ-8�:�܋u���~U{s�k�����NA����V'\�U�w�uL%�yLF+ϋg!"q���7�Ŀ�0E��U��uߴ�}��염���vOZ\@o���~�ư6����r9�HzT���k��9����D�I�N�34��-���8��N��NDT���HT9@��&�+ۋ�̧|���Z�H`ܓ�#���-���x
-�b��D�I`�6��{�B	�K����I�3�����^`)-8t����6(�E%�29y�OD������U5�~*RI�RG�	�w�6�$=�&2x�pKp�ޙ�24r8eLz��5�U3Myp�x���x�g�������F�B`�Sr��Iu=�fE�ӗ�I�'�����>���� ��9IK�g��y��6̜b<ot14xϘ��C�[ �Jbr[j`���S9�ן8\�aY�Nֿ�;j���[ ��=�\,�>kx'QtZ������|�;�u�
�R;~�Xo�[����K�"p��b8KMH<���)�K�����|����%���+�Gx.�&�����������zߑ�D�n��`0;���{э�?���F�TLY�_׈�v���>`y�W�������N��:3��/D�7U�_�n[b��zj�RA�g�F�����~���]�)�ϵ��*	l�da~an��7�hTy��^�g6����2xn˸
'im�����a'i���3g�e���`��͖U����$�((ɠ�r��S���U	.ٯA�b�6g����/8�9|���ǫ��n�%�7��9s;�u����V5cj�~��$��R�3B�V8���{�éhu������c�掤O�=��~��o]&�p�'�:H�{�ǡCM�IF?�0u�>]�����47�mG[ݎ��^k�>�UJ�������+ˋ�mǢ��z��q����oC�����v���jfEܽ�+�=���|�у��^��_#z��ܚl�Q��Ͽ���x
9^��� �^����V��gNI	w��ಌ�3�NDssW������2(k��� �i}���_�sC0r���y��� �d��~�5*���1i~�+u0������ s�ݴ=1��u]�z_�OD�s�Q0�y��n����ln��e܊�t���zI�#�~�$�k�g>�� t��ڂ�P9�J~�́Ć�h�2��lFcS������&��c[��.�G�Y��z⹀�Ŏ;�k ���o.�� �l�-�(��d�Q�y�ȕ���7Y�1;�:+&���k�"�V���z{�T�hJ��,{Ȓ�F��1i�,I��Z�~����0tmn��H�T�QϠ�2������e^�m}��V�B3�#�r�1$i�ۡ�=C,!Α���ځ��p���7���ƛT�S0�XS�����*} "���f1j����=@zA��p�P�������:�ܼ6����}VW�ɲR�S�u8r�7/f
���M�	Y�Z�B�ùT۸�C�~�%�Uܙ
���ݾV�v*�l\��G���?U_n����pV�]�LW��y�p�6�y�3��TGֳغ�������}V'�b�=������ ے^��vV���q���F�9\=]��Ǜ���:��*�m!턶u�m`\x�^�s�J��k
}Ѵ�Vɹ����>Ҹe>fW�t/��6`��^U77+�z�DMMmKH� Q���)�n��2m/_;�?��Ư�hٴ�zr���f���嚪��6fe�c	������c9}�O���d������	��P�1�B�U��Л9�Vg�����*  ��K�k�����BTTT_p�'�+�R���+~���+�>�Z���~�*..�/۱��m��-,�L�"��z
�D�5ɪ�h5 _q�+//?�����N�ş��̍gc,�认��CwQrq�q��Q���)�t[��)nf����f2���3^��m��UNp*|�^?��qb�CÛ5g��.���i�c��"~ Bt\��B�I�Ґ��V�_��u�֚j���Ό6�)�W��Ln%j�/%DEC�v��n�͐F���$�.����}sf\b����
3�9�[R���5A����$���GMVI�N���-+�B
�S8y'NNI��z�
<�p�����-���?�N��S9�v��uf�D�;lλ�o5�7�R=~5��
?gH-�8BM�qs�Ip�-����v��Ru�Q���cdB�A os��5]��ocI^7�Zgٞ��V�=��S��:����˛�Ξ�}��+����2$�#�gK�m�~��U��2�J��GU�0��:�����J]����M�2�<��؄�G)���Š��3ζ���BWשX���l�m�=�2=$�K��������@?�V?�m��~Rv�{'B'm�9؜i�!sn�@0U8p�dacc#�B�É*�����l̧	�}����������ߗX6�
�^�����1�R����#�W�9���`��Q��>�=#*��X�c>�x�����b+��E�+�<�:�<0���@;�ug�*��싞�����l�:\[��h�8�d��v�K7t�<\�A>��i6d��q��$]Ӻ�s������J*ԋ���ܹ��d�=]���.�jv,��%]sY����C������q��B�l	���sQ�K�9ʹ%.<u��������Qr��4)B�v��=���n+{��&��2��7m�L�m�3b�ʶń"�E������Sљ��AZZ����z�ӊ����DYTLlع��׌��羅������!c�Y��������jDsHp�:a|����8�������RX��y��́�'Y��Y#'�"?��͔��4�*��x��6݆�I���RYYy���8�tB�����M��v5rI�4��yi��7�_f,y_�/<}Qy�
շ��j�`�׈�/�{��s��9R&{�g]��t)�W&�ʎ
U<@tF�Z�o�4e�!�����nK ��e*_���8�(#���*N<_5S�����g��|����X����G���r��*!^n~O��/�iw���T�'���2�e�pu�fU8��7c�Z��S���=�O��!	��E�S~e �j�͎�OZ�w*���vǣY�=�Y��	Wם��f����IZ�1K�A۪���;�n���Dz���e��ñ[��c����Ӻ� ֺ���S���ӷs�(�3���*߾�da�]�m|�,U����CzfNM�hN���=$�8�{��rȵ��u?�s�z�����B�rӕ��H{�y�VPљ�洵�32�!FGS[  ��H9Q����	ݙ�i����g9��������@v�l�����J�v{�\f��k�.����,,���ݲK��6��8OЁJR�*����2���b;+ߥ���u���=G�Éҕ��m�����RY	��fj��G�~n�z�:��DY	�@g�T�b������[	㑟�nm�\�8|��ƙ��On�Vf��x�d�c�v�oL�b�J�S� )=n�R<e����.η����1�k�34:��m�;���S�vf������#+���e&)�E���ǲΩ[���0�z4���	|��^�_/=i^1�Xvd��c{=����|���l����腶S���ں�Ku�����N��>uW N]%c���7�6��/IS,�.'-��Â'�� �k��1pI�6UG����vO	
���J}�5��_w꽿�� �6/��;e�5�8��ƿ�K2��"��XU��e]8�:Q�xM��'����jZ�jh��j�&D��K���S���G�SAx+� �kڔ�����c8��õ� ��yk\+�[�(�3����N/g�7����%ܖ%c�Wm'�w)�%�g�Bv0����P)W2�nc��Ґ�]wrDFޓD��҃R�h,�C��g���:��O������i��B�,g�be�ј�ũ��6.3T���׉ �M�%�_����<��+��qJ��zR���y�'?�G���E9~��բ��U�cK����������Z)�=I�p*�EX��P�cojaV��M�*�#cD��&"2퍹?M��Vt�aʭ���4�o=����Խ<��C��&s�Ȣ�5�����j�p*����/�b����g�#Rq։���$o�����6���Z $O�S��:�hy_%%�� �~�B	���XP����Tu�v��V<����LIu�]�e�{k�����;��Z�	������1��R��|x���3_I�1���[j^����6����8�*���-���_�2t��[��z���o�@8g�ž��C�8�RܪSe��RK�r��M�S\���qK4��������MJ=�T�+v|�Mj=�b��~#����� ���Wn��hH�H�ib�B0�G>�ͩ�,1v�����b/���߹������J��/$��S��Ho#�7���ܵ��_(�e1P�c_z���+CZ�m�(SO!�lz�rЮ���d ����<����_�`J���N�0/O/}�T�Dv�h4�;z�>�a�"�\/H����jk�}I�w��Χ) ��v��{�6��4�Ѿ��Ѷ-&U�٭-q��tBv&\��b��Bi=�P��5x�[�F�	Ug�<o|z�b&�9��C�Y��G�q�n�|� 7���6]�El�סw�c�r�ǯ -�L��9q�;Y��۝�;<�}���6���Tn��f�M�)E��1�7
��tk6���:�Qɷ ���^�w�#�*����Wk��qK� C��9L�I�=齾��W��s��(~��ĩ���>�zrL�[V �e�㥒t�	N�gcN k���R�#��Eס\L�R���A�����fkv��\%��3>�8�KwbA�Q{���}���_n~~1�cRP�A$�.��Ս�RbЉ�:&�e�\�\�o�x�X��>���K�JH�!�}��Dj��+��������+�6ޝ�{g�s5&N��s�0cf(���hI��0�v�P��]!����I��U��N�vtU+*��P�R}�W9~7 ���XΤ9Tp=!���*Z�/���:����E��U��k3q������6^=�'Rʥ����iQ��<��f�V[�WZ�N���y<��p�:�u5��s��,wy!�f�Yb(H�!o��"͐]��r.q(W�M���5u��D�;�����ۻ���r.�n:Av/�ĺ�,Y�*-����I?9����m�J/�Gu��+VRm���=Hs�R����S���t�u��U�?��^�af��J�c{��:��8	TC{��C��u���#q�Y�'���g����E�~��_�SsM���C�iB�v��2�$�c	�����V�/<���`f��[��E�l�^�����d��H1�Q��aN��-F�X�hoE:�\�Zw��wc���6���'��ϧsm碃<��'�o�GM>J�>�#c�;�����c��DRH��/~����T.���%���M�v@�R�.O�Ӓ�`��cn����'M�S��ͧxm?f�F���/
�*�=�-ڂ��z�@ϩ$x�O������k��0_��z�����x8Ŝ���z;��R��� ��/;�@s��F^d�2;��:=���ykn�@.F�r �Sٚ����,mx�C7o���әtz�t9dc�%�3&�����)u��|����.�@����ka�#���^��s+�B�mc}�54�.��/7�r*�9܎�Y@��<	J����[7��pt���Euk�=6�:�%���������R��8OC#FP|���vqc�y�?!O�ڪ�@mԭm;#��*�E`��oOW����Rd\�./;�y>���zE��)�{<	�X�"-��n�"M��5�#�@��R5ᠩ�	�[X�&�3�Q�����H��"�Ӓ�I�j���M��~���%d� ����Y�(������ ��>��;Y@��lY���C���g�s{���Ar��H��c���Q�l4r
� �D$��}�]K�yʺI���m|��o��g�����S�������߁R�.��{�rP�]������~�y�������4�ב ��ڊ�l�4َQ�i��P�q�Mx��T��QJ�淇�zƱ��yV�
*W��'�Ķ�p�xy�mf�So��x[�l��������ކP�6�!�-�þ�P�AIP�� ���~�����!#M�џ�T�d�T�T��|�뎫��8%ů<��/��%�F̪�[��f����禔M�X�>�z5j����׍�v?[�����p��}Mp�U��F	��,S����m�Ej;�-G��n����������pD#����o�� |t��]X�D2޴]ІK�����O�4G΅�S���~�H�����+S�føĠ���:�緅d:�$�|�8���H���p"����3ox���%�<�s���Rc�ܞ�Q֯�boq�*�Og@��UM�F��i� ܪ��[��xe���	oW�W��s��x�EF�P���f�	�G�q� ���a�{��&�kc������=���XF��B�>�i�e��?�$?5�S���ތP՞���v��]dN�_l'�^p��c�=Z��\�+�;�6�'A b[Ĵ�,%��3e��+��&����)��؅Y� l���i�>�*#t�@>`�,�ʏs��s����֖�ɍ7^��١��z�F��~ϧ�M1G�!xY����G�D��RrZ0�p؝��KO�ޟ��h�
�.�*��@,ö1��Դs6;tW<@&,W��deeϑ�O�<���B���3\+���Ԟȁ���PQ�$ơ\�
1����"������������[�w� ��_��m6�:W~pW����� >���$�Q���$÷��ͳ���?�`�b�l�ܥ��3�Nnr�-�pt�옐����>��=
���J(�`�"ں�ܶ��v�^�_d*>����)H)���\�||�>?| ��%W��~t*����B�s��N�.��[$�Nﶟ��F{��B=�60�Q����[h�`n�AR=����@KN��	�o�5	���i�PF����S73���G	h����w�{?�zw�$;��������|^6��~g��O��b�o��NP3.$�>U~�i�ݵ@C_���j�
�,��7��y�pр�6���=�����s.4�N�_�]��2ͷF�I7�x��� ���2�M�vK��L$���u�Y��:`7l2��tMw�@�I��\2��}�+S~��N
���ag��y��r�*���tSs�����| �Z��լ��
$�8Ri����n�Cz�6�]�	��/Qg�+gH�mED ���!�5��Ԛ�LĤ5��
q���EJ���%^��	���m !��#����R.!{t�����5�[����j�@Y��K=c0^v�b_@^�_rmOY2�^��8M���g+kT�r���Dt4s$�6d��ں�T���:g��Rca�t7"��yxxL'_�(;���d>t�؞�!3�$�N����Ǟ�x>;�U��o�u`� ���)�L��ǜ>��D�u�W,X�SK7�Q��^6Z���q�j7�9=�)���� N��kϭ�ў2�@�qժ�I)�PSξd4�<���q<����������F?J��p6�PeM��v.3�D����Et�L�;�D-y��9���wd�)���@�+؟�T�{�|�u���[|+j`�oX�Qc��M�Ҙ!p�=����*ǻ	vN����1��?���G��n�neZ� a=�s�â��ׯ�Q."����&j�խ�VNʒq�t����r{���G���O��BE �[���4��k��T�j���௘O��
�;i�'�g�w)ֶ��k"�z+�}}�v�Tk��=������v(����� ���p���*z��z���K� RaB'�5�N��]�\�yr���S�?��$y&�4��v߂�d�Tn���S	�����c��7p�����7�ꅅ1����C��{xߤY-(S���d���O#��J,I���צ���|mƙ���$�Drܙ��������'r�b���t1s�k}�'���F�񌇋�68��
�������.�J7�xQ8����ܳ�F��1Vy�H�߯;z���w8h�Q&9M6�<�]�F����k,�-\��@�A����fk9� z_u"��a�wW��JH��)7Ag���V?I({�������{c]{�n 4�*�l5zZD������%A����Ĭ����Ҏx[@���$� ~I6_���V���d�������߼�ww�$�}:K��4-Ѐ�{s^K����L5��6gv��\(w||X$�}� � �z�OD��GN�я���j����{�#傋}C$T#
��\��aY���g�d�ͥ�)�1����NOt���4���lڻx��vi1�=��HEx������IԖ��؈��cf�70�Q<\hO9�ٻ�c�+�̳��6��N�Ɩ]��<���f!�1�"��/�aPcDo� �j.����e���D�\U���JD����E�\`yH9�L��KA?�NO��C˳��=�u7����ڻa�'��a���m�vª -_���C�\��p�l��}=��g���f���4K�����X2;&�Ű>��6�;�ձ��r�-���{�dP��v�b��SN����ꗟ���Y~�<��9"�0�\���>\���w��;[����S(��fw�r��Y<�,�PUJ~� dS��5�1��G��~|愞��>���o�io`8E�L��;�'�k~�w�=���D(q��K�6?B�׿�Zn��L֦����H�v�U���~���!��;��MB�����L�Н����_����IX�e��e�EuSk�W5�X�s$zt�J�Cl͊���4�e1�?�*���:�+����,�P�a��Y�؀���F���oT<�[�ne_s\���/�,��K�җ����Ir�i�}���^�����O �i�.(Oz�1!�g��>;�o�(-d�l�c����#�A�Q#�����ZO�*�	A�$R��]��l=��&)Ӄ?�4��2/}J���{� ����a��ۼ����i�%D��@�,�t��V#�(a����F�%Եf�)�l
�ߺ��@%{";���N  ��h����(\�
� X�]�ͯ��a�陰��&�!�2�D��x�k�9�5x�^<p�_�]c}f�<�P?�t��a�M���W���o�9�t>�-s��\ S�sw�~YD�	�g�B����)Zm�b�@�2&�X���)�i��w�P���<7�G��̚�۹����7S�k�ͯI
�@d�B���9V�Ց��q�e���2%1VY���c�M��1ͷǚ�7�v�c�+Y(�27�/�����!tA��o��l��짲����'�ާS�lz���X�g�(�=Q�;Q$%�w�e=�i��C��
3�jF�~��0VZm��.�)����ذ�5�ʮ$��,��V��0��JeX�"�u�!-�cV��M��:�����CgV,��ge>�<��i��ߠ=�BG���&��ty��f�xG����̐����I,X��㪛j������H��'��ǥ�>n (�0c(��f���9r�����7Dܖ]�$<-T�q�.D�rT
��opE�l)�(p���m���OW�޹��5��u�<��b��, �����G'ʏ����	:(��<�#�؅�<�	�:�?z�m�>�H���-{�E���e��t�ڟj6Dt�O�\<%�:�������{��������k˳��c�X�vln[`u�6&�Fb�HAI��Xl�ae��s�;����^�h��o������g
o��x��f���АJ�{�%�_����� �?�`ػ�$�[RI`k2֦M���`���gxO��
Z�ez迋����
)-��c���V� �_�g��rœt����hrU��3�pM��徘�~~�U!2*�Aj���H�7>|Si�|Ǹgc�0HI���!�}���OT���Ӳ�t��k:�t*��S�U��ƫr_į_ˮnr������F����n�r��Y�}/|�υtGM(]�?�[���R��SO<j(%b#,�@t!xR�-���Y��'!�7�	�����e���,'��A>yش���6Gb�&)�����{��7wí��[�-�tm����'��j��mU)��e�U�1߸.�"� K��C�z�[����s�'�l��;���}3�)�v�"��,:���Y-j��7@��k�����z�!| իL�KE����,�;�\ɵ@fD� t���VhS��=��i?}}r���:����Dc���%�'�Ye�s%)|K˵�y�iِ��	)'y`��V(Ab����
�"In6vp��,��eRe)�-�I}��'aJ�߿����?�!Ȳ��mS�'�'����~��ڕ"��)�u���yI��q�*fa#wC;e��w�V^NW�.�ɩ
Q;���
k��I'�W��
W���7��D�1��H�Ԍ-^�^l*�>d�*���{JU�@��ڒ����@0%$�İݣ7���ӭf6�����ί逪pt���8��:�-���՟��,�Kܳ�o�sJ{���x��5��GL��h�W*mF)�P r'>G�<�<b�3���v�(�5Ta8��;D�@��6�u�/$�Ig����|��e8�qh�i��Z�M�R4�ip� u�tak�;��Z�i��a�UwFk�&X�b7���I"�Eg�Dq��?}���C�a$�CfeS���v�ҽ��R��w4���������ml�Z�����[�A}�cɝG0����X���_)d������&�(��/�&I���u���<���^ڢ�{7���ZsA�l�]0%���h�8�s�P��X'�m�^�-����Wў�Ȇ͹�B-��A��1;6g��@��%l�d�׀z�@��fX�x��vl�K���,O"r'j�H�����<�~5��pl��S +ſ����w�V���4[ �fe�Ti�}tC1D9���)G������;�e��E�����l�{���L��Ћ��|��50��X�u��]I��K���b�\���_��
�7z��n��;�j,R�����<&C_OA[�I<��A��"MnC��0_�⤻�و�ޮAZ=��$%�N����19���ؓ	�ՋwW1�����UH�V�I��m��r\X_uI(��?����+)��*�d�壙�$!.zNذ����N=�ǫh�V��ϷR�������k@���!�jG��K* ���u�߾�$AX��K����f��ϔq�B/�p�ёE������WdK������	^`-8:���xl��K����*��ɔ'8�:!�������7�!_�v���v�'=���F���<w-;F�p.Et����[�����L-�%�''���7Ypv/�'VU6&���wR�!�)M�7��Y/��r��Z�V�\�_�~��?��q�?���(s�sn`|�$��6U�JX�z�H"7e�_�б��5�e��Ӛ�D��;	����]s���G���!�a�P�������f߂%�j|6�j�^p��%��R5�S�b����h9�j}����Ȑ����p��(g�Ō���̼�ю�g���E�ƶ���<�&͆���һq`4q�Mf��,yBt�a��+m�ڶ@�cў�i�iX�h�$�v�3G?���<A����e���'�Z�Z����F�ō��g��`f�s?
��]�� |�6��x�]��a�ҟ�����}���z����I=ˬ �չa��Y��D��*t'L�?>�棎���=I���	N_\~ݘ����v4�eSoHqDZ���y�z���PDU���5t{��>H�\*1����z�	�*"_�����L�!�����>��~��eô�pȦn\�֎)������,5�R����}�>��kI��kt�BV�ɫ9���1�;���@gvh@\�=��(��~��I���rOOʿ�����կ���߿��]�6����C��mY����������5�d&�X1ӄ�'����⥵����ݏϤ�[HNu��ѫu�!�����M�*���"�Fv&��������8><�/5�-l�[�m�x��c���!�g=0  (�*<��X�0`�(%�����(��r��w�xq����|�v�<o�J{�;�A:�/�ܧX�����Tf�1�����U-�� ɛ'ɋ4ck��q���������,�L���Uz�u�PVN�k�<���/+:D��ߦc�Ñ��Z��lO�4�`w++(�rzY@@ to��
Ao�<��%����>
إi�3WK�'�O`���I'���5�a�n��̥�I���7�ă���ݝM���i��+����SЩ�9��ϰS1֥�_����3Ks�*,��e��h�Kk�6'88�� �e�`���NVz�=f��������G����<���?u5�	���,,T�;�N���{U�R67�����6��A )�E��ޘ?�J$E�nZ?)C�e��8�&3�U��E
/��Kr��K��S�U�Kz3�Gi��o������&�/E8<=�b��:8O崹q�UW��`�o���}q�'ؙ+3�����M���ރ��߸ͭ��S�S���~��u.��.�R��k��H�)�륚��G��T��lݘn��[��<��l��+�*��3���=ϸ���g�O�GVH�6�9���C���`���?�p��x�rJh�|���S�h�aW~��.X�)4!���7���1�=�7��c�mG+xe�lڍ��伴gnE�K)�[��rV+�#x���T�\��'m��ڜ<ɕ���ѱ��X��Pӭ��Ŕ{9��H-+����5�m�ޖ��/}�Qqϒ9ޚU_���t̃WOZ���$C�g�_����ض�)�X+��(~� ʃ���)P�?r�$��_�$�|b}�-�Q� �nҀ��`[�nҚ5Β*�`sz6��`{w��{�e�|�(� 2Ra�V�^~0�3�xkM"|���g�,jH�`K�#��g�,�%�=���#���_�&>�A��O��RS&�N�1]�h�6]�zٱ��v�{��D�f1��ef���ᚚ��܂f�F8�>�6���cp ^p*��0jedݖɋ�y=~*��:E��'!#R��}�YҾK}�x}9W��,��'�S�q,�������wwvpڪj��.��~~�M+���*�V��J�����X����1�_�Jg��#�P�S�D"NPWBϸ{��&I9'}N�Z�_��DN�����=۹75�E��X�E	�ã��o��M��/	w+���Oz8��X��'nw_�,?T4����@ҳ��%^`��@���-������V�����#eecf}���l�9��t��T����x��	�Ϥty��$77��F�[����Ҷ�2����[�⇗:�~o6N���$.]ힱ�t��&� ��v�񙛝��M�!9���AU��Wh(�~U:`�)w?���A����K(�"����F�+�	;�9ztfV�k� ���֚9"}�	=NRH�����V'�C'���)�����r!��{\�d�t]��g�|Ɖ�,���sU��j|������M�)N�\S�hXKW$���C�(ljk=��u�I7vxl��@���qi�<��%�������2U"
���03�A*��'�r)y��n�yV$g�0��gF�&��)*vmo�4�(N�����D4�i6F�=��|)�ȷ=�̄��]nأ��T��y4�o������o��g������56LY��z�3��'��\>p�"e���������yR����u�H�ǲ�P�1�����`�Y���o�|X��I.�,�5��O����/s��P\0�F(��D��^dqdw�,&D�z�`��C��� �h���q��~m��hO�BS��C���]g����,�45$���jғ&/E��s<}^M|	^�l�RZ�5ڭ�;Bw�$��	�޿�(�X���iNi��,�D��TN�!��8�#p�]�Ǫ�'�J�.t�&��]� 4:ofB<@���rȪ�����ϖ���6��A�Ӭ��0��Y�#q#���K�����x�s���w��~cc���@�+ �N[�vͦ���.u�9�ۘ{Hm��xH���(��v!�I<��!�"ծyRS��
2Ƚ���.@+�䂍@�d_d�P��t��
�M��-���Hq��Sخ�5f��@�Z<ՏWK�+G:k�ع���f�^�%va�J���$��9�Wᣱc��J��
a�p�)��/H�M�΢��|���X�X R�����՞ڗ6���Z`�G`�%���� 﫥D�OF�þ��k�}C�Pg휳}���w�<��� �RϾB~���J�pF�lM�z��w�^���9y7�u�D~g�J$S�EH&;�z�K}�6p�k&UD��Kb[c,t�/�~6�
��3�_�w���<">��0�[}���x���N�E��b/�����$ih��O��>���ϖ�����u�ik�%��߬nm�8�������p��NL�݈ryY��p�	�`-��{��HQ�C���y@Cx@n<���<�	ߗ|�@:/�D>�M+��C7����#����qH��A�3���z�>�����SV�����_��M�|�gr�Y8�iD�f<��p���@�D��ט�\e������썴]UX��|d�-D�p%b"X����k��D�������Rɪ���t�N}�����u�������V�x��u�n]5�|Yp�VF�8�܏'L��F������i�<>>�}-3���<��&��歧kN�Jwױ�2f�GSC�xJ��� �K�
���|M�lT>r���]�>�S�ߊO�J����w\A2c"�`��	�R3R}���f���`��UY���+��("N�W)��?_�*��
VK��֤
�5��[��\R;u��%=�q����ɹ2]Պ�q�F?Deܻ���מ.��ollB���w��G-^>Eʰ�8����H��t��{s$^������v�*���r��F��o�E�6��b;���$sڷ�sD��cߟ�bV�	��~_[�?��;'���ˑ�?��#ۥH��i}�[�`!���g�B	;r�TsF����`/'dff�~�IN�o�C9�ݱ�l��[-W0�WhO9ŕ)��_%�zqmm��t�y�n�R+x���#-8��u�N�V���D>qS8U�˒0�2�ɥѵ��4�/��[�l���NIc��$d�V������im!UUݕ�N��m��7��^H�]8����[U&�k�`�3���I�Pơ�0-���L2�nVœ�b��Α�O#�
(�nƶ*7m�#�O .���8݅�(��ڎ�VJ���U	����`kF�؃;oi bV�ɘ��{��+p�z_���"f��fi��h��\����yQq:�/uU���p���.Q�D���LW��J����,��_��U��E|$*��
���&��v�� l_��݄�FI	���v	��m�gW�8�� 5�q)�B�����bDMG�S���e`��t���ڍA�|3���������G�y�|��\.w��*ɮ~N��w���R}��}��A�W���\^������@��*�η �a8�������m(�\�;�d�nǑ�vaF�R�n�O�Z����h�M&d7C����ɓ��~aa�YY�i��p:.�3�S�D
q���6P��s�K��S���_�E+�Z����`e�/�/����!�yQ5��5�T\�A�撩4*��>%zIY�SUJO�����������%%%�R��t����T�M����"s��O>G�������."�t#]���HJ����K����(JJ	K/�t
H��.%)�t/���������Ν��<�ܹ���m��+ݜ�U*��ӤU�4��>/!d7���,s=������N=����D��s���%C��͏��P�CS��F��$!pw��N芧r���[+��������Y�v����D��[9����\�A�dmmWe����>����|��s��y�'��<�tg�y���N]��;ő'A��#��њ	�� �N�w�(%���(���TJ^S�����m��$ţ�ǔ��U#i���+�<{cs��r� żK� ��@�C����#V��E��i�F_�|���h�vF�}f�m/��L�~���%����<_��ff��g��9oծ������(� ���2���D`�CP	UR�)����kǴ���f�<� .�K���(3$nB#4 ��?9Ҕ �Y�<3^X_YK͓>�"A
��9x��M+ �%'�Ɉ��=k���ѐ��8G�6��q���m(Y�o
�a�� ����62:�M��xՆ�t{hӝ<"~�g�m��%��fXy
q�X�����lz��O�?��!�x)7h+�u*c:6�����SuU�'�#���;R�o���A�G� ��?t��H��6H9��ʳ�Wҭna����<�?��7J(.�կ�o���J :5~��?�Imy�˹q���.*!�Q$�������U�"la�;����a�u����͆RI����}5933��'��X����zza�W��-#M~���60d����2a�ZfO��5��W�?eWQ�dP��~�Ϩ���;9 I���QOn�H�G���w��z3�=���)������u2���'hUm���v;�-ak�����ηtg��aDћ��Br���k)��̵Y+Ƽ��,f���<u�$�'�,g� ��_t�اII#�]�xj���]��ah�t��A�%W�I�,�4 e�rU�Ҳr҅�V{O (Y8x��YrETP�3��2���q-�,|���W�`}ǧOҽܸ^
��D�ԩ�O��)&2�D|�p���?m�����⽹P��ĽO�=�8jc�?�
}��ocE:ٹ���G�ăc��ui;�ރ�#�k���Ԩ>�Շ��d��&�#�v�ф���|S{3�0��_�i����qEk���8�7=�$�ɕ� ��~�lb��q���$���ؘ�bE�B�Gd$2A��t�vw��*B�æWUQ;=��QaeWi�r��f��*�-P�C�v ��ƾ���6+y�=�b�hSr�-��T_q�_��squ����Q/d���A���K:ܮ Gr�N�7���X���]�{����6v�� ���v:���0��+S7�J��1�ʻ>Z��FrK�*z�|��8����_'ߗ5�w�"kt�aMlC��O��d��mxi>L��&B��Њ��?Z��C��=�� v�߻ᡷ-�~y�f�X�:k.^Iى���sI�G]�n���XG)�Zz��'���;NN�aE�'���}@x�D����"9(��(qp� D����4E�|K���bW������|�0.k.�Y~��^B�H��~�<�¨|�(H���ɣ��7�/��Ytէ*s̟�O��xƺ��+=�`33�A�י��|��6w��!�H��d}X%bz�]ߠ)9+aO�&]�
Ĉ��+�%^�����r��gB��&S
?l���S<~���[�^�?�@�d�|TPƜ�����4| ��*�!�s좭&D�U�����e	f�w
ǥ΍h.��4ުCުH�}%�妡R'���^z���.��	�_�I����D�z#���r�E7�W���{�)�\ �����3��R#9Vq���d`��B��|@�d�����AP߿�v?���IU�7Ӣ�h+��������3�Sv�F(w��y�f
��eh�kF�;��{��J�,_ҹ����%� ��&hfN)9������2E紧�*�ԃ��KJ����������HK���E9���O+�:i�wF	,M��$@P�f u�L��Z
;s����7�(�d�Y��y��a+�4�b����_��	P�a��~maى���Uf�=RaQK����U;GY�d����w��uH@ǉ�v�]��CY�T��-��4|�K�x��^1���۵�=�����WM�$��.M'(��I�U�����yyv�@��=�<M/�aPnq}�3�����Ig�}��ϟ�6���ĵ��{����;��J�����	��q,Z���+
3���h��i�ӺP�=��gl�*i��8x8Ƕ �����z&����H���Ŷ��b��TBDz��a�L����Ǚ
���k��x>�\�z.<������F[�,��Ǝ������b�YCw�V���c�������t��jE:�L�y�\U�?*r
x$Ɵz:%1c��:g?��>����=-�'���$tD��E��I�GO�$<��� �����p�2�"�Pܶ�X����p��/��m�_�����{�a2����Ј��?i��,�P���]�^`���ͫkj��-l%YDBL�k�YN����O���Ɏ����:dV�1��'C�#嘉M*�:�xc�Fۘ���04�2�"�M�iRۗ��'�]��|\ҟ�di�7�Ѹ��jt)�O���̢K�A��5�0��qҰ�Sp~k���/�<q���?���"bg���u�P�yWq��s!������o=&;�]`��J UB���^�O 6����Ğ���Eu����}����U��|������L+MM�i������ע�F��̃�[g���ʗ=�ҘWnKz@����s�RvK崽�'=�h�h7�~��������������qE`V���+�O!AS����A��q�".�����_r��<=�c0drSS��\T�F}'�-4�2�n�;�S�$��N7__Q�l�{����>���˦��*��]H����|�z��L�~Dr��X��̚8PB#�ý�s�A���0�|��+D� �L�3A�5���g��5�}aa�k� ����,/N���NY��J��+)V��6�!�;^��7�L�pXe��E�ǲtX��q�t|o�~�jH�V��"S���M�#R�C������v�V_����!�5���i"�$�瑀ω�1~�l��U�~�qC����B��x?%��٤	4�z����+׻/V�W.�S����g��{k�@J��ʠdg���ɐ��J;��pq�����|���m�т>@zk��e.ψrB˳ ��^V��	��� w�5yrR^(���	�����.���q,��������zl�̽�TE*47�|q��N|Ez��y����m)��e�k�X����R�>�91
�i[���ߜHqw0,�֧�|:����ߟ�<���B]���7�jb��S�I��-���R�8�k%O�;�6�=*�$y,IIh�4
� 8�*��K��r:3��(y��(�LF�F�����S����f�`�_�f�6�]���0�(��0(�??���a6�28��b}1��"��c�X�"�Ƣ9�x����V����n1]f��ͅ�Q1���7U��9�?�f]I��!^�E��^���D��e �����\�2^���	�	~@T��.�4��v�3I0Q�7�ka����0n�����9y��������q�ύr�B���+�Y仓�(F>+����zXbzdjj�	��L�*	����!X�G�/# w�K嗦H�����=@������:׿�V��l3T�e&��8J��:M����]}�I�Q�ۚ.Rbv�P�"_a��[z�lk	�i��|�$�%�R�{����[���Ӌ0�N�v�0�Q+�U#��l�*66v�ތ�V��fo��o'�]@���W9�K�R�����T��hN����>͡���U�w:��2�S���2�� =���Gl����R8�Ks�9����a��EQ��'�z��nP�7���]����+���e��~J����~��	+��@X*���b��̌j�#P��[��)rξY��L�˒py{�C����U�i)����5LZ�ꬋ��`^����M�=C�����ќS����2�/p�,�]�8��s>���i�k �2c�@R�oR��#s�����U�E�S�{�o�]�1c���
H�_��+�<��/�v�N#A��a�	��'���Rv��1�A��'�޺���]N�ԙ��U�t]|��� �NL�Tץ����������{�LE�j~��`F��7WL�	:Ó�X$����"[ת�k%)4�P���P9T���@��a4��OV��vi�Lu|;����t �?��պ��*c�d����~��܈���i= ����0A8�{�+ŻK���baqr0SA	�E�>O�?�:����%���o��_��) ��97U�D�T��!�������S.����W!�,,AA-���a��ʡ���-�s�����L�y�~	����5jS
��N�od��kMh�</�I��*Kj�Fk(�=�׫_2s~�|$�'��!�euZ����D@�=���;�� ?v���~Dnf���i9cy[ Y��239r�f�zv/��[�1��݁_�E��e��8
�
��K�7� �ER%q�"��}���Jo�nE�*�n����P���o$[�/�s�붖Fz��5�҂���r%kٔ���^U���h��v�$���{�/8��yl����KD��E&x�0c�بa���T64��W�P����8�L���A�ǫ����O!c6�O8 =���KO�Q�~��VwT��kw�;�m��	�N0c�z�Q>3E�p=@�u�#�f�}[ΰ������I�N���c@�)i%9��rty^�4��K@���V)��cwW��~��+ϻ��~�кO`��i����c�Ba5�O�"�����z绋��N���6B����jT�fNg8�W��[�k�A�W�߃C��8��"���c�l��F7{�X��I(�3�x����]Z���Y�Ã;L��2�@P
�5;�HM<�����x7�;y�9�c)��j�
�X?WQ86t.��\�~�~ �e Iw�P/zIpx�w�D������2������ȼZ3�#�+Dj�-���Q�D���ŭ�`_8�ց�%w_��'�>�`I���""Z��YP�e��췾'�=�ߣ�{�����07�yF�K�9������	E�Ng�Ӻ���^R���B�tk����7���Ӗ?5�7b<6�!���)Х��fu-gV���!�3�1�}�D9��PX�V'C&4@�O�V�D=
�r���a�S�a�X�V�$�ٜ��|�Za&�MJ��잼�~�?��M�\�~V��''i6�ٍ֭��Z�4���D����I�
�K�S0�S�S�%��Yxy�V�"+5�����&�I׻��쾂LjOAb})�y��q��>��C�Ahs_ޤR���}'�u��t�n�����@�7~$_��G��NF%��;�T}3_AW=�6��OW�L����z����R��}[����P��G}��'�޳W�y\s:��I�IO;7��4}'��᳾�7|�W؆�VR�e{1��Jw&�9W@#C���H��G� ����tjJ����c�֔��Ov�p���fn����T�=9����Z��R�`\/��y\�wH}�j?���U�N��%�@�y)���C6����w�T�\#+J�m�ɽ�K
4�������
�N��~�b'�ؿ3��M:� k=�Fퟔ2�[��J8�U`��k��o[]����Qv�z��vmhh��z��_�)Qh�: �����!IlL����߇�o��J��_1L8
��J��ޫL�̣�p�bX�s|a��Tq��AՎ���{��l,���ߧ��zi�W��''�PC���C����
ܭ��x!���o��s׳���?H�7{p;KCތ�RU�iKL�N�yw&!3h�d��%^MC� �?{#�֣L�y��t\����I�ҵ4�>�pQH���H���9�|�N� u�V#��Z�R~pdW�l���E'���������?�����F�=���hV-��I�X{�Ի�67��D�b�cV�\3&�+��~����>�ݙm-��q�]����a�I��x�576R����]~�/����CH��x2�~3 �	
��rv�e��|#U~���,��H��r|�>�@�#������++*,n�TG1��n�77�������
�ٖP\\�u��HK�,����Z'346�K��{P�T�C�N��;/.���3��Z׊���s�-�M�훭��r� �!�rd�0�ef��I\��]pӒ�b �n��#ŒGY���fN3S䍶�|��\�[{���c����
�~=O�������+N>��\,xdu��Z�Q�R��4���~��� �O9H6�+��?['i�3��Q"&Ǥ���z3H�cI	/�����3,�B�E��FH���tI�޶d���,A3S��.�T�/�e���x���UQ�ˉ�ç����ퟥ�9�~O�� �PYWgW������G���K�����o�������nN��}�1���Yh0�z�5�r^"x�9xy)�U:��S�uo!��S���C 姫'N�6N����Y��@uuV:�uR~(������X�����H&Y�_U�����o��"I�S��u�������4>�U�4ޔOv�N����9��1��[__oPs�tJ����m�t5(8�X$�g��9&>9'��K�!d^/��2��05��xX.���s9[������9��z����W�K��qo��c?��=���N8�������`�\ӁM�����rv���]���U�{ɪ���eѩ�0�A���E݌ȣ3�!�s��5o�W��-�P�^�1ˆW��� �wSk��h �h33���,my)�jSUE�cnBf�%aJϺX�����?>[�-6��y�j��q�$%5u���up��"��
d2��u*��1\�,��I��v�X���4�N���J��L��,L\:���t�O��m��-�_����,	;���R��F�u����kà(���iW��v���]����5܂Q�{;54�8\O��fw� \�U���듛��K���e�����_�������egd���p��*���,��I~_��y���ȸx�B�_`���}|0�0�l�F���<t� _�� ߢ��ak���!��n��u���S�g����LO��]W<ovM�H���W���x)gn�U]]m��Է��i�e�\�>�A��F��O��=�h�?Z-8|�}Ju����Vl.���V�C����.w1���5�>�;LF~�)i�_F�sٛ�3=}�r_:Y�Ԇ���who�>0���\Lpq��y��q��{�b	6�7� ]9���q���	*�~���+!�ĻS�j�Rm��ǘ�"��Y�D��r_�+P��X޸�?0_avј 4�0��������wB�>�݋���ܤ�̵����R�w%�픈�봪pH�;P"J����k~�Yq�M�f�h���"�i�JM�V�e$Hօ5Id��#@�]Igu�)@�n$:Z����㐬0ˁ��Q]�̂����U~��-َ�$J떿.VVO��7�1<j0��~�����-��Vr6�!�a�S��i/�~�5c�4f�/al,���"��⽼�	���j:�j�kT3���M�Mr*��<؊}f1��<$�U�~���jໍ��+s��8b��aW�E�V�6�6��u�R�=?2�x��M����C
�Emu�ѧ_���=%��3.ӯl�Y�l��B��4�ÄOH�Ŭ�u��[Qxs�*�XF�����I,<������,7ifO��T1�=N��F\�s�Ie��-,�����^�qz�	��䋪oP`��OSÑ�3�F�����&�dP��](KF�(���m�cg`ȹd8�v|�`:�7������q���^n�D���@rK!��>�8Y�ڥ8���7��q6r���Z��w9�������z~D"�h^ب�uʎ��ˍ�F}�_T���%3W5��>�q�Lv��
��7� �����ͺ�(��،���#QO)�!_��Fo��/ˮpN���z�Y�F��9d�_�����ir5�"�L*�}�!����bɨq�*WV�s���?0�]�N>2� s
�2�S�6�mM]��ߚ�:3s�'��	lD��S&v����Zf�P=���1�ۡ0�+u�ό�����r�;�˙t�ΣA�3#^Ϗ��OF����
����~
�N���I��D���`�?��	&p�H~	���}A���q�[�b��:y�.U�6���'
x���ׅ�~,��2+�h�@����XV�
�����y�% (}wqʁ����,IU�QH&��UDЯ��웤��Mp����(��X���o��(]]wث����⫊��(�R���G��>��a���i
��b�����o��2�Scs3��%>���<FBL�$�}�<6�ۛ)�����_+�$��h�JL�+mD5���w?Cw�lW.�F4mL}Q�?�~�8�>E9�G��6���(	9?cH|>��M�v�@�MAِSKuI��މ���c� A�T6��	���<weSv�/���Փ'�� �^��4��mZ��5#-�h�tP�-��o�ow`����ԄW�ⷢ߮z�W[��tX��$����vǫV��MLlz���n�F���V���R������Jl���h�d���[v�/u��o�i�]zV��K�@�̄	H�~�NX#cEA�ew~ff��kYk_`q��R�/�|�-<,��/P�EAi�Sp/�7uE�50�T9��M/�M5j!��R����bfH�Qc��pH��i(7e�!�� &S��˨hu��:B�qH[�0M�BYO��R��m�ST1�ԯ��HI�޸�ΐ+A'��O��	J\)�����`:���a�H�Ϋ���{�v���1'����s��a�8/nK,�{=/@��`�4f!����c��M�Y�"D�n�<vs�?8�?Ľ��� X�DM3�مE�39ʒA�_�vM���AU)_j�OX� nIE?�*'���������)ۈ�����y�ۍ��Fl��0-)z�cM��?�L����6q~A	K���W$'�A��T�լ;a6�N�s�[tV����xL���4��E�!��Sl<1��gݨ3��k���а��03z�q�D�̅��7��ք8}0�&:\�Y�eF,S:~������x&QrV7�.��zq�����ܬ(�eA>�"��#͐>�T#�i�HB5u#4�,�n�V�u�6�:�����/p���z�t!4#rG_����!�ɂ�~��z-�u��"� ~�a���r�/�Y�؀p�WElU:K��NھbR R�C,M���6`���<ڝ���j4D9�xjM���y��t�8�+!�l�m��5?�[�|�K��:�}����vzJ�����"fØ�F
��ϽI~ҳ)���y��b���3��0{�Y�WލT%�^�~%���m�����3{��H?�½� M�uN�!<Is�#7��JE! �(1�#奓@|�UݏN���k�'!�]�c�_��DQ<��<S[�|���d��Ӆz�j��J�C��$3Q��r�=���}�w_�EQ�}Ѡa��#��ݯ%//I0{�oH�����q
�v�:�?�t�"`����
௼��F�c9O���/���܃v0�h��x� ���j�]y34 �ϥ�α{	\V���SH�;!>#�,�N�|f�`Ԇ���8���^Պ��/�Y h�v��j+_T@��W)�
GuاoiL�?VCRA����G8x5�ix���M5��l���sNz���
~����>WN�-s.*f\vK���Ɠ�u���%%���b`+�o�- ��]HS�`d~��W����T���D��)el�h�gz��׽癛�?4�M:z{f����4�F���	}}�'�06��v�|��ڍ���z�N���F��^��*�a�mt&�S<�V 12��<�S�/�
}`��AF�8�35=@��b��P�H���
��O�dh"9A� ��hz���^�pE�#=P7I�٭�Yn9g��E	M�7�D���?��4��V-\�}�dH���_�=�
��l/A��|1�/����Î�i&P'�/�t�^��]:fw��^~�b:;���k����9�k�/�� �����^0tZ^����� "�#��i{�[��;���]J6J��O�(E�E���L�͏��Z5}���R�
Oo����l��p���i[y���I�c`�;��Q=$ƥN����ԛBPqbCK温�ow�H=@�zn�ޮ֨#�hs��@jx&IB&=�3�a�����}�X�*��ԭ�QRRo��C�t0���~�l%D���!9f�9�Z�3��a��w��2�nÈs?��)sw�:;-�Ћʉ�����y��v-��O����^����Qra��hhX��׳)���=r2��3V9�~��Ǟk�& �u!N���פ����I�MB��Lx�Wg����Y^��m�z|=G����n���(*��x����M 5��k��� _N�
���u���A��!PX��q� [���b�'٣��a��T9s��׍��9no:H��c'Γ�RFْ�l�����}���Ix��,������%a��ӯ�E;�hZ"���r��8ā`�I�tjv�����mI��
㲷>9�^V�]��SoY�.b.��Yj���l��>p0�>󇉀�)2���(��ӻ���^k�鱃Mj���d��� ���2���?�Ӷ�����Vr�{�C���;q�����g�9�;�_#�g�+KR�[�W�?�Y�����6"�$�Bd�Z�*�Ӭ~��@mo
��؄�֊��X���b���_����Y`B<�ă��FW�j����ꄸ1�)��̸kޱ��V��������h�}b�i,�5<O`�t{���ʐ당|�ԉ���)�i�\Y�Y�����]y����{���(�&�S��9���va��ڝ��x��	KKr���2�=�K�>�v���2T'��� 4G���T?�F��)�zq�M���VE��$�e�
F�_e�rUmi>��~o�pѩ2�$���A-�qߔ]Y)`a�/��L��'>��K�E��Ta�O��P��E!�2��'"y!@���L_��'���y(���'}����;9����؟�/;=���͵�e������8�B�`t�R
�wM�Z?[�U�v��W(�����F�W����@i��!��ay�[�����0=W��q�e\J���d�ȸ�a���WAo�q���G{g��R\c[�M^�>��@o�<�I<1^�`�ɺE:��n�����H�+��cE��֌w�ý��-Wq����V���{%3o�_�P+ao�����ݴQ1?r5$vss}~6�I������bo�z�G����q���_șJWJ�3����ย�GDj��BmS���+@�Q9l�KQ/"ԍ�.�ՙU8���b�5D� ^�"��w�1,���[{5��?VkC�n�Ţ�#��O���7������F�C���}U�҂�E1QM̽ny���C�l���O���%]�8�|��JW�ٹp��E�7������=���.^���my��=N��UQ�B�lTߖ��KcR�Xw�p1ԣ�A��.Ja����pzo#��i�&K��`d ���媟l�gGϭz`F��-�vwZ��b�_�'��k���5��'�fsw�2
�`-�w@��e�ט�$� ��͇��ݷ*J�Q4��l/܀�5ݛ�U�>�����z���t�������(��?�u�;"e	��qj���7(vS)�.��ʶ��:u�9�A%5S�P�bQo���ׁ������D`I�EupK�6���2���4�Jg[�l���*�Q�$������Z�ZiB*�r�91�iq7b�u0<�<�f2u�"uڱ�G;c0J�)hv�MGǙ�x(u�k�o�"mo�b{���n�!��L�gV�]��{A����(�~��p�K�}����S'�*B��4l���>G��.Ԇ�˷�k�E�t���m?m���E5?�S�e��S�[��_]	}y}�e_�jPgG�;����ț9�e]�N�3�'XI��@��Z��(U��Z37���SP6�DJ�8�\V��"=�$!D�CNL0.k��cO��툐?X�ϬCsJ�a���/#�E��݄l�l��vq��򉱘-zl;�LŪM�M�6׻��J�ڂ#��7��>�	V�p��-u��.�J O;p��k����ٛfx-�2o`s���n ^��ڹZ�ǯӀ�^eҕc��73����ڷ�J��r��2ɟ�|�J��?˙�Dg%��KWא���f��dG��3w:��*j,��r2i�E����]P�m�L���$�)KP&f���
@F�^��6CR���L�b�u��l�&|ѱ�V�� x{
"9D^��fG"d=�?�"w�a�&�G�%����Z��.]��mp���O^��=��Q �8��<�uN�؀}�2 l�+f#�m�:�ރ����J��3�2?IY��M�
���ne�/e�!˾ŝ�.84@aw� ������PVM����kO��^�/<d�N�5s�9N����e��O4�Dʹ���C�&�[y�D�@�[�(U3d�	)- ���wgb�A"����Л�o%�����>"������C5��]�N��b���ŇL����:(r�����%+j�,����SH-��_q�g����G�����m\�ƒ�H�tV:�5E���CP��X��c}��ƺQ�UyiA��an�ū#��+��R����u]* �{�: ��3cv2����bTء/�&�<�"�/eP#é	��+��UM2 �a�&�5�vb@�p�]�dB��MZ�)P��������2(��8���'E���T!['���f�ɪ'@I�X8`�{���@�t��A���[ǣ���o�9�	���f����X5�9�/f,/����]����f�J��Q|c ~��۰#< 6�pF�ӂۡ�I&r���ȇo�zxx�DL�Ɓ����*n�@�d/� (��5$��q�b��S����̤s�#�䝁�,��u�K��MB���-g����r�M���6�ۓM�p����7�S�hܦ��i�����g�1iN�fH���~�/�����LlaQ��L�.b n��B��i�UZ�0�i�_��~�V$�q��H]������EIxD\VXԣ����OJ���ǃu���dE"|�?wށ��[ZϢoR�����ֳs�i�7t7�	�-o48%�u����n�YH"�k�Gks7�6�~�)�� �jR���/�FP��ԓ�,��I���c��csĩߎ,}lo�yys�4s����4z��\tw��l>��6���+s{����$����A���!��ɱ���ܤ���9��zUX3�q�.�����_���n����o���2��S�Z-�L��,�%w�:+���O��S��BXi�;�����d2�P���t��X�R4��L�Q�/dL*�.[+�د׉k����n���g��&\ ��Z��-f,Mcv*��u9�l,ǩ"a �x���,��o���Lihii�|}�
�T�C��+U��RC�6d[���\GK� ����1+�f,wsiqY�[����	& �+l�
<�"-��9.b[m��[\��^m��lP�5v�$��;��'������U���M�����	-gK�W?U}�7��Z����BSO�Oa~�^���_�%�W
�[/���w
@���A�;l������>����6�y���S2�Ѽ5�Uv���ԓV���bh]7.Э3Ίy�?7�'��c��O��K:L�7;���,���� ( G��bo<����u~Ŀ�;����Ŋq{e�͙Ok~��avO�BK��yuKy���IɎu�s���A��Ϫ�G(��vC�f��#��a��L�^'�\p]	q�yk�����rצ��W=��s$W�jM�Rsӆ/��q�W����_�g���Gm��Ϗ�Zm�r3Œ�O�g������@���E�e� ����C�T5AT�"��@j�;�rx�qY� [�L��P��+00��u޷���-YdksKNj����,Utu_�>q|� 6��;Ώ�B��|yjFo+��*PR��o���82Nca�%���sF_�G:��#����rc,^��v��r���Q`�s�������]Di�����l��YV^A�#�����[�_-k1�@�{3��������(���;�ަ:}G���A���<ۅ*�N���~�D�+P�1@��o!�o�P�S�!��f��ld`R����ϛc�wv��]�5j����=�����E>r��b�&t֏�9i�[�>3_EQ�7_��46��ޫ��I\��F�Uߜe/����A��7���k�V�����S�Q��DkCC+���9�֫���`��������:����	����� ��5�����ǷA'�}�^�|{6��=�8D����d�,�ۣ��.::�����ͧf��c��v|糭�s�Yǝ��2�jtB�l���1Qr@s�]��'��焪�VA�ˤ��*N��A�r����hu�q�­s���EG6fj�꓏=c���n^CP�8��sٔS�����Y�;or?@k���@eOA��e}�'A��o���	���?����A��M���Q���-�2�m1]�n��Q���w�Z|u������͑�H;K��_��{�-8�J���Л��sް��wD)�!��'yo��Zi���
T�}�&����K2��.�܇����p���эq���������a�K�)un=5�Q}Ae�}p(�)ߘ�zĸ�Ɲ���UY�Y��T�5�C������8k��ě,�B	W_����=�����1^�~�U?�(�c{���7�:�L-~TGw��R��u���I����+#��d�T c6wa�e� A!vD���{@3����At�����ʟ����~�ũ�=ٓ!oU�ۛ�>�@�A��^��~���)u���O[N�8>@�6F��҃jbﵲ�������X����'�N>�X�����0�c���,���wCtV9��7��4j�v �_|Y}-tn����n*������v큸����V1a����G>v}�2bZ�G}�?˿����Ϯ�������0�N+�&Ű��҉*t}V���~�O3�Ker�����'@|=��V�矞��kL={O�Gh��%SdT׵�N>�yB	�0�`�v�����m�T��8�DԚm����S�_887���MU����F�o��!q���Zn�aN�e�@w8��[ҿ�����Y����R¨���vBo�%���yW D�!� �eQ*	�gi�Y��9���l��T��I�>O��EA��)��U����^��7�C����#[ǘ�Ҕ��{e��,`��rL�����t���Y�!"+�ɱ�� ���ڹMQL�B�k^�߁����5)T@`��n�8�'�7hZ�&�J��l����Lwd����r�H�{E⢽7���.�&s��K�;��폤A��=M�� r��H���Jhe^:���s}�A���J��e>M�I��E�P�^��gs���O���qv�`ߝ{��8�^5��z�@�D����nM��R�����z9��^�8�;�+��NǶ�)�2 ��5{Sk��9Tv��sӶ�=��[�B������nW�$��;�x��=�#8�Ы}����@�|�v7AVs̮W���C)�}�ؠ�����#���n����4r��$$�இ���?�k�R���A0/4Ͳ4�6E:� 9�p�fS����_z[母�&�;���R>>�ݱ�'�'j���6�E2���,o���H�Ɵ�O~;F\�_8��3|�8���^�`����ǽ����P�K#6'�r�7����a��а����o(���Rvo�w�02���Ĕ�2}7m�2����i�1b�qT�N�EO��{�gS9_���N�BdM~D�c�E��9��O�F���@|8X��>`j��k��jP�����+���a4n i& �4&�rs�z޳��̱\մ��>�ϱw�������wCYC%�����B��5�-�k�n���0T�ԥ��v ��}���I�߽���NR�M�k
�g�����:���t�X� E���^7'�r�L�f���8�{��wH�Y�q�P��mw߸�C��z[�ȿ�x���/%�Ma�CP���m`T���ז��1�O�A��/!������ 2���q����ivM�t~-%���#���i+�T���\ӿ{�a��kx��lnݐ�c�Q��n��q��ފ�_��b�,�L@B�F<8("�x��P��|,��}���ا���������`�M�IY��,��DN�X��4��E��.����*6sA�x�n�w�B��^��t���	�鬡ʲr�l��C^��*����ܜs;���l|@>���W7b�.�,l.����ZB5�p�z3x�ov���V�jZ��\�Z�<���ޖ�`�O�3�f��A���ֆ�f/�9��j��4��hNLv�$},���-����=��ٜ��k�Ǣ���L�tu�b��ih��ʷ��_���.Ao�%�*[�"Pe�+H��rߺ����U}�!�PO����Z�sV=���q���z��T*�L�Hk�%��hV����~g�.�����Y��L}uT����"�H
()R�A7̠��tw�tJw(J=)�� � �5��м3������`��9w�}�>����}�T2j͡Wf�\X����v2����1v:˥��y��F��\��䢒��#Th�)���a��F���:�������RX֪�$I�y����@���jB������YU�0q&��'%n,�&O�[�qm��YE}�:JUdX��*�|[z��k.�uk�0\�����"�x[���5�0tR#��CW�j�ʭ菊�	��t�'!pMdɭS3'}e�L����a�_~�v���O��ߠI�Y_.��z�i��������f�%���V���pw���:���Ҭ��u,Z�F�Ӹ�|��Y��!���60�L=Z{r(��ߒ�/��67��n=�x�V��4��e�+L��^���7�ݭ���A�o�F$�a�e�|�b�����28����m��>�榬�Qgǿ�Ԉ��Y Z�	�/��H�dE���dG��Չf>�Gc}�\	I�k[�?>�0�c^�R�?�0�%��
Mŝ��F���
;���Z�ɚIW	����]���S[UEw���[�:V{=�A|���f��:H���Ϸeav�XM'����|�3;$E��8j5�t���Q$����l���;-,Oz���(��ߏ+�7yR�_��r��(��=l�ϧ�:c�@ZA9���������b������骛���ֹJ���-�iV�e��k��gk�+�%�oht@��h�S������<�u:�n�q�[�u��߮7o�J���&��W�!�Xٙ��e/��
i�l�Lz��F�W7�y�������
�ឥY���	�_�[�*����5R\�p�f,I�b4�S�C��o��29�b�3�*죪�Ϩ��5n��T��P K]鋫�G/�S�]fb��䡿��gs`��ÏF�5Ė�<F�,�E��mN��� ˽� ��:������v`�]�_��� nR����ǿ ;6���?ΤčVٖ����e{�x\05�1gL�x*��Z�w4��c�m#�96D|hG�:fѲ�k8���mp��#j	D����ԛI�ߡ��EQ�ؘ�i�ո��=��Y���9�moI:�6dI*�ȁ�"O������(���'���Uq��7�/��#s�/�Ф�D�`[!g�肘�*�Ǽ�Y&n�,7�y7���Y��uhh�Ͻ��.������U+��=gF]c%5��|����䣦�ԁ�����x$K�[�6���cZ�Wώ�ל�<-)��|�٪a  +8h����`WD��ݿA��C��[��_�&ؒ�cx@�!���C��5b�/�@kX��Q�*��J}�ﵓ]��f�{���noq�U��;24����U�d��H�E<}���R]�]ޡ3��r]�%�4��^v�����X�Y������9���pr!����rB㫈C`@7�828Z%����y�1���]�2��ܙ��ӧ8��h�����	փOl�O��a��0�������I�g{�p���}	��V1���Cmƶ0�`�u��+�ž���]@MP���;�XO�\~���'�X�n�R����l����' i��^^�#�^�a�ZX"���	f# N��}��*!�X]}|t�"�z�*��f�N��1
]8�����FZ��/� ֨��`@t��A��������b|��HxL	n�S�Vd��e�%%%��t)B���en���/�F��=�4��'�f��A�#|Gw�i��(L|�~r֩}���N�5������槑�9�G�7�F���)>g��O��u[@I�k�7-���x��i�q��x����=�D]4mZE�����C�.�=���4L+�a���9
�6�P���W+�k���BEmDM���X�ؕpx�O��J{S+|LÎ��n���t)e����Yx��s�Rٲ��-���u���G�<T��Gއ�/��[�o�լҍ��1�u�o�2j�d��;�]?��t��k�H+�J'�z���B�0k��u�9��{Ew+3�b��3�m��I^O����@/;�ܶgl�!>�H�磔K��I�A^�(7��jQ�!;�&0���i�a�Z
m�nǅ�Zl��o`�Dg�f������p�z�U�"�O�k��%��Yg&[	b��٪a�����}T���ly'=��2�G�.��z�)�ߑ�1:+`|��tf��B؏m���ڣ#l'��&���l���A�,f"f���#�Uq�[�� \n��4�S�ssM>p��~BG�Py���Y�W~���\D���$����aQ�>�:L��(u.~.�N@������Tzr��<㋕�U{ʕ`ԧ�|?0��t~/��.Ռ:� 	��y�k��Z,��Z��w��D�0N��s)�=iB[.�S���J��1�V�sS�j��׊I��ϛ�!�[6��вz@�����&���7������� n[|���F�����6?��cG<_���Z'���6�(�^ǑD<�j�X�-|3
8����G�^\l"���w����_]���5]�Ȣ�!�c��|�$Jq�>%i��5��%7Eǝ15J��:i��$V= B�~���Hi��� l8��Yny&	w�e�΍'c�!�=�^&?B�"�mw�33�����i��s��g���%�2<�Wj�Z`u~���'�+D��-�q�4?��X��)�I���E-��i|�S%��+�r��`qs�P�vk} �J:�n��k�����[[�/��w�)�����9p�M�n��L�����2��WSl=	.~����&�(���>K[#�SO���]�q�<���L1	^rzg�"�țV|�Ӱ��#��'e�ʑ�?�K��u�a�ͤLҦ�8�7�����J���X�t��d0ʢT?�q�_$Ӊ��Kx�bRw��� ���&�N���G��tMW�<�5��U�;P��)F����b�*>&���il�cV2s���L;0��n�d%Qm�r������@�M��η,�4q��B�_~g�^\�	f��x�V���*�p�$���ʎ��Aq������/a�:�x׈gmEƔP���5�| Շs�̈Z$���zM	?�}y짧e�n���n�� ���HB��׹c^�]�*I�h5�.g[�Bwه��gu.��ivT����d<�0-�/�VuU ��C�?^����=?�'����'�[�����M�ͫ+������̒��{�nN�*A&��'������_�<s�l�}�K�M@A��o ���~�J��e�qB����^��=��y��M��ViB֝k�A���4��_���GS7�e円��<�>�>��{� !~1�H�`�_�(P�а9Υ�ٙ�9��t�J����n����B��è�o�TU��cu��Рgs���7]�QP�Q�訿�-���}g�����|�pSw�[W'�k-.�����I�瞦�.��G +�p�A�. �����}�oޛ �K�R�&���y<�����0kk��[/�D�*	-B@��0���>5�du���$�S~��/�*o��/5g�[�G��BhЭ�h�0�YJ?�tȲ����a�� ��U1qz0���D�$w�����<����.�]2Fy���_ZT�t�t�Au�Bg��oMS�q�������y��7���Zx��z�@��������νd�(�̼�pԢ�I�N�@��R���ɹّ���2�z�1w�2F�1z� �����	(M(���t�h=$�J�N�n�nad~�O����%h�����f7�B�ciQ�y}�adEr0��b��1]�؋�����D|�{[��$���*U6�rs��\#M�BA2C�c�o�\V:v�m�ў&IJJ�� zܔv`Z��j���;�y~��:H�S�ȍ8)=�n�5�q8&4�s��Y�?|w�+K�����ϝ*�V
���:�I�ѡa��F��'��%Z�"��,YY $Ȼ�'r�6�(�G��B���)�f�zv_Jό���w;�������F��%�ЗB�.-2���kNCQ��q
�_	'U���UA77O����8>TyOm�*���S֗��jA�P��-0��Z�F����QNH����\�ék��~��D��6��S��~ܳ�H�����0�p�,@��]$!y�O���R^��%�X3Et�X�l��XԞ��^9͞P*.��o����6o���<iR�4����o}�密2���1�B �-o��|үыjHb��A�T����c��]/�Y!��op�4��rE	k�I���\Ć�2S`���D5����$/��'����/�B�{M>����B����g�W$z�l
BD$8�1�:�Z�=��o���l�u�P��f��!9:�q���?_u���B-�mΛ��L|I�ܠo>��( �����4*���&TZ>�K��4�My�Īc��g�ʻ�xJ$~a������C������aBD�`כs��N���B��L2�y{VIT�,����t������eG�	JV#9
*�a�hG=�*��!�j�qs������-�!ۓ�wH�|wO�
5,Zd�6
&0~����ʅ�S
\��9_�?�&X������<w��uKM�6ۃ�=g��7j��ҝ�M$ 4V�4�F�D���[���Q�6t��'���\W�����;j����ѐ��wc�پP�׾O�8��MB#��J��f�j�j5dy�G��9˝f�س[��=��rݝ��HY�E�rt~��5�J���*1?G4_:*����������p���<��,�ou��Y��*\ �4!"vp�W��&��8#�V��(fm��l=%�~�PK��v����K��D�0{����ie�ת�<���eb����f �H��]��7e���g����GB��h����g�-Iƍ��[T�]�x�@[�R[�W����Sǻ�MoZ�&�7.�����N\�b�êUw�c=�rT��H��o��pKM�$!��ɲ�@��L/�ebv������-z�e� դ�!�J=�{qAq	X}4�Z��O���NDp�?���o�:bj~Ȑw�0��9[A<���fY��dY4�Ӕ#�zb��P�ypV�y�#a�̏��J��x��;����?k��I��R?/���ލ�POc��2T��=�&���9�)j<�1;�tj ��N�?���/�X�t?LR�y��7C_c������z�ʹp��L�ʌ�Ț������~�����C3ϺCe\ˁ`sn%u�xL�n�����Dx�fQ�};p��k��K�j������)1u��E[�����;��)��Zx����^�<�ѐ��E�kv+=S�q���d1�=a�ng�28�0�����	���8��>5���a�&�qL�.��7ޟpӵP(��3ӥ?+T<W�B��6)x9u��H�CK���°�u�6ܽ	��z�����+5�����>*[�ʾ��
���%��g1���y��s��%U�����<��Q�V��(�{~6wx��dόώ2��^[&s����C�Ky,��|p�����7?,Rˬ�g<m�gF��������n)�9h%�� q��_nU�66y���� �U�޻��е��93|��]>�A6O1͎�n�9e�Q��ez<އ��OE��3�kAXXT�o�2��9�~�OǸJ��W�{oy�N�KSML�!؉b=}��S���KE���џ��@�gȚR=n@�x�����]��{�{Κ��A,�>�&s��� ��O�7;�}��\����<��,��ȉ����D�j��9�x㣧��i����h\�����u"a��� �(��V��R�������1�.n�� @c�}?c���H����@ �������(�l>B��bPq��lg�툱+�8�����)K�R=�'9��K߅���wZ�B���T����J�>�xy71"��w11̂�7>�~$^_��j�BG4w��3��*RE�|ӈ�
���>�χH��b���^�Ւh��`��M�PQh���@�]ԗ��G�p5�p	�$y�D����sx75�P�(9!s�:P�|N%j;�@��|��,Dx�Ӏl��u~L�?�p�T�3Y���/V
��q����뾝X�Ϋ��exϸY�� �R'aQ�;;�Bl�&���g���6��,�۞�TSB���G�:wE=��i�����,�`ؐ�T,�#ۯ{�8���d����\>���ج�Up�b��>�ي��ؾ�)�38�w~V�GM,Q�=���S�.��um�Xvi_~�;`y�R����x@>�z---�!L����9��:@&W���r������O�i����t��Yg���E�AC���RNyN�.���Z�lY�][��aZE�!V��2$R2fJ���2�%��yC�
J����w]���sEP(	
Ձ�ɻb�J�a�q��zP���-Ň|��� ��;��Ѻ*�"�^���Fk���f� 
d��	�z9s�F(�\\\�"����PBv1(�=i���<�[['���h��X?!�`�a�<�nXn�?�+��gI�ob�ɲ�	Lg�Y6�����k��s�N7���6sc������+�v^n��!��"�������K�����F���	�����H.,$us�'���$��y-�$9��z/���t�u��e�K��,2�GZb�jn�_5���sRF�?X�ϟ����fR�;�*�L8�_Г>�w�\����ͩRx�pM��)��0h���]�<Y�B�N)0e>�� �sq�Cn&���b��9j�k�9���&,ӓŶu���#�?�Z�?)��P�+K�w�j�v����|�Y�Uk���:	��A4�]���2r(g� ���~�1;˩����)z�p�N̅�U4�=|��#�Ȍ�V��9)K.Ki�o�j��bS�����)��-���و��ʉk��lnŮ�[p.���)�T��ц:@���O��]@c��Y����������V�]*��-��8�)�Tio��K\�0���!�������}E��w��=�j"�W]�������?�<�y�(G�S})���9��6�&>Z\������&��J{=be\s����:Gs�X'{�F�^Nϥ���\�V�~=g<��w��}�����]��	F�Z�(Jם��"�c8)��w�Gq�.��۷fmEOWH\��5��<Dx��K���id�i�`v0ȐH~�����?��^k�fu?;�������5��;z�9��b��\����Ms�w��;N����Q���F���Z7�Nm1.�88m��E��ǭ�p� ��z\?N��csmqX��<���pԬG7�.
?��3�3�!/gý��F�)6<�B,����:�:�%���6��4;o~�q{۵|�����='�]e.�����[/B���F�����+�7�W����D��8z~��P�<"F�{r�E�L�^���?��,�"B[V��M���k{�Q|_v>�4�=Y
ן��K_2���G���⠹�����}�$�<�9NgrҜ>�|*[�8ⱗ���\����h��Y󉵰�BK{,�z
���\�����{X7�z�A��9G�-wU�)zF�֪����[���VG��n}�efu�Ё�;(��B��!r׹-���հ�\��s�+:!�,�*V��Z�N%����qxo
�hJ4�����z���L.���8]juGM��ŮL��Le�y;� O'J����~\�-�y҄�*kZ��XsXY�g���=��_dJ��i�E
�������<��6�r����r��T7xQPNFf�Ƕx��k�y|�~\>�{�%�}��9r���}t���V�413�;�Vvo/;��Ȉ|�	vV���Dma�	?�,�-pk��3)**�\�Wr�I�#U܋�{�Y0�GQ�K[[[?�>I�������j�Uk�m|�`��#ח�f ��q��]�ⶦ	��Z����t��_�IJ���#z����J�۶Y���� ���%w	0X[q��ȄSF��ԳW�"��x�'�
v���������{�w�4�x�t���Z+猴ܳF�}cw{r<�V�*3��`�h8����W��ӵh���sW�k�-��M=���Zv�+$�NR����j�rA�	Loc��
�Ə����(�;����D}���3k�Y�
kMp1�NY=llB^Sy�Ū4�en�E)���A��Ҩ�}�	q�kY���E��N]Lk�X�l$s�.<8::��(����=���K�C�������q��tT9M�"�*��1aĈ���G1/.|�cɩ&��kcm�[�X5�F���7p��+��\��t����7:oȟS�?T]n���'
(y����5�d4����ܖ��C�y���g�%��Gh� 6�2,k��۳����)��nذSF��K�x��,��H��\�� �.�l{�	��p���H�R�~n�����rlIRNG1h�7�sb�+��uH{���I��v� �de�`T���j�6n�����Ȥ��7_�܆4oA;Nw9���Wz܄��g�ٚK�Ӽ���y�Bu���e�$G�^4.�"��."b�%B��:������S�ݯIVs̽�iim�Ĝ��bBk�"[��O�1��o1�I�{�����aHwq��s|��-sG@�3�e����cL�����Q��05��u���N��.#P���3:{�����L<*����2zhХ߼N��!�F���\����x]����ɇ�|�A��Lm����cqB�V��bd�є�<$����$m�I���d?'����&���"j���`��1����OQ�K�`��\���%��M����s4���Ǥ���4Vc�ǵ--���r�+�Q�z��d���wA`�Ne@(�7ȑѡ���(۟%u������KZ'����Z~f��R��较B�x�s}�c�s�k�"wj7�J_Ǧ���.��/�kI��STId&|���9��u�J���f��\B�T���v�J�DAþ�yƤ��j� N&�ŝ�^j��NO��p�(w�{���tَ3^RCx!�������U��t� ���q�'�X �2p$���~��ӆhU�R��Ɛ*�O�efZ�t�W����i�4꨼=i��b��@k8�E"?���=<�*o$�N4��n{s��Q�mM���K����v�ræh����d3U��.�J�Y��A �aB�/�;�9t*�c��էMLW_���Z�@��n�95!*r��D]mm�|L:8�h��V�o�������-��~h���$�V�}���͌ڄ������ח!A%Y�1qH��"��rЫ��gl��S��Rp'���8FhI_ɍ����#���H����Y�׋���8�L0&��q��G�B���u�L�D���u(�������5~���7V*N{<���*I����8)J��4�r?ܶ�bL�IEY�W��woV�����]\Ȋf:E{8B���,8&D���݃�7�,��D����o�~����)u[.�)�c�M��4�K��"zB����:H�4YЋ4ϲ`N�����t����ͯݖ~*�z�<b��5�J��ɖ6��-��/RA��,��g��tw��d���o���S�L{e��������]��ZIp�<�&u�r[���Z��y�ڿϘ�
&�~��Q� ���.�۝2B�{�\��� ֖G��%u~��@�lrÞ���XI���×&qbP-��A��������V�(��[ac��p�+�"�ֱ$X�.�+>���)60�r�c����j�V�l{�Ԋ�$ ��<>�q�s#��:� �ͬ=�!����m�8���c�߬��_���?�t�#��j���~a����^��гB��;�i��v��?z�x#�ECM³syL���m%�C^��u��B�?���O>���Ů	W��0��n�E�wH��_f�t��
���.��>C�6���M^9dW�b�L�Ѭl��F���<N�܃�(�El�'bca?��a#	�"^5M�8ڥ�����8_�nv��E���!���7���l3����kK]�q���y Jje!��f�/���=����u�Y��"���#�F(ϲN��g�``�FX�"�A���|��孖��J�v���0�I��B��i���'}x�gX��E���h4ѡ�j�E���4o�O�rz��{�������@���r�3Q�)5Q m�ʊE�W�{3�V��[0Gq��0ԕ�a�R��̓
N����q';R�U�~g쫃C6f�GHG;��(�����Q�~W�.)�p����?_h�O~���E���`�3��ˎ���Q~1x��=~����$HLg#��zܞ��]�F�q������h����tꤨ"���^!2�7M�%1$�Y�Fʔ2š�����z��s��uB�}���6��qf�o�����:IDt��D�x��l��2_"���FV��*�����7�o��z�d�d_���j.�d���I$���"���?��J&�]����ڲ���uXGJ��j}��:&�ydV��6�QuM���Gx��BC�=l��(���-��hS��2���9�yD�̆�6I�͚�4���| ��P�ըOW�D�5��ߕ��OT	���Q�]�GW�悒�N�0�^hŽ���9����^�'!�������B�~oV[n���?g��*><��q~gE��ҥ�1{�WW�T�<�@+��ot�
�|��I2G[��Z���d�Li	G���c�:
'
3';���Z�$�>x�V�;�����| ����\h��lڞ�6D�9����R�����=ȎS77��e�jq2�Of��p��ޯ���;�d���o4}���K���G"�M�3.�{�a����=z�����F��}����8I������j�h�Ar䍻�����KS�Ompk���W��Ï��D6[�%ade���Q_���lZu1��E���]�l�����w��
��a1��؜C{k;�v���J}��Y��_ǡX�ѯw�$�����d�ū��B��g{��J|ۀ0���o�}QϜi3���Jo��a��!N��r�JD�DKR�|����V���Bq�D�Yֳ�jɚ'>����	iY��K�R0X����d��~|R�+��ڿO�%|��s���}ٚ=��y� �?��G�c�i������X�(M�p�e�f.{ؗ��(�ٰt��><_���]1,!0(����� �X��ٓA����?�Ur�=O������Wz5�nz�z.�@��v�5�]!�a	˗4��N�2��)JN��RO]TdO~�>\�A|�so�����4��Mq��,^��]8�>΢�f�����ǂ�$��s�E|�zm'�0�S�]4��g��7��@������l�K�ċt�'�v��ݶrd#��j.J��a�bv7���+��sr8��	u�����ڸ���1���y~@U����\6'ɏ�� ����Cw�s���0��5S�K�(yv�o�ML�}j)����e��+UAn�맫�ǜM�+[F��!;k������6*؟�`�p��B�L��*W��+�&��p�ϯ_�C�*����Tq��ClMt��-e�kϤS��1\T[fwgtu�c�GH�"�J�(:�C7���T��W${$�y���h���A(k�h�rB﮶f�A���矍Q�¨O%�a�1sa���`���c����?�um>��9\��;E��J��*�Ԅ�2� a٦��)R�'
k$v����e/��u��62r�"��P�:�Vs�	�FG$2QQ�Y�i�yr�BU$E:!��Q|f���:]|����s��f�����q���}�u|����,C������}zU�s	�\��9��m/J|*�����j��(6|���e�_�����Q��U�ϸ1O������_��Z�t�M����7��X"+�CR����s7�c,|�t�*�"�^���ǽ��X�K��l{�|8W���i�`��?6�rP6�u�c�6C-�?���7�.��υ!C��vm��	�B9sp�Z�b�q�'��� �����!�+�ytH;|l��*���һ�4)�N�w�ӱR'	����[���(ɛ�����z�K�O��?�@�`�t����'����>U�Sy]8{�ˍ�X@Y�]��ׇTmΰڊ�/�ܝE�y<s�Fv��c�=���)��- ^��9�b�e�� Y;��3�u�?u����|�(1s��<]t��Yg��_�i�O�]KV�,��"��7*d�5�?�o�Z�"C�{Mf�+�US��٧dh:��(ج����XA>����,�7���م�?TeN�I�G;_*!@\QKi,؇-7�l���w��ͦ��q�[H��u�P)��Y� �d�d�� �0�L�=�d�Ȟ��m�8�����r���~b���!!2���=������_�+!�g���oy�92~})����M��<�^F/�b.37������	������9�a����#Ł� m��Ϊ�(�E�8D\�S�U.��*����mۘ��т��N�$u�����ع3�y�P6@���)��om��ϫS�d���Hѕ�8�W��T����u��q�iw�U�QD�u-g������!�໷'&�����$t�g�~�r�l`S��w�f$�p
J3�F�g�녀�H�c�G������v^{���-n����rm`�������t��)s�쬎��xAL&��a�N���0>��̯������p���nVgK�t��%#D���Ƿ^_v����h�����/�J-�s���#�|r��X�{w����.��1��͟�h�W��z���e�d��M૸��]�uc�
�ɔ��Vp��u���֒���ЧJ�eɳ�h�������'���u;�0����Q�V���ΰ��	J�a[w������u��<ʱ�Sq�ʩ��(4"+����wg�DRl����U�`�;e���k�{���x�l�{�I���I'듨q;3_��7����鱒��4�(���j������!{=������%s`��KTug��-�{Rњ(�����p�=�����K�pX���j�qWA������&��Џ��Ct֫�~������h�<�s��9� �H�H.cnV��>.!� � {	7ec,Ó���al@�3'��R܉�;��������E,�b!"��X�ɛ���\-�o�j��Z������=<J���I] y����!YcG����9Ӳ_�ON�a [>V�X�L���+!��=�	�(U�:�p0�;CW�Ҫ��mz����V�n�(�7&����v���{Q����u�D�1�Cs���w��(O�C�c�^A�չ����?��;+7w�\�7oBE���\)�D��2%�s��n�5�A1�l��:
YZxA���c�Ղ<��7���ڊ�w��C�T�5����v^'�d�+l�]%O�sS��ս�P�ި90J����طB�N,�h�vɳ��K��L0�<�~u�>��y_@ό�5��$�����%���+4]�Ⱦ�݃R!��F���Ӿ�\�wD������6�����]�/�����17d�E� u������s����Ƀ���Ҽ�읍rJU�H"����1r+�ą(�8d���m������c$��͖+����D�¾��R�T�2����[�u݆+�LN�H�L��Jr�W�y�+���>&�gVZ}%?�>�z�\Dn`�N�2����!��A#��3���G����\�q�/��v�J�J�p������zȶ���u'�i�������Q��a�������j�z�u��}'�J]��l����[
YZr{m�+�]�h4r3U6ڱw2y�vny���	�Ő��X7֌p�<�����o�!{�r�tn��9X�`5���Qkv&)Y�����XA��: y?�A�o�,�,�3y7��1tE(�U\OM�E�[A�^
n,�����M�K�(>�P�Fz���Z�鋮y͏��5Lǘ�Z�8���T)7Y����O}%����F�60�_�3���V9��skS����g�m�D37f�-qmB��"ĆZ��_���.��"z����%랥Yi�.��^Ail�a����F}��իv���\;1v�e��L��o�!����Q��v��y��d筕�7�z?~y��&<|�{������Mw0��	$����M���Ȯj`_믁��FA�k�����3t�OA���e�(�w�;]y�Ӕ��c��{`692}���D]� J��,	 �DX˹3�f���9��N{f`�䌾>��-�������F�Ǒۻͧ)�{-±Q �����Z;+��rW����o�g�R��Nv���s� ��YK��A��w�*׫�����D?6��S�H��{��{�%d{+;��z9��m�t��U�jd��������-��K2'�����ٚ�p-]�nİ�����.C��㸯�6<�_=3�?O��Z���ע��ڕ*Œ�
=ht��r�-�m�w�p}�p��z-�p�CWeJ�j�B�����d`����ܓ��:qC]ݟ3[�����X�e4�o�oG^_ӓ�� ��s1-xݰӐ:pxprJ�� R�0�F��*%�q{�{�S�����uh}g�Zn��{g�O>6�hiߓ/��~�0\!�96c}i�������*�	�LW���t�?B�z��;q�Ĉ��~݀��\|4%�5���Y:�vԧ��s�Β�E���^��U�[ݐs,���>���v��@aY03@e��4U/�y��j��jb ��r&_�o�~v���|���*`�᪖�}��BV5�ǤK@�+��k�����58' � �9����d��pF8)�_�_'_�Zε��-�A����s�Ng��^b�O��Ԙ��^o__���lM�4\ː���M�D{��5��z��L�Z��^�����n]�O�{�}��`o�L$����5�`�W����E�H�G�?��z	e����|�(�h��	����(>cuG�HoQd?�A�����n�+���\C������������v��n���Y`�۟f���W�ep�'�RÒ�
j��>j�{b���f 
�U���N�Sb���Q<�T���@�k���F�QƧo�/�;��z�Q[P��j�&�>6ӽ	�A+��e]@O.N�h��` 
y����������p�� �ba6����%�ݔ��4��/E�ޚ�
�z��"���5���WjL2�˛ϊ��d5��\Dx��˂��a��1G�B{������T�H��j<��0�8D���4C��@�Ã�/���9�쥯��1����z�����q�%#�m���̜g\��:İʦVQӛ���w�*�%�	�Ś��ry yS�J��xD[J�^���Z����Kv��n���"�[=*�;��Sc�W����k9���~K��^�0k�O��ռ���1'��1�ҟ��Ő�J׬�l��k�ix�=:8�ŏ�_y|��&E�L,����(i]Ŝ�kߖ�䥩�ܶ�6s������;�� ���x�0��/������y��B�l����:�ɆQ=�Ō�f0w���,wm�"�r�)r�ss�KU%����!U�?�����_���zQR�L0�v�s{w�uڻ�%����������]D�jY��5m���Q�/�^�D�����(��>��S��ˠC��:V��]��e0m�,Y24R�#�㔉b��F�����h�G�yO
RD)����1�^��ॕ���k��.ׯm}���H����_�/"bQxm�JMIᗒ�nk�c���446q'L��1Ȓ��FΫ4�`��j1����+�S���Oa�L�M���P�Q���/���0�������R-U.!j���/E2����{�x�5%�`f3S܄��u��L���͛�<t��ggg�|���4V���]�t5T��!�k�A�νϝMv��u_)v��^���~>goP!܁JYu�(�)����[@=7�~�;f�s>��bv$��}��Ȕz�?�^�G|���#lT����X������1!b�U)D��ƛ݆�hE�0$�>�X�4Q\y�x�\���Y������ޜ0sC^(<(��˲~�n�FS��S��G+O�4;�{E�E���Y׃���"R�Y�ec����`��_�K�fu��Z�H�)R=�s�M������#����r��U�]3\sv�秳��z��إ
���-T�-���~��� 5L��[�o��/�����<�I�OGd���(�].xܺy?F��;��m�02�G��-�oaoA�Ӂ���w�ߍ�+#�n�����-"���]M��&|��!ZvhR�
[.^r'���N��Қ�����Qi� �^�������s��Wt}h9�Ӷ6�k�� <�#��3ٸh��������%�}5d LR�q���������r��o}*��W,\��:q�?�vK�$j�3v�9����"Q��_#�|a!��t��9��
�U{��_TT���,��~b�7���ˆ.;3����:h$�B�����tb>ӭv��vfS3��C2�P!�!���XqK��r:��7-Q[�/o9*�"w��ܝ3b'5R�����K�cm�5���9�_��:˄ֈӃu�3��u��~d&�rl|�`�b����Z��mKrwM�d��F,����mί�:�Z��-*�c������=O��ҟl��n5G&���k�O�i0ƕگo�R�����j]�fn��+�D�`��D��O�7��No�j�>�Mi���c��~���P�,{$�$G�Ǌ��lG�
��������Q�&78{�P�q��͝��{_���~���ǽ_���9^����K��k�r�R� 4F@�
�q�c6���e��j���`@�A��/�d Y�㈆�4x
�'_f�����+��ѷ��R���ܑԢr�Z-.���6ǻZ�w^j�+|�bjsg�I�� +"��٠1qgh~Y_$��w��=�lj>:#x�i�3����p�����
a=r����awF�!P�٢��Bi+��x�bd�z#`B�\t�X��U&?:m��djju�"�t�w��Uϭ� B������S�OvF���rNk+/oA,��o�7{�AU��v=F�)٘8>)��Wy�'"���W��eQ���6�堜&0��("����k�'�^=����m��^N�`�5��t.�ez�0}� �:�1�:��vM��q�`l?�z�3&���b
z27;�U�~�"t������wL7�	?c5��h�Ey�5���]�5�ps�q�[C�7�z-88�{@`��N��()��F,qᛰ_p�&�f��t����F?p�)۬�v^��%N�
.*���@=%���<��b[�C��w���(��[Q����ۃ{��8����5�nL}����ks��ppt[�U&�߇"BF�O:vUPg�	����m}
�=xx
��M߹���Y�0�{�]w�����'�@�xi%��^���3�>G��m[�\��6���������xT8cUd5"0)���OS�P��`OvΎ�����ي�56O��|x���9�Q��+bW��.�c�Z}����Ib���N۞��牄�y�U�RW�D���Ү�-�L��ɺ�67&	�
BwM��f�P�K#;�K#^T�.ff橄�׎yE���m붌���L�L�sH��;���Ҫ�G|�K��\���kB�M��j��/� �c%��͡���|�Z|�c�f�G�e)�<��p�������� ���[�%�r ��&��K|�tPI:�j9��}w�7���kH�{������ĕe���8AO��%}��x:�DRR�g��v��K�e��%4v-������(4>z\�#���r�bp���q���?�?2��cʭ;w�K�t���p>:F���ɪ)��4aq��G�D�/"JEg�F�5�`1O��u����2ɼh�\v���9_��
jw�,d\q�U�n��;� ˙)��CL��ΜivKл~����(�2x{,�<c�r�de�c����|��K?�M�f�S�l!����I�����х���_�U��N��~\)N0*e/#�}G���}���]�"Y�u��5�rR\�	l�u�ǡN�j?�5ߛę �`cs��U���xK���3�h���)/B&H��昂&A�NU�	��z�6��)��Y���X���JF��N�_*��Av%??���_1A�ߺkP�X�Y�]�*ZhR=����;�|S��EsƢ�8[���]�hp3�̯��f8S�Z'CW~��X`����fDF�����y��:?�#y�^�L�F�L�ɒ�~B���?�<����m�3Xkc�]6x�}v��' �:L�q�,�M7��^�*±�����)�mb�A��W
ȹ��0�(����Oޗ#��s�J������#Z�`z���A;�<6~�)F�*��ڜ�����$� �v���L/Ek�!e�Ҩ.{��ٷq_�B����	qa)|6�`ft�:iO�}�'%~>���� E����ű3�+���<����WY@��O�>��6.�Oz�7�H_��}��^��{�w[$����ڟ^�Vq�u��_�I�R�DF���kE��CQh|�����QL܃���(c>�B	s���+������ ^����܇Z��~�~4���S{`�E�(�#*t�Q��ʢ���^&�y���d#��El<
�i��xG�/�Z�0&b�_{�����U�1���h;�#&m{J-�Aޟ�,�M£�C��J.Z�1Ny
�8s��$5՞�@ϲ�]˅T������Ś�����(�V�ᜮOw������s`����|�n|~��7�`�8����cR���U����^j0_Z�TRZ��un����H�
���S��҆�k�)xa}H?OZ����f*��67 �ޙ.�B{y��x��r���:Ϗ>p`�!��:o�L��:����*QK�w�h�����[�_-q��U�!�HR�W� ��C�0޽�3���?�xN�4��.�����35�� 32�Ѝ��O�8�)�$NGV�\@�5����U������5�^�k����,��ٷ��~ʘ�5J[/��27&0��ǥ2��ON�+X��g=92B"¾s褂(�>^`�r��*Z���ǚ�|������$�ӨL�K%𶼾B���"�U�.�3�b4��tKw�Z�N�򭩈?������<�v�4���`���qm�Qz�\��z�����w�6kc����z;y���L�-���.��'KL�Ψ�8f��Y��Z�k��*6��������.����;��AmRW�3/58��O���q��$���V��&1q
$iM�W2�R0��V��1
���,>@��Z�s����g�/��E�·�*���=J(g?���#=b���)VJ����ˈ�z�nP��;��zqO�����U�������z����_(��1�٭�_�:O������?��t�3(�PB��.�?�@T�HD�&2c��R䂞R�*|~&�)��*h�\����߽�<�<"6T�����[}6M�E�`g����:`ܱg��9�ò�,�m7��ŔlP����u~7]$��L�<,����3!�BSZ���0r6�5�)�L7H�!:T��������gTA�P���CËY:�_
�Ҏ������x]�����,��)�/���WN~+~�+�$7�&�wvH$d)�̍�^�^��U�b]��&�p+����b��j]�v_S�,��=������"�K+����H�{<�l�ȳ��2�GS|ɫG�E��ڦ�k�nP���YlL����c%��޻TO�2����U �������J&�x�q���4;;c'���m�U?0�	�?A/m,���
'����
&æF�^��K���,���I��˅9|�#ٰm՗xȉ�=�J\�4�V�h���)�u�|�o��q�0��W��K���ޕ?Ыҷ�v�5�թj�u� c�b�6��^��_6��>�떨he�/Q��u��20:��.؟�[���o��qx�T���uP�#vǯt�Urs�B��X�n������<|��g��V���z���jp����/�� ��"� �͉_�Z�����H\���=U)#P����~Y��>��ű��n.m��i������c~aP�>T~�����"&D$C	hM�gS-	��%WG;��t�z����<K��*����y��������~4ӿ�W0���\B9��u�Wv�JDH���.n%�f)Bq�pw5�+��[�!��I�^�/�v$�o�ؒ��	�&ؤ�lT�C�8-��^�{`f�v��p�\��i4�d��z���\�d�����rt0�:/s�����!nY�G~���OJ��@ Y���{���L,>�b4+�������X�%b���>1�rD����%Te�ٽ������{
445模��/�C��L��R<��,*��)�%�u�%p�%�b�����:����A�I knOxnv+W�ݠ�<��;		r���v�ZdLV'i}n;�e���V����[$�F��Jˎ�l�q��e�LH`E����b���W,�x'L��[Ak�xy:����Z��n�⋾��Wz��f*�!�f)��t�c�����ܫ*9ε�]gˤf25ă�c��h/mK�{<�{��'��9�Z��:�9�:^{�솿0�$'MCIi���G��|&�8s���b>����l�޿�4�*#XJ��0���\uF#��=�[.�ӼW����ٜ�_y���c!0	��:��&��C�f����4�_:�����R�Q�!/0|&~��j�^ �K\z(��Ԓ���E)9E�?~3���*QK�P�E�.�3�/�2��`8��-�#9E�Kz~�g�� iIڮ�f��-��Wb
�uS�vj�
�XkO�X'ݻ����?�#��	 ���2=NN>c�Ab���~�_i,qbRe�e"J;V��d�J���e�.�o���ުI��7S�c�h443)��r++�u��&�p�ґf�5fJ-
w��KCo�AA2���0���t,y�z��t~Mn�\��ӽ���g�E��LGW@��e��۴�	CM�Z4�����&��~i��.��4�3֦�����86�X,�=9/zC	�^��<���2U�O���i�Ğ �����IX�^��]������l���M�E�~�h����G�ZP�T�׬����L(X*H��mQr5w��J�P���\H4�7����1N����L4�\���k�F�0����:�s�W��,��k�?�f��J7�П�Td���D�0�'��^A��2����w?���n�t1x%�VѶ`V���~�ʕ�{،�TTUZ�ku��g����E_�2�Ӹ{�C*�+I}����J#��ϑ����ɇD�*a�wp�>��q;=+�6��PSU� �{��L��M�a��'6�[y�T)�.�}�%N����)��(���A�4���[zf|���໘�A��7M�$��*��:8���y�*�%���uXu�WOȻ81�%'C#�Z�m��u�����~�]�p��
.J�S,⳵�U҅<Cb2Q��������bn٣��Ɵ��:6�9i�3e�S'�CDYbM��S9S�����1���I��وG�&[�V+�B�?�����A��pgB�v�>�Gƴ�Q�BnΚ0p����E�2��I������X �1m������adG��	��i�!��~�f\Ԭ��w����g}	?~z��]�8r^q5"��S������H���+�}�)�K�g�ӯG��M�W�Y�
�L�~p�}�j�;�U���(�7�\�C`�->˾��w���ƻ�`��o�E�i[t��D���P��Q[�7ӭ�$R�T-�g"PDm��$0�Ǐ}�R|z��W,�'ф��%=�$�rZ���6�B�d�G�ezQ��n�҇�>ɚ1נ���A����x����&�3�1�ͮ�y�%���n��u�Fw͔�rt�3[GRɄ��Y?�@����ٓ0�}\�d&��j�S6:0y��/�]��6����l�;�E<DוM��s,�O��(3���v��<O�����<`��<��mv�\���f�D���,�2�]>������<'��>�gee�x?���8�D[�
�9	;ji �c�<t�B����lUJƚ�R�/����jg���͈MT�!<;g���/@�A�Ģ���<CKɕ�gz8�T�f��IP�}Mbؿa�s���|I%4��Ϧw��Կ-/ȳpGݷ�������s��x�3Kk>�LZ�Ҽ�x�r�@��^���t]J��{v���P������L�P���xX}L�VQ�c'���`�}������3�a��O�����o��'�ՑRJ~í�@L��`�!�(5�B����d(װ��%�H�Zs�ʩS�i�(zL�̲F8�6�$��^�3������LNP{�6)�\�X��P�wF����ȁ���|��d�`��H��2��7��@H����|��8nHПB�|�k���A��� �nl����o�X+�q�*��-lvy)�GJ-�
�l,�r�6�[���S���ZS�z��^!7ЪlO_�ӈ)t��A��/ʞ����_��|$�;j_�F���Րj!��k،CH�H�c�+�r���i�T��P�嫻�c}���
�>iY���Q.t�7�u|��b���#-cp�kTϠn�,������Ծ���I
@�<h����}��go�D�a���kk�d��w6����q�����6�U�+o�FWG�a�]��ۛ��b��0��[2���>	�[�T� Ŀ��?�D�k�YzMV����v�9M�����Bt�𲊊�o�y.l��9g��V��Bg����n�K�%����ӣKŽ"�#>od�����X&o��[�Ք�T�&4��X�8#����/�F\�Hiw��_Hv�>]���������dm��;:B��.����A(eE�_�Z�2���P��xQ���v9W�]Ffk�
�1ͅ3T���(R�O�]#}��n���)�k�-�w��YC\"AK����<_��m��T���xBʥ�ndH���O~d��8qt�Q7����n���[��w�u���X���e�l��zJC�W��V�de��[�=n&$�����msF�O�[-�8]'�碔:�j杍b�g/f��"�4�t�kBc&|0�Z�#NS\���3ӶN�!*�/�9%�ۅ��յ������U��u����Q�e��	����,+r�h%�Z|�L
����e��Z��_ؠ�JT�Ko}wI��7W���		�W��X�Qq��~��Bnd"���s+5�~�0AK�SO���e�!�Bc�'�����Q�#�F"�n�lo�U:Ϙ������H���?�y��q����t!lS�9
q�\N2�?�_YW��$������Z8�����[����^�A�!��~(�f�ؤ$�Ms�2�b�p5�-M�O���-h�Sud��9�-�HX�����+�f�ip���;����;���'Hz2l��ى�K�nݜ�!�3:fO-Fc W�DbZ߷��!�W�m�.{
�ʮMQ.gr����߸������G�;>�(�H��KMO�/����:w�Zg�W�����d��,`����;�ԏ-޽�?p���`�Ǽ�wGGd�c=�?G�G[���������\s��>N��sM�
�U��7S2Q�~hL����w-Ż|�'�^(�n��͢>���VnU�r�H�_0����Z���s�z��Y���HF��'��f�*!Pj��戹Q���B�<������:=��A���Mۘ��������1��Q�p�(W�d�?0)�N}Y7��3ڻh_�,�]1�w/�S�O�1�y+:񼴊�9�ش��.@�m��\*e]����m���.i��@T�}o�DUF莖Y6���vp�H�����B�f�kQ6p4K��ZD,ېm���&,g�<��}�FG���I�O�����[���;����<#t�c\����S�t��hm�:ky��^0W���H�$�ΣΎ�����@�*�������I9J��8,�V���Y(#�_��#�P��~�Qw�Wֽ�-�:�cYgh��h��Hpl���\L^y��B����n��>Ș��$��'��7�8�j't�A���zA�x^$����g6�@����i�e�I�^���q��]��ǫ:c����UI+jQ���m�t���B8�����R������z&y�Z�0�Cjd�V{g�?=��.�q�TkSX���~I�":��]�����4���lUn�v�����~��B�g�̕��5�57�Z�fF7���VTk�3�,tqK��ܸc�}��xS��>��n�}>��H{3�����J���k��Oh��]}��D�d�ݎ�<=D^����D��,�I����<9�<وQ�>U�j�\6n�I��[4����`j�t�O7�ձr�|��j������P�M���ۻ��7���I,��ׯwI��|����2�܎ưX�Kم�o55/��&�� P_�~tTқ�jl�^f_�>�>���ע����S��4~�p�uM�{�+MKP��z��0�>6����^ŷ��{O�&���ϮlQ[�ڹ��ͺ��h���{���%X����^Z�ܨ��SEc�Y����q�Vj���ՌC��/,1e�dD�˙[+U+ˌ�A�����3X���_�ZҤX7��CZo�nD>ŭNp4=��/��UE�� +o��5vr�ן��3�O|irE�nmgNj�.n�z��@��x��S�C������X��)VcΣ��k�mn�jЀi�R�]�T��+&|��h�d��������\u�B<���;�vǬ�LS�K����OhR��~%�u�����'��)���L�����OLd�Ĝ|�_\WB%(��О���.�殛'On�1�>d/~U���:�}��y���	��z���(+֔M7Kǀ���/=W{v)|f���l�&��!���g�Q�q��ɵ��w�5��h���2�0�qb�h�V;��[v���^�w�v�KS��3���	���60��=�$�O���I�w��b<�}�,k��S�L� yUv����#��� ��a/�wV�M��2�`cG:X+�_�������PF����v-��p��Ȼ�N�$N`�n��Q8�;�A������=��\������}�MCC���F��_L▨��β���E� ���!����㎎�Bk$�5��`_�kaaa����@J��ɫ�������`aU?�Z��/���IR�l�k������P��p��{�n���[Ωa������u?�\��G�Jbe���M�z(��*�˖���5��LqeB<�,��/+��٧����	�������L���8$������o��Oq,I�vFu�LB��<�ݲ�@�_e�I��a�U͑���wզ�{��S#��;�캎���>k��o�F������w}�(�>���11μ�8{���
{�e]F��7�ag��X�"ʋ��s?
����_cyn}/����N ��g�Iq�����/����5�^Bl��ޛ׭�b>�ǟ�p�p���U���dMLpQ��JA�=���C�2���U��9�>�$�ײ�ob @g�R6�n�w��,���Խu��v�:�����=#(����7��|e���
�o=���:��I���1�G�#]4cS�y���̀:����+��ѶV��*�rn��i�%�^�[ �AEW��	V��:&^]N�1���l��Xκ�FO��>�V�~�ա77K�Q�,��7���րs���G�����*����1��v��U}s�H����	u��S������RiG��j���$X��LÙ�wD9�s$�?�T�xSj�޺�	K��~�7vav�����~b#��nŌ�u��������K�!���6�׺V#9�o��e��0c�>���']�u���\{l���������B}Y�k�AS��B��F3�ޖ�\)��Ҏ݋[��i��Y�5��=-�G���'Gʯ�9�s�eB�c�FK�K?x��I[N9Z�o7T�d[y���͵*��]9h<�K!���	�?�fF~E�Tp��s�ظ��X���;U\��Sv�7�7��ه���;z(p�KSn�����<�/W�m!w�y?��J�ȼ��v�����<��0�=��������dGњBCㅫ�%=&���:<}R��$N����l0RQv��眿ˏ�^i]��R��t��^�4�]��3	�K��u��)��ąg��y����Q���X	ON�'�w�"�g�:��FWVƐ[����Xb�yQ��ҩ���j�KV��D�ڌ�΅ɭɆڙ�W��6�pZK.��ry�p[�[��*�eLT�n��np��*������µ^���?N��岒�!���%[
�����\�{yC�?��R����L���]��O�U%�Y����g6�.")�aU���m�^��K��F$�����p���������Mc"<O�ɸ��:{�9�*{��w�b�x��<�)╩�����!���(Og�<���aE��]�0JS����%oF�`��o8(Z|u��#ా��6�R�8�LMM��Y���[�mlX����['UoE�5\��=2�e3e���:1v��c�3:�����ks1IC̠�*�8�ޘP2�g�kФ���M�Ԑ��v�t�tRu8��Nlm�n������F����΢��N4#���B͵��~�!:�����f:h�2Qw��|�'������i9;�h[CI�����q��ӈl��}����M�z���H��*��u����H��brn���;�~�����+�̋(���<��4��Dy�qǎd�
��-�u�z;���'_����i%@I��p����T.E�Y_����#/|�G��+ꎫ�.zډ�N��-�-��'�#N�ǆ����}IWt᣸���*������[3ʃfd���«��iae��
t 9�|�	<���ã[��,<���.�.�5����7;�N�]"����<�N�?��V%:^�U��1a܇>�k�� cBr��3jnH����E(��]<�[�°.�J�o�Nxa�r�V�ت򆠡��߰��u��
x��[=�D�'��GGzt� ��>{���<���O8�-Ğٷ��Ϊ�yK�h�Cj��X��7;/n���(��x;L���  ).�kŬ��%[V7��͢q�@�Ѯ�R.�A���kllM��$>N֗�a�G�'��'�����������Rc�Q��)�; \[�l������zK�4�%>t�l]}U���l����5��b�=���H�t�E qg�Ýu��hc��6>ԏ>JD��o�X����8ʨ4�����[�*�D��\����\�B|ڿ+���)Gue���_��Ǘ��9���(g��d��#QW0E�@�{p���m����.e_�?�Ԯ�<̾׎	>*�c��aqy}��$vi���1
��0���V�ޝ�C��ЙO��s��]���LqIm�dۆ�UD�Tu�po�_��dF݄CY���%��{����������ki����Ķܛ�8���m��{V�3b�u�r�N�������zM��dz��$�͠��%JZ򺤅S�� \�m46lK�]���A���&�%��_\���e#�D�n���F���m�~��P�M�)�b1��������&J_���Dr�->oo1�<#.b�q� ���f�E��b�0e�8�\����;�Q*��%O�v�����aS�"o0D� j$s�/�}}B�����Y�	���_�ћ�Ï������}�D�PȐ�i�m�T}����&%4O�!B@�/�{�%�3�D�����
!��� ��0�xf�����	���J8�<�|����NA�+�ؚ��g����Ͻ�����:6�׀�mu�m�j�#�T���;_9�x�����P�-�jh�!����뒻�X�A����I#CY���]�%�B��1UJ4\Z�c���Ո8��"�$��sgy�_h�4��U�&��ϊ��|�P+�����͇\�F<�ے�?��EN�sQJu�t"d��d`�qsrОk������.}�.&�;�&�(*v;_����n�Ϡ��%!7���*3���F$�	ߏ]���29��?��B7��՟}۵�W>���������:�)��eYdy�'�G��Z�Q·������w���ƴZ])
�oݵ�Q�z�6t��oߘbۑ������O�ֿ$��l�-8�{_eo���vx|�(kM	��'�]�\0�ǍjL$%���]��T�cQ6NF����\+�w�-g�x�_r��`�fG��l��߆n�'dU&�a��ٽZciI�J���Jۂ�Ș>�]�C���t)^��sjs/��"M$�5�(Ux/ɱq\S+XELMP�n�|9m.�\����-�f�+ rw)7�z�;[Dd$tu�T�6�/��Wڇ�(��i0(X��|����/b�a�g�Ӥ�^����U�G���L:z��ç^�>���3k0����
�� ���%��F����!
M�?FЏ���+�/ɫE�ql�<��4�o� :�2n�W��H$\xX>T{���˼ǿ{`�>40����\�fD����HL��<��=�sz(���MK!�s���vaycK�f�.�据�S��
�{����hm��Hܺt��]Ϥɿa��@�(���Ӆf�Z���ǭ2n
j~�;#q�$���D�}<�{g]�"j�r?K�`�x�~8���"�\����
��bL������w�������x�L^l`����nc7��|/����>�\�܌�K/t�W���W2�x����ݬ2%P����1��&�P��˷-�cy���ê��&a��"�lO�Ѯr�m�Ye�-�HTR;̝����0�k��eC�|��҈�q��<��P��p�������a)����=�����\��5gW;��I�x��oPo{�|�U:?��I��=0��}�ECp�b��u�bɀ3�&Y���;��z�������xN���O����OpD<���P�|�9�I3+��4b���j�[��%�8#R��%�  C�,Qn*~�AvMM�RRU���^^2�u�9񎆄�	q��/j�#��EQ�o��:��SA~[��1�Tt\Z8�i�J�Ã�+jjs��Y{��c�W0�r�Z����oN�e�������h��k���/>>K��f!5*��k�`�PI������Ơ���u��C7=]o�O�C�l �B���^���lr�I%N��W,.k��kPRg�
����^O��㝈�3>X���q^�B�Ux�͘����U�>
�����h�k�z�k�Œ���S{q/�,�����a������:�1�AH�b�S���-��W�erNghNWn~ј����;�X�.;�r֐,gIr���O�Z+#`��!Vn�8م�fg2���������%e%���|oƋ;/��R&�X,�=E���r������$��<���s��{�'h�2g}<�����6 $��Oj>���:�������׆[��1�~�� �$��,ʪ���[���<���ݚR��:9�����m�'��r�8Y�HJ�ƾ�\n�q\�8�#k�Qh�֍D�.�BN�rX=E�$~��-]{�L:à8J���Nk�Ew�ID�%�0v��g��;�����J�lw!�M��#��� :�s���E�;�g�mW�5��뭜�|��kG��+s)H�+���<��:����*��p׋ڤ���h���%9�:?6A�Y�|!v��}��v��^=�����7��:@9h�Z#_��<%��Qg%��(�ԭ�*j�sP��o���o.��'8��'̷ߘ��0��e������-����V5���> *166��ge}�#,,�́���<y�9��z>�IȚ�m�9F  �J>_�M�TC�3�+��a�;[H�s@���7��e��T�r�P����/�����rU"�h^� ƭB�ؽ��簀����S�ɝ>w6�0���:�K*\o�e���>����2�	%�G0��ҍ�?t���Q&�N}����1L��Ŧ����T���ᆚ�L>����^?���2��_j��i�߫N>���/�N�x�uv�V�NA�g+��{]��� ����u7��3���t���I��&L���.��������`��/m-�a�%=�큡�8o�뵻�a���㑬�@י��&iiIh�^X���OVso44�%��M��2F^ |zrlp��"=���pJ
v[��N�t�0j��M��f�0����� �W�Ltv[�!���).�ɚ�n�	۴*��[�+"��v�1SI�L��ص�ʯ��&8-�S$���7_�6�t��Ӏ���Wy5^��\�2���*v7�/���?�h8��������byw���I�΂��v�	ֶ|̈́j���MYgb{u����U�~!%)��Y��t�y���� ��5�Ny�'݃qq���z�5P�4�4=�5	 SBئ��/��aEWF�_��i߂2tm���:7�sff�]�,|�����-cšt	X8~�����Cw?���QF8U����L��J��$����O:�-��e��4疤��У(�J���1�df��	�v0N}�,�VWp�|�ݢoi�@�iQ�8]F$��S�b���<����]�����dU)����1|�1ǤJdd�I��aУ�����M"��C��L�V��{�e�D����ƶ�Ł?�D�u# �#�w���Hۦ�û/��$��Ia�h��6}qN���+i���A���� ;=mqQC��+��~�Q.�S:��W���­n���%�1םlp�����C������q���" �齖81���/�(��Ay� �}��w�G�!QQK3��f�bͩo#��;��n�W�5na�<��l�>�{aռ^��8܌�'nXO����cN�/��w� י�h�)hc����$��Q�i�G.�1G�j����KS�]ryE���ۋ��m{h������+Jd���h���C�i}�G�ZR\��+�ܙ�+���r�9���r#0YC!&]��W˰?�K�]L8V#h4Cjˎ78��N���3�7�F��7�&M`�D�3x�&K5����O\�B|ef�|��qS{�5ccIeݙ;o�gbV�o��bŜ�3�!տ٩u�	��P'��y�ߪ���XO��;����
�<���Ӱ@��l��}����ON蠒Y9!"����4���r}���B��{%�<�Dֹ	q�����5�l����m��i�?}b�=u���ϡ16f[�艔7���1ۙ�ƙ�޺3�n�71}c��ڙp��* d3�{A�]N�w$�t��!~���=H�t@ۨx�����`Wr���{��z��8��8]����?����ȷ1s�
��V�VFk�[0<T�0I��*g�z+r2 ��I����%��4#�8N��\R�����K�Z��/D!�;f�$M�\P!!a�ЄT>�Ȃ���{Zg������z�m��ڌOO��-ʓ��*Ch�����=�[��Z�HN�'0�d1?k���F��;ߍ�ݕ�bv��SPF:�af���oYZ!@ȊJ�Y%Fά�v� ͤ�n����x���_< �kĵ�\���/�9V�Ky��o�z�����wOS������o��3�Vi�������'��������G c֬�+�sqW�к�D5��n�e݇��o9�7���\9:�������$���<�Nh��o���C�^���� o�x�݌r�Y���ַ�g��K;���s�,&i��i��L�D��=3�w�F;�ϔ]O[���>�!<f\/��'ػ���o͑tA�-��h�6��x�/[>�wvA}���ge�p'K$T)�C�,>oJY�K#a8g���h���e:o����]�����Ŕ��JT���8����H: �ڞV~ϛ�;p���n x���&G�����������"1}���Nv��Q�����kyt�4S��<c']���5nn�;�W/[df�����3��R��^���+��� �0�	(��E,qR��ٝ�pz�Ү�
pX;l��&�(s SG��� &�=�;��P�9�7�+�8���ªV_�VP0�2}ǙR��8����H����[E\*�l�l���_n�פ�A7%���㫞����g_}�]��1~�����	�� ��}�Xb!�&����NDo�����7��X����;�~��A����"^�mk��e�?�X�碌����98�By�?�b�g��1��s��v�6��a��-^rh ��>!�RF�"@�Tj\���. 6.ކ��S��a���i�@��DV���~��g/��n$��<P��y�q����}p�J�K��u�AE���VX(��"΂~1��1�yf�>HDAx���l�$Df�,*�%*Jk"��e2G���3�	5���1�����*��e�x�=�׻hD�74�ԇ�<�C��2�B�ԋ�@�]�M볁�4�In;q���t[w2 4@�(eF���>=@9^�,_�{��M߃�O���y�Ω2�C��W�s���5��~��
ķ>]�I!��	��a��D��V�t�R]%�Wh�`�'�AkD�l�#c⹻e�\NS��2�+Q�M�
wL�lB�γJX��Һ�[�)�@��R�Z�>�L]�U\F�fF(_��D�m��5�s�:u�qq�)l�5�9AR��#o�A�����tϸ������0�Ah���<̡��T�$B����/�%�煡��������'[ܰL	����	\Jy	��n+Q\�?��g]ol��[�Y)J�\�hF��d���	�g�mD'�G�{xٝ���vN��_J2�����\|0ש��ԓ�w�`ΐ��㞧�%�1�|�jm����@�_Ƹ �[��C$E{�=�57^//�R|6r�a2�ϋ+-
� ��F��	-���i����P�b;/��W��6��㹔#���:Ƀp9 ͒����0Fmf�ώ"􆈐1�̡�[n���e�5Q%��
��9�=x�e�.���IA��Ǳ܆uwK膣Ezd��a�w�l�={��YӍ��>L2�z�xl�|D��i����%,��kv�QG��t���n��J)����`��l�n8e�Ϻk�'|��ځG��|G^[Ա���L���އ��x���m4��(r�xU$��O��A���8'�ثD����k��?@҂Y_h<�!4�Ɨ]�/V�+g���>�4J���J�}�x�VPF8c���±zA��̋M��g�|d��d����~FiL��cA�j��%�@>c:�+��Fk�0{�,.�ֶi^� �(y����>p�sSx�=;;���yѿ3[+X�qo�Hql^�[o�gvGN�uM�/��f}���Is��F�*-S˟F�}�H�k{�}a��`"�d��OT����3��A�hy	O�;g��ZlS@�D��Q���;%bo�6ƞ��hg#E�U_��F�A�tH7�)
H)�).H��(]��t�t#���� -Ͳ�t.������;�2���>���|��y^N�:>�?�+�mi�|��eA>TߠT��~0??�̟�o�~�	��~�>�������d�;]���W=���w����Vɳ�zKs�_�F�,~"`S��u�kRA����4�5>���%	��_���~b9�+0_u4�:8�h!w\������c�졏��'�e]L?K\��5���vN[<�u��H���ʍ���{�gU�L���b�PD�#V�	�9j1�F�|���qv̛���u˪��Of��fQ-Q3�)����QJ�T�5�t�lR�]D�`qÝ_�Vۗ�O���,n��X4���u���	h���O&	:e����JZ�$al�}g�H�#iQ��@��3I�����F���&�7�lFq�	g�5j�Ky��1�&�z"����
Oz��^(x8�%� ����+�M���%lm�}��N��w�ҍtw����r�C�/�q��̖��Gs���`G�k�u�!)�V�z4�����j�%��+�д��f��/���j��K��w�����nj�l���ߴ�����+�W�x���2/�p�r|�=a�b��'��g�����*������d����o*�d���x����f�ec�
`0F@���]�_cZ�i����=<���$�	��>l+}����7}�u�퓍�U��(�.�OO؞����0ER/�`�0^G��,���Oz=!o�X1��r�z�g	��ڊ\�����*k��K/K���/�g8�����{�./O��O��`n�&M�ۃ�+W��ʬI����B�0� n��+�
ד�F���ʌ	*�~��3O�/�G�J	�1X�-�����A��nͼc�zXF�i�7�C2�/e�6���N���#�6ǸfS&�_9K2*���9��PU� ����pA	��oO��
�6wB7��xK���3�TjĊ#��0y�H#*�[����.�V��v]�x�>r�Ű�w,L%���G������*wh�QĜ��i`vl�ߛg�k$�=	o{�֝��eo&=�.�g&�Ұ�l�lﷵ(/���4��+O�0l�Rݥ��`��$S�V�<�LtҁtWJ!�f�9�o�������bf�u�&��kjK뉢�̡L/Z���0;��L��������+שmwZ�2���4xl�;)�8{e�'j ��ۣ�M���:=�.T�Ѐ��H��0�.��������1ܗ�L��ó�?�/�F;׍��J�iᗕ͠�M�
��-��J��	 � ��1J����ܢ��NJ%Ծ��4M��`!�>�>⨞u~қ�)��S���V@tt����:��'%%7촋F׷�F���}Q~@W��٠�lXǏ�A�Ȝ��j.�Q�'��y�����'%%a`t)���	RNz�1���?n�>��*v��b>��� �/��1������K���l���p}���r�MҪ��؛�-{�9�R��S��﬎��Xzׯ_�5]rH$r\��֜Q���v"--��2�Z���}P+n�&�=�U�bV�}ʫ��yN�7��zh3�O
�Z.�:��̗�Gmٔ=�D��o\c����3�4���18��;����o��?�`��>�>���B�s�(�]����ǃHܦN]$��R���	�!Ѓ�RD�G�/q5k��z�$�L��zj�3�5�t�%**ՠ�}�ֱ��8"˞�c�Joo���`8]r�E�� �v�e,t3B�sn���\Џfu��ҨX��9�0��>=q�Oc��7��/�(��j?r�������I`� 3L
��Sϱzܵ�>n�
 ���'ω~h�9K����$��yм���U�e^s	����,�b��u�+�G�Rn�<A�m+�F�V�3R2�9D�:��̇�������桁�\�G=#��R^jglKn���w`խ���+����w�^[y|�(�SU����������6�����+���er����7�.�&�m4�wu�5M�^� v�I�((��}�ޣ\���=n�)���-�L#�h�dۋG?\����4�4O������
�	�*s|Q����9��J��~:��^��ߟ�Z���$G�G��]��Z�.3�E�_`����O���,�PN$=��,��4P��y��u�K�~�;(�|m2��|!qT�!_	�gy{7�� �^:�1{`�J7!:��'��\T�zA��İ�����/�N��*�j!�&��xG栗RP��=�=#�aΣ�W	J�۫NT���Y�z���hr'/It�J���T�{����u��@j|�;��N��b��S��?�ң�?8��f0g��t���%�d�s�$*����ћU���B���٭��?����5���uӼ��ʀ��r���W�Ύ#9&��ݗ��]�ß(Te���^���qG�E`T�Ys�Ik�Pgp���B�L�rt`z�g�h༖������ך����3Skf�ד+�g�M:rHZ���l��'sxyw�5��< �d�&br��/���x�߈S��Ⱥ��Q�g����JK��CV�V��)��e�u*�҅�02�a�[0����c�n��hz�|(��@�9�/��^X0=��%���x������.a����m��UQ��&0��?�[�yy��� ����	fMϵ�ټ��<ݩ����]8�Z����������fD#���I؁�ɺ���8+nӆ7�X����α z����D��yL����L���ͪ��S���� ��������(2NAQ��#_,���Z1=e%��;�QPS�ۯo�@֤^���Sֆ�&l�(�+�O����hf�W1t�J�������SW��-�]����_4Н�a������"��/�;;Y�C��4��0CTf�-���-%��L����ϊ�`�.���I���G򀿖N�>V��gK&����4mx�x�j���.��5p�J�^�)帯�A�1Pm�?�	��QjP�֫���ο1�4x���|�?�d��&�V��cA�M�IR������)����f��ͫWM.	/)�<znӭH�uuuj��[x�����OA�WC���˽_ ���lf�bIX<�_~��
��������t�)�b�T7��ñG>�{~s7}�1��b����W(�+˿["8Iq��h���	j����n�����@M�/��c��9�*"}�/��jS~P�8�{���r��o��
�K��^���ٞv�K�Z�׎���(�����	$�ڟ��6�_$������	8��TZ�d��z,6Y蘿��	�#������kX�BЗ@��g����=_�0˩�p�KJB"y�/����D| �f���u�sj���t��s)�7��U(:�֪֡f��ww���M��l��?���U�>��R=�~x�zG��W��~�d�e�ե���s���6���y��p���d\=QB�_B�d#�L��3��]2m&�i;~��2Iqѭ˴�D$$p�����i�&UC3���.6��Z�!�હ���+�v~�X��o���O�N �P��K����$��&S�ne��25/�v�$�q��az��ʾ�d8eU /�iT<��bmt�%H�M�����Ә�p%oP���k�|�8���m����qS�4H��^��bLb�2��Tط�nX����?�u���z\�Pe��U�<�Ү}��DZ���C?v�*!��4̢t~j���E��O�?���2tG�F?f�T�avW&��\%��B6q_W�L_���B�ޢ���ۈo�vj��X���2
�u�x��g��ҵ�ǷL�C�sS������q����8��|	.�mX���}�D�u��Y���mʃ�K��[2�d��>���;z�J�����?7;�%�htf��y�j%����=Ce����E�0ڳ�clek|��J��b#�m��ҹ�����A��]��C�[��sD7��j��;�)H��^oMb�����Z��w�U�x��Ȅ�fP@`1;�L}��mp7�A�����:Qx�9~��i�8tvLH�˔���t�P�� ��)���Y�㍝�S��ț�N"Moӛw���ulm�"��>k�x��AgOlpr����I�;��u}�w!\*c���.�(~SV)1�����������t�O�V�a���`��8�����,9�+����z����sA"}K�n<pd}?���Rz��!�&�t���b������So�ĢP~���ë>$c��M[�R����=���k��'���G�`�bg�����\i����B���Dڂyn�R��2K�Ϗ��Vwn�����2b�a+�`uˮ�o�$H��������ӾR�ܱ�D���$��%��G<�R�fj-���X�-�RJm�H��{��8��XI�$qj)9�A�/�~+�(y\2Be��=��@�5O��J���/�9$wq`�{�-����^���0�vzv6�{{��+�I�[�rE	�y�s�Z�G7�z�$�[CXgwQ)��C�b���B�����P�u�%Fq�Ge����)��usV|�eCRB-n
Ov�ަ#���y'O�}��	]v����%a;CD>�S��[��3�RN�!	$�:����XR5�\vI\�t�/��*��A]��<��}��Ŭݞe@���_Cg��l����]m���Z��YA2�9:hZ�$g��R�47��5��(.�@�XtJ
~��m.���s龺ݹ��$5���\J�1�Ҽ#`����n�K�V�Mq"�X<�V�9�8��n��/D��6r?��J��gV8޶�V�T�z������"[lf,�'G�����U�����Խ%jo0k��@��hM�"��Na3��s�o�x����a���1�&�vv.05;{�	o��q�r���Xս�7aByF�\�W/�Z��vv�|�C�(K��ڸGts����Z����0�c����as�}]0g����	�{�@��KM��l���lr�1rx����6��e�r�JL.Ԯ!�PBϩUpxTi�?����_�*B1��_"^���~�2��fO� ��h�~�.�����8�쵺=���V�K�6Oe�%�e���(I�#���t�t�!)��"@W��oN�6��Do�/��J��o�B�,��W��gBKʘ2�Y��<O���/�̓�����Ѭ��� �_[�k|ef��;�o� E��]o��2r���^����y�߁z����kh�~W�}�LwG�݋ɞ�M����^D�9�M����k�_����~Ҏ#+w6�(1ѿ�]����+��d���Q��L�X<��Um�/
w[4(��CR�t�@L���f�.|o��VO�A�6K�IG%\���Df������ck��)_*����4�{���k?���j��NrЏC�%�o:��(�xH}��fX�:��I]�Z���sN޾�:�����������o�LDtW���r���;e控\�wk��X���l���w��l�����$-����v�;�J�BW��!4���H�S5��s~/���vg-(�^eċF@I�6�NfȞ�l�>�>�kd��9����z)�������JEOO�{C�y��ig�6¼���rglt�I�ުZ��n]E:\�3�<�j���6�s��W���I��M�qK�"����e90����W����c\LD��g}���H��=�`O���o����)f���96v�S�ۅ��%�>$��-~�?-5��1��E�$��ޡ�&�8��9���ou2<��U�lݔiH�����cz�=	�K���c���'��d'E�F+�WM7�0*iկt�I�[T3C*��~�	p1���s��v'�_�|�u�:�Y���u�B��T��T�k}���Q�O��:s�����
r��w��)�wf"�^E!�C|�&��B�J� .��.�}\X���tB1�៙��f��W�L��U���*wPki=*�3���q�i��)�rN`m"��3�$^3��X�d�����o��n���<�����x��,h>t���� MT`�W���0%gp|���Ԓ!F��}�ao� Z�^!�Zx�p��-�fM�U�E#(�����˦`����&)��沌�K4�h�,{~d�ϫGߍ������K�m�^NVA3>����D-����Sծ����'y���������([��88h3�h��`@lH�o�k�P�шG�@U�y���k2���U�D �lȓл3��,�!���������ZR�E�-z1�_NT��؎��De���,5�$�����z:�g�z8����į����G��j�'�tuu#�8B��p4G�f1m��ނb5oW���s:Sc�Fm�|�D��эT��^N�Laʣ��H�x��є7�u>eh`�j4� !T񋋨ܢ��%�������C_���)���jC�+�J��z��bk���H$>�wû�➸,Z�x���K.�lV��D�� j���W�BE�6~�e���Ncͧ���Ks8xj"�KՈ�w52�
x�&6���yl�P���ow^�I%X�#�h��ݨ��W�B?�͘m���pOPH��+6�����L�7��[n�Td��)��C�௦���3:���/}�Ĥ�^��!���,7�譀�E�e�#g�̯I���.���S��6���5�c�<K$��0mI9#u�����?C�ȶ�٣�B� �m�����\���Ob�wIȊ���L��+(�dw߱���1���ߝ������0�r�n/{N`��s��r�~afV!E|%0P�L���+�o+$���I}4�mv��9\�J5~jB�vk��q��;�?X���ᩒ9/�ð~H�7�((�6�6w�����W�'�s��	���Iț�?�7�B�T��8���o	}7yҏ�_�qR3 ފ��poC����sΤ1��E�x���8%d��T�Q�[B߈��tW��8e���	]����iS�I�� �Sv��U�Y�$��5��0?T�
I����^��UA��^B���K��׸��R��c��K46��Kw��4��`�+�
��'����튍�8���t��N�4Se{�0���&�^����8�ק\��EBe��0�����,��!����
Ǝ��\B!���&�!�X�4�zw���>�|��3ڬJ��H�-s���g�/���=��}Z1������|Qbb�]�k����ڡ��|���N#��+wr?�
�i�����`��$x@��!�mEg���1�,Q��f�1�dswY��.�an�'\�;b�,Sh�dG5FPL��v���0 ��H	WVV�Z���[5�p�L,L���Q\�'=YIH�����wk�kD�n�<����L�j���C�.ںl���ġ�UvP�Xp�s ˩���qB?��� Ōf���`����6��^S�oꪒ������h�P�\�鿼���;���f��
�s�����}���y�PyѪ�.y�������N�i�+�Mxk��w�<߯j3C<]<��O�p� ���A=��<��ތ12�(���W!����h<d��Ӽ��.�̭�g�?�Hgc҂�ؙ����d垝��K�sʬ����)�rf6!M?/��3|�g�w<쩤�"1Y�̨�!�������@P�ʱ�$��}das�2���Wפ�w�M?E˿ҿ�a:�4�ů�/��L,�����G+�-7�@/�~2�ؒS>�Ǧ������;c�=��Lݓ�. ��"�ܦh�J�A�d}-͔�ʔ�k�yF_�l��DRٺ�G�3������1#vc�� �8��^�6=��8m�.A
�4oY9-����q�_���l~��:���k�� �1�_i�|�/.���"��Ռ�?�c�}���p������_O�x����!�6K��5wqQ�5��<���/)���2$%L+��������ء���L���RM�޸��g)����?>zA����������r��m��KL�c�&<��s)`݆���.��r���6mI	5i�D��4�_���o��x	�bO��ʯ�av��T �	?`�c�?�$K����KD�ۇ�a=���yRm9�7�i,���n��oO7�j��Y-gH�o)K��D&�q����#P�f�?��L���Q����C���}�7��$\��ր�ш���S���,���J��oʸ$�g3�ŏeԌ���}��Ny�����/h�HiU]ޥ�W�Na���`պ��o�3�2���]l�/�6"���V��D����o��z�����Ï'��<�)4l�
n��{H���Ҳ�+nm�^I�?����<>R���}N �
xǧ]e{'в�U�z��ן)M���+kt*�
#�5����� I# *��:�L�m��#��(����)jH��z܆R12�D�-��y Udx�cI�� ���6ZA7�s��\����/�!�p�=Mf+�9h0[2��-��u8�y �AbT>G����Fx!(㾡ߠ�`#`��[�)1�p���̦���-o�ct§`O��YT`��GTM��C棞|�򋷵�0pQ*`t&�65�T�w��I����9��B�����I
=U�;6x3O)�v�����cD&���כ�ұ���5���r�z��l7��s/3�r�J��0�<������������"TC�"'�p6�f����(z�q��m�N�;�-���/�a��W�����I��t�pf�HQh'��*�2��%���"f���;���������q��J�	`,WJG#����RO"s4���"�/H��Yl���8�������("�KbY�{�ۛi����a�����]�|ӆ���ndd��~'�!��D�ˌU[��ޔ�8���8��Z64d]���fH��S�D�����J1P$�`u��5��H ��F" RS9���IQ��.�Q�砬�2�:B��-�ȃ�s���ܾ�K���T��x���+Aw6᲍ݭΘ�!@Ʒ����"Z�}�rM�@�]Z��Y2h���٩A���O<���!�S�d�Ƕ4y��##8g���<j~�f7S������C���5X�Ϟ�Ȳ�ʝ�g ��&w�����N�5�X���lܯv��X0��M��-9�}yԫ���&ɦ���T&Џ���x�î6�	��hۼz��\��T�#"�xҭK���M�gI��p�Ͽ��9��Q++��B!�"��M���|�b��h�*O�J��f��ު}}u��Y�@�M�!##P��]�b@�um���O���DT�FKG��*�VH��|�L�=�نm),:�5l�E.�L�7!��v�������vM�ߩ�c�S@ޜ���-,:�MQ"B$���@�jo����DG� C}��Ϟ=s��.Y�t�ś��ݑ���e��;�O�x~���K��y�x��~"�30�k�e�[�$���(�_�--M*�pH�����e烏7 6�����,v9G\�{H
tJJ�D`�"�W�ؙ����Եy$�;�&=���B���A1���CNa[��"�s��u��}l��2�,�C߻<ȁ�����|�s�>���B�_Bߛ��W�BNr{��Kn��v�zV��`�@�$Ӟ|���90�j�&��F9x�[�D
'I�S��|RS~��N�;p�>kǳ���fj�����lѧy��vl���
��q�G��|m����ǂ��̬%�t0o���۸P�<������p���MyQ�p�^��V��M����pKy��'M1��A��������صq�٘���Om�ޚ���?��b%K��ӆ�U+�d��O���Y������Ŧb3D��L�����FT�3W)���̮o<��c�
���|�K�lh�`����FF���|��26��L˛���'�$P���CRrZ���5�<$��l����^
� >j������
�@FMV�������f##����oU}�?c��˪w��о�A�s鐮4�����BI����F@+��T�z	1Q�>�U��o���z֒����Q߬�iC6�m��(NvT�� ��U����ɴ9�����H�k��W�I��^���8,��m��}X0��F�MNB� &=-�����d�󬏪�yϛ�5����������
NQg��ɰja�`���:��f��,f�̀!�Q�-�q)�'fJ�4o��	�-[���Yb�O �T}o/ i���Ч2���ÞH ��^�o�f5��� ^B̩dҧ�w�^Ǯ��������
��`���!B_B����.x?_��Ĺ��_�'i�_�����Ʃ
v?��]����������q�o3|H��P��2$�|��[kl�iQ9�,�������&J�@U��w̌�Nn��un�-����[<�����x��^'8�����I6��"��V������`6$��0�������G����U��3Q��x&�}B����ǂ�� JbXV=)�i�/F�[��8��7#�cF[e�==@iՁ����u�/z��M�6�PH C�C��p��~{�g�n�`C*�s���$5����͕�`��T�M�wm��Kv���)B��٦ |�$ގŮ�"�S��N&[�:�?_驺g���H��
rssf�YL�ͧhYA&{��+aǊ7�������e��-? ���M!����"�r{f��A�������r�	�"���6CZW�o�7f�!�Owf�)/hz�gQ(�r��{;	@����}Q��8�)-+C �5�*��z��iK E~>(8R�r��3�'����|��M�6�T@���1m2���R��.Z^"*����N��IT���y
*e�\����K2�u������/�4�*�����j|�}M��n��6��Y1T
ȯFR��	~y�a�x+��裢/��biUl?�E��������)�uo[�����Gm"�˟M��O,VV��;z�؏�b?���&�l��^�'
�'{\>�6�f�H8��&�}������F$-�,�	ȏ�����]�S��;�Q�,�.����� bLj�&�۽���L���1"���T���2��0���.���TS���s
��;8���sC��4G]���L�[����ҭ%?�խ�ݩ�h`(
��w>�f��	��TÓ��[ǭ���'{��8��dP�55��C���<���� ����U�Rs¬�ͻ��/FEBI�r�_����P�~�H[#�*&�y��^�{H��6 ~{�{�%�s:V
xN.���߭�X-g�醍N��iܪ�g�T㕁�;��h��xG ��[�UW.}H���߁ر�IϳۢӾ�������ls���V������"�Ņ;&�+OƏZ�o�I/��<�ř��G�r�j)�S�GP~��d��~f֋߂�~c� x|~yy?=�ݭ���-,(�����	�3�2���KVD���.J�����Ӓ����V�l�;�H��1�Y"
+��Yj��OX���uu�B���b�t�����!ֿ[/��Ҟղ=�'�3�>9�0�$�pf�P~_u�T�����񛚇c�N����9��<mQ}��1E�&�V���uboM��gk�-*kg����MQ�� x\sPfq%��ۦg�,L`f�V$g�&�ܴ$��cg�KcQ辪ݒ�C�����}��<�0M�@����v�F�-W&��sc�A�M�����vo���4�@�S"���ʝ�����۟Ar k�2�`?%��.����Y\f�mDLazd~�َ�w��hF���F<�]�)�O͡������Q�Qp�Ic��wnY�w�W#���gC~ȟb$������4݄�0=T2��f��:gb]�h���_h�/yJx�1}�ʹV�(\��7i׾���ѥ����/-/))iW1[*)�4:���Sĵ��ig���N⓸����������}��G&"�+s(Sq��:���`�����]5q,֥���B�i+ݟ�~���)�߮�M"�koW�t��dsT�KF �	�lc���w�"A�����ˏ1��}�Ɇ��z�-��h�!�Ϗ�"���y����A��H�ڏ&gC������F�v�n/�5��W�69.�ǯ�oQY�.B�[q\?�P+d6�)굿����-�;���v��bs1���'X��-�<�,v�������)�g�Y�H�Q����4�B����蝧���6=��O���}��?�O~�a2�WPX&��'C^�S�b����VU�ʏ�+�"yg������2�K�Yg�z
:aP�"����_m?ا2b�r�'(�R���*�f�r'�f>[HPP�X�Ր�����qR�������r��J�Np  �O�#�B2�AQC�S�����P�ϖ[��s��URҜ&x>���}b�gsl�'r�7�y�Ec�IM4*wt����p���kE�G����"y��\B۹60?XK'��t�H�����ة��B,"���	�^�dcB۴U�Gh�+Iw����,������g���l4���a���MQU��-���Q��f�_�~�)�0�䵴�]<؆�g�ZRߎPK��Þf�4u ���Y�\z t��(�g����c	�91e;�x8j����ڭ���.?`[\�(=J��rRy ��q�^j��F*Δ�@J$��rՙ�+�
�Z��ׂ(ORH���-q��+��w:�l�D���D�~���층���0�`]�J�i�VG6�Y�Q�}#[ku��FR���wT|yy�e���A���=>��=tc���[-����~����˦�"5�����G����T��)ξ~~�W�*�ff����aJ+6�����:%�:%_?��z����=oiKPT�M�����o��XN�˓�A5<�u�Jj����E���,''7���}��}f!y��Ԟ���K�'�O23��1��?\�/���Zj��kp�ڥ�b��r�PJ/���p���ۗ,����#	=�f��d����^���!�����-S��j���O�@����>����s9��%�kF֚�f�L����[�d�PlE(���v=t���B� �����i{��s�0�zEG<郮V�Ov�#�Z�6%�פ�7Cm���1��
�ϩ�?0��/3��T�n��=U��>y'-d׼Y�*Ruj*�A������cM�����b�WɈ�( �$T56q��&'�/d���c
W�uzcO��Ч�K���Upb�ׯL�ϹȠw,,���\�5֐Xܠh�&Ƨg�В#�77�D&�9����_ۯ�
���1�{^���e�T�B�o,C���빼�#]Mc����D��"EϮ�~�6�vXPN��
� �����OGp<�����*X���(�r�\��,��¨�s_�����R����k땯���ŗ�KKK�����U��V�����C�M�66�w�?�u���z<�e�{�-b�w��G�uuq����匎��g+Lͼg7��I���A�%�1��	b����2q^n���T.��R3���K�-ǎ�����L]ZZ��:��?���=$@s��!�pe��kcG�]D?���1���6��9�˝��������I����ЫgILc�h=�A�>����1n� ���h˵g_qZf���/��F<��M�>*Z��eq�3)`ڝ�M�@���ƹ����:���;��|?���[R��Å�e�����,x-N���'��k��Q�M;�i�gҧ�>a�HABB�����]�Ԕ�뗠�guC)J�;?�X	G���/ܜ�<��d�+��:Y�R�z�6����p��������4E:%\��x��  f��s�gk��;z� C�*#.��/�]Er1kBi��!�o�&��[���ʅ�I�k�Z�x�̃a~��	���a�2�d�,�Mj�b7�����d�@��O	�����e �F"���V1\��=N��o�bz�E�/�J��{��D$ͧ;ס�/�Q*ϞˋF:î�n�.�b��c���*�������/΋�D�T�%.�uי�[^� \�w�4�q�+/�i���`f��/�49��Na�D�!5��b�&<���,�mHe~m)̀��ڿ�½3����'�wƖe {e˅��ݹ�G�FMԀ�{�7��	ikV��*G���j���b���SE8��e�>�A�uK��5�4Z>m{HϠ ��4�Wċ�5����	9�J�`+�����P��B=�0867���N�[�P�^�
vo��3f�L�5]%i��)���m>^HT4��p����47w��@��C5^?P�^��ş㶢:|c�3�O'M²[?-���g��o}}}	ZE��9��NP�dSII	�Q:�ysl�p�h�H����$����BM05(J�FT�319L�"��Q��>^U:���	N֐q�0e��ƚ�6�E��K/�:�a�xF��@R���3̝��a�X���H��'����L�s�=��⦸IE51)�.��p���ƷC����<��q�E+�eJ+���p�}y i��=�M�.��uN�3�9�r9?�?��rT��SЩU�"Z頳(;�F�*\�j��<߸�=���q�|w~�G~s��8��5ݿs��1Y��㞄dǑ]�6i8M�E�?��2��ňw��v�4�9�S�9�>���)H j+�"�GMO��Y�0�`�h����~�^;ȏ�ZWz��M�Ǿ�Lj�^��(뾤��Ѭ��*G��	�L����m��#t������+Td���Y�Y8�8V��ER�`lQI�4�g�7��!6C�f�o�j@�Xח���
���W��b��XϓO�`G0�b�t�a��e�.DMٳAĜr�+++�'�8�
����O�%�h N�:�F�?IO�%OP�b��j�
ʪ�x?;*���I�j��� ��W�D2���Kdzy4���!�)��IŬq���1�r���� kq���,f�љp���u{۟)Y>����oB����{B��^��[ �A�w��v==�o���ill��*���H-�W�@���8[� �]���F&�r������#�2�+<�S��_�4�Fv���4`�6�t
�j!��9���#�{��_��+a��.��X.�~ᴸ*�������3ҩ�e�pi��=�,�x��B��ژA�ej��2N�_i�(��R��M��1P��㸉��r�=�r��� ���ݮgn�M�YJY�6*d�mK��[��'���;Y��4?�����<��LK:�s@g��il('?�*.¦���6���7kw�BJ��Y�����݆͔gw44�M�0�&R?55�>���p��6�dQP=��e�g��%�&E&7WCX__���O�%UU��L�΍/�FZ�*���?�����W�@�g��t0�ǭϷG�x"��l��.+ߘ��G�ES��(�;ȝ^<����LO���'*�~�Y[����%x<kb���ic�՗��c�fy:dmL�.��)��x�b͕�߿���o��:~�B�z��3��%�_0�'(D��)�
6b<u�Zm�)��,ە��nk[/�9�c�[4��E��i��JOX������s���5���ڤ�4�Q��� � |X\�no!1�s^�C�w���'-�C��k�>�l������pձ��m��R��~b`<����Xud͵��W�i0���L��5Ng����5�E=?�h�V�5�ޱC��W/�,�~7��$�U~\ss>��$QO�|1*�x��2�JD�J2����]�XW���}�͔�'dz���Q��g�Ⓠ���]�fл+JyK���N�&�c�b{?s��\L����w�s�^H��I���p�T��������V�~(��խM���s�4����m�`�y-���P������^#�[/��m �%矁�=2l�lp���'-y�x���w���]/�Fm��w�% ,N�;�Ⱥ�ե�'>����>�=�z���߶�xk]������s�����(K#�H�Ji/uj&u��]�P�dEW0&�ߙ��B�pz'��|7���?��U%Z!:��Ѭ*q�:ؽ/J03�_"��
Z��Y�2��<iA��)&��ڛ��iO����o�,R�q�t�cv"X'��ɴP�py�����I{��g5U/�elT�2<�b2��������0��ppC���v�t4+«���LsG�FU�.�A��q��*kj>���M����3 �F��#ej/TU�[=���z��e�N%���G������RS�DZ g�7a��{!|��p�R�޺�	� ƽi����1���}{[��&�$���pJ��B���C2FG�M�F\��.<��6�rlR�P����\ �����6-�~��VQ�'��O��&�0�,R��Y$�.� ��Q�����	|Y�Ђ5/�x�YB#,���q�MD��Gإ5�t�+}���P���i�������ƕ�uz ��q)
�o{���5�c��qf�n�TgQ�4k+� ��׍��Я"�w�ъ�[�iŤmt��ۅ��B����	tQ�y��!��g� N�U��EY׈� 4qȩ�_�Q��;�ׯ��y���'��ǫ�X�Ť�]�p�;��K&I�;N��ޮ��ωK��o߅�H̶�9��ɛ�F���D�oW]^�O��TEj��,C�?	֌��z�t{��F^6@u��b�jH�H�-���~�pK
����
=6&r{,&�i�X��tꦌ��5l[�,�U�9������v�, �l��K�B;ś1�u�l���MgVzU��W�"x�o����Svе��,�����ͽ�{��&p����2U�C���XO��A�������چQBR��Q��NA�Aah��SJ�N钆A:��.)��n���������pf]�>c���M�5�*Ua�~�p��2#�wJ6��1��,:1�$����
����j�i�}ϣ�A{�n8!��x�J�ۿC���)�CTXXX�v(QktD����腩l~�}�����d�d�Q�:���U
��?���\��e��74��kqc���DFm��a�~��A��",�
P�b�p����/,��k
��\��ٮ- ˲��|�.���2��sV9��|�(�Ӌz�nd�Z�ۤO�c#}/��'���^������f"m���hd��V��s C�}C���sD��)�$<�=�>l�7��(�1~�8~�ȝ��\���ƀˠ�ͫ?q������S�z� tt�!B��2���&Y��Z�������z������G�#F�E,�3n�xe)�w�Yۄ �)��]�B
(LC�����L����I��e��F�+�'�xiv����OmZ��C]����`�v�G�\_v��a�y)��{~O��H�	F^��KS���/]G�l3ª M��%�^���ῥ�n_�Ev���pw�?T���N1�2HǨWR�gv��z�A2��W�bM�$j�~����n��n>�b]�`�a@~��`o���l^ e|a�?D ��Y��1�`��N�8�n� �o��/1v>�Q��.� �>�_�?D�rQ��H;�cK���i*x��G�C�O��7$����j�����6
��(?��\ ���bo�&+"� lD�G��\���֣f��;Q�N��v+H��ijc���$��K��S<;D�>V�����R^�Ƥ ���5��(�p	�����(��ܕS����,6}k������?1%�9��j:�t`2��h���!×��:vuۚ�E��Nc^#q��P����Q#����;��B�_}cn.B��V}��A�
�%�77�l��Ǒ��|��.߾���"����������>-�ã:}�#��x����HrWG�B322�N@	�^�H�\.9��\I�^%~	�0-T�(l����d����8�?�KlőD���[��d��ϼ� ��������Y]�}6���O���D��u3i�`_�j�vM�?)�HHͣ5ƿ�,+32(���3p_��ӊ��V�O�%�+����ܡ������ I^	�(@+�%�;K�K#~�}����9Gʧ\�b5������-eaX��^J�wP���9�鮀=ےW����S��~q�/���킼�CAV�^w$����Mwg\�:��g����'�i�]}��#?m�s��']�N^:Bۘ�5.�w=�7�� U��X�������"|�QbW�.�׼���wp��4<<�1����I���&�
?7�"����U"�U�t��́�p|bj:T��A<)Sx�Y��c/�4��Y�.]屫Ӹ㵐��G�X�s�]5��'�`����wz��},��n�|)#D#��J�%�ġ�X���������>R�W�N�Y^!ۭ�U�b�z��H*��s}�O��i��[^����k����s2r����p���*U6d�����g��ݎ�_�W;6̴,�J��h�zNj��y���&>����`�u���!wiZ����f�߳1�i��اy�\��4����))K�����:	�K���kR.�@�>�����js���K>����x�JD�"���R�����M"����!u!�����^� #�����l��2���Kp�Q��mX��;)��xn{:�����Z�%W�B�	<�����}��?�1<O뚂�bk�&p�@���/��eCJ#�]*��<�A��p�P���Р�!��ɰŕY��M*K0�W"��7#c2:�l��ڬ�6�}C�OX���^�.'��ه\��5:��CbJ9)L*|}}b��h�C���j�N�R,����y�^���e��ʆ�c��k�9�X	 M|g��
nu���y�����A�?l�Q�^��\Y2u������=6��ʑXܑE������vw}3[G���U���\�ZR\�9�j��Ď��_����`v�do�h�NV��:P\\R�Yri��~�V8,�Xh�7H�T/�w���د��(l)a�h�Q�s!:k�-�fe�A��yV��
�B�))����9� s���H&Qթ��3M��g�B��/�R���Xt������!�j�d"��	�N2S|b{<����&{c\j*3���ij8@���	�A��TP��r��$���Ez7w�N��+�6�9+�TP�7`�x���ޅ�U�#uvv6�R��U�^���ڲ�aV���q�������O�L�
����&����Y��;dz�����O�(&��Imgn��Nt�C	q;Ġ���xmt;70�ۖ�D|�)�|�d+�;��c�75mk����[[X	���с<in|!S�k��;{�}�|k��h�aq��\�PrU����Q#BG3��3Mʞ�"2p�J�j��L�%OS�uJ�c����vb�E}8�:����4G��22н�I8i7���R�57GS-V퇅�C5����+�Lcޝ1���jG������海Eb�^���|��(�*�Qu��E?+c���y�u>Ͱ���ߐ�ޒv��sVF��E);�v��*���.���p>H^7l����t/+!zD�G�l}���Q�2>
��a�cz�oKf�-���N޶��׽j���.��z�����a����m�or�\��LyB�VP!��ۿnF%Ir�/�����;���C2%.���\s�ejCq�޳9�j�3����-��B8;`y/�>��6�M�T���������蠹{I�+}����J�CԊd::�KS�,r�WQm��lgY�k�;h(7\�}�ޏ*�3j�M���8�8���$�i���,:j��Y;<j�2K�KB�"?8��xHR.�,�(���yO,�h�+�����g=}*E��\�rA �	���_j/�Ş����QS�j�5b�]���4��/}7��>V�p_s��D���2��4�@}!I|� �Q#ǱUR��_]g��=�E�&.�v��$�=�׷�������.�il|e��y	�b.����u�D�N��9��x�6vϯ�4���rrr�RR��N��c��T༛@>��0?S�>܈'�)���p���V��̜5���:��켏K��
�"mU�Ǒs�avz��f���=��=?�낣W���6$�E�孛ە�K�ҳ&�N��z�\�&�.�:���}��T��)��-�iN����#�|A����k�N+Z��3���ǰ���;.S���G�8��$����q�6<��L�[����p�t2�>��|rQQ�S77�)g����T��c����4K�ٔP�	4��4L�as�+#�@�К���r+����7�D| 5����6]�r�SZ��)�M�l<=u���68��6ihZ���[�:x�O��ZB.a>�Ɍ!x�ū�UF�?�Wχ+Y�z|q'.�u<(z�्MJJ*�v)�n[辤�xȬVX002��ly5�w�u �,j���'ʴ��I���� ��_<��^��&�sY8&�K6�S
����ċ���l��I8m-�$*�n�!�@��-���
L�����"�_�fM������P���.�/��D�AP�E8�);e���!D��5�9�n����7�Qÿ��F��8A��\w��k��Ri��#����Ś��)[�B�T+Q\&Sab+壼��e��ι�n���w�B���v��s�ۿv+}����?Џ@,�WF��}3�b<��ϛlq����6��8��g�$��Qj�h2r��Q�Y�P!�BXճ" j%�XG��8*�� r�̂[���j8����}��W��P�{�P��ޖ2`�A�7��L<�o���I�,��w�aN7a�v�7�˝=g���(Uݶ�����y=ޤ�7h(y�MF�$�Fx�Q7�z0q�Cq$��5�w�&��4<�J������]�b��3�#�]i�ۡ���Ն�G�/`������(��3Ieī���<���^��q��h�\ӭ��/���+����_{}��2��)��}C��E��ݍ��0_Z�a�4��y�\Y�X����L�N�UTT����V�'rx�Ƽ�O��!u�	�<�
B%Ǘ���>�kǒzt�� ʧ��IbX;`NZ �ą��MɅ{����2-�GU��g>��ʒ#�(�]Y}�.����L�%$sPS
�|p�ԐD� �M�e���/���ĂJⳀ;S'�>�9�� �P��}���ǵsm� 'ܕ/�+%��3�+۔41jy�O-�7$e�N����y���%�E�S�g���C�	�����@3tA�}��͍6͞�|����A�~$F���(:T�d�e�L|��M����	m��i�^��?��ݹSGQ�!S��g3�:������X���.hO�o�p�[c1سu����WL\�8Yʢ���b�?�	ND�Ql>�:jX��
q��?���%����#�W)���W^�i�w�P�WZ
�d�5���J|�ŭ�QB�� .~8	���A���6��D�M�Zc�ޔ�Lx�vґ�6S�&�_0F�+1d4�q����,�	u�P��}��� ��5-M�6m�7Lk��1%,b�w�'���3���zF�^��L���&V?��ץ�ｦ����=4��m��N���I�����g�������ܐ��UF8z�-���V�E�Xi�	IU[��M��;;�5F��۞��QĶ���ok}��������.�b{�,9����{�v���,�%�Dh�^��ib����CӸ�3������$ciy�6���P*����O��t�[\��������<(���D��m������h�ֹvy ���<�Se�594�4X���C�Dͤ���,�)HT���Iw���}`5Q�?�=B�U	j|�/f���^��q�A�Sl��p7+�_�4;-id٬)G�
"}�A+<{� ~��as^�������8��ͅo��6ܦ�c��G��BW��7�}�J�_J��8o�+ ��,��r0[.P�t��Γ���v�J��(�S��PoZ��"�F�Ϟ��\-�w5��E���F�C�� �':��A������W+&�i����F�bO7L3���*����i��,����>�޽�s��UZ��I�n��[j�ZS�CU�H�	nR�����(X�/��X�k�f!��j��m}R{~�Ph����2�,ږ�!��PvU�*�OG�*Q1l��s�N+�I�������r�$g\h�sYVq�?�@qb�aA�D��ʝcn�|�f�W[�gV$$!]������V�{�Uqw�����]���w�!�c� ����p}�Zlw��锠\� ,hN��4Zt���V�n�'�W�}�	�U�-j����o�t9�1!3X@�
#a��1ٖ�;]�Š�b,�u��z�/�Ď�fA�?~���˽�O_�9f/"�0!zC�C�����j�X�`��O��ڇ��u�,w�]2���j�a�����<:��Yu�ygNa����),���FcxW���{+����jl^�xk�2��ޚ���@�U�umi5
E�gQ>�K���uH4:̯}�-�>�S�m��r���@E���C�zuj�:q�\܉MLA·�9�j��\�=1)���V�
"��<��«K=������L�g#��10��ph9'�.F(�@u4 Fh��Ghhe?Q6��<�����y8�T�5�`�o�|�/Rd�������hz����{������o�+?�a��RBF� �$�k����j%�w�"?�� J4)w���ͥ������g8��l��k�S
'� ��^���W����}O�'��~X7a.5����������脓(��P�Hdhoω�_.�7!0�D�w�jWB��kB���F�ӱ)�����xyq�Ț��<~�Jo��
��	�8G��<�9��oT���7�����:�YC~SD� �����B����m������Lۘ�_�x�@u���Ńm,�˻���!��s��LV����j�c�o��P�cC��`����W�V���n�y�����@��ނ�8%�Q��l�U��j�E�Ǜ�	á�i7�2k//��p������7Y������^��iȲy��Џ��t��:U���}����H(�n=n¿ ���]S�:�%��0>4�/���7i�Wx�TR��뭾�x��K�"���f#
v��_3<Ű������H�!)s���Y\Z���dڀ�|x��y쐼?zz�b�%e[���0�ipg=�����W|�:)魤��M�vl{&5�֡�G�*ax��&�(p�ٓܨ��6��-��/O����N�e��x ���vJ	��{�5���q���"d�æ�mh����k���}�G�������uE5+�Ϯ@N��ЙF�?�8���SA2�X��ɘ6�|�7�Z��!6���g��j~:~f�޸>׵�j�FΏ_�Gӵ�6�r�@<������b��\׾�������R��" P���8<'.���0yC[<��:n�B�/��O�zc�1f;\E�aq�|DrP���j��*DϏ�s��.#L�~DF�;�+]�����j��פd� �3n�ՅøLos?l5�C��5���hnM  ��-�t�oG�x4פ���=^PR=��H�/S�3z�!��*�޴�����;#-�A����^���Ō����\|��¤����`�P��`0�ө�����~�@��3�I#��<�7'��jAɹ��a�d�]z`��� �+a�و���OC�#���vy��fV,w�e�%(i����&*���rz��:C�h'�12r傿�{@�����XJ�~�Vd�h��4#�j��iW�s`VCN[H�K�{<��\��Q��TfV��]�m^��όc��lF�!�9ل NF�5��ԧU��~/Q��������ʱҴ�.��|Rz���5z1�k�����'Y�7o�"�R=�����|_�4��^�+�!i2\��I�����p.9fW�&ط����DOb>��ǓXq�zzH�&��	4x�d������1e�K@M<�E�p�x2utgw�;Ԕ��/�x�5���Cq�{q��`6%^�(�2̜.[���t�ƴ��էO�+��,ر"�b��U����fy������6E�O�����[�9�8����~��}!)��$�M~���hnc�q�v�L4�����p����q�D����Nh�1Ud`ꯧ[py��6Z�� s���m�J������=�����>����6�ΛՃxOˎ�t�+������ҫ�#��ڠ�Ј��w��x<d�DHn��i��g��o+g��m9b���nm���4�����Q,�iba�\�SV	寰��Jb���0���e�zx�+����"8"�M7�5�����s�W6C˽���%P��Ύ��|�9ʸ�����T/����E��=��`�6Ϭ9�
�8 {`��_dAA��Ke���;F��,Ow˅ee�lӯ���I�{v�fFSK+�ʁx�d`�z��}�LM��~�So}���]�l�\�p��C�gW��?�_m�0�}�y舌~�pZ�@������^�^����T�4C�:[P�e�ih��M���݁f�M�ZZ&��X�k]wdQ;����d��4Ѣ��}�͝�ͷF@N���������J�u�l``g҉�ߥ��Pbv������z�� Ը�Y^��Ϋ+��_=���~|{žv�3N�C+�Fڂ�����Q���Ғ��"̎��-n���9�|x���|��H������3x��n�-��*�����T���i���_��D-��w���{5F�=4�4��ض���kT���������Y�6-fU5��9��ן�=o��d�u�4F�!Л~�kH���O����m>�p��-8+��\dl/ʔ�J�~�o/���CԟZm�s�_<�1��0��yZEM^��:�c? �����K�I!�u��#���LRix)��qI��*x��j�T���O^������ȏ���)��u�~u�i����v�d�f[zQ0���q3��v傄"�d��Y��<.���qR�|A[F^7b�?~�D���{�l.7e����t~�?[=�H�O�)�.��,���r?8��^t�p?��;V�{/�4s!`BѰ�j���V"�U��GbQ���k�%o�Y���B�}%a�O7q��Y38�ٗ�qv	\�v������f0�{���ЋY���<�D�b�>GJ�6�������������S<�F*�"��ݝh_�-�x���x����a�5�h��"��`n�Mr�'�MV�c/���^��@��)�6 {Xx��^I�On=6ru���;lY�l}� \�)y����K����<w���)�s�ۘ�-�������}�A�yۢ/���ꂮT�p��x�9�L��@wJ ��d��}�)#n��4�ڃS��=�:�X����r���k����ύ뎁aa�BKo`�~������7d���:eDj=ss�L۲S��BQ��-n�ku㒙��^�s�]�c&�E^W!)S퀽�y�s�5&�'�""w�Ko0��*�$ܑ?���lʴ���mtd���j�Kf��p1���Z}_i�M\Je�w]XX�=�7�J�R��)2I7r��&�;k���H���h�x�'��i~D�[Z�j!����B��F�[� �D�w��e	�'��(�e�jO��6*��+���N��8 Q�&�a��&Ҧ��{ۣ�;��p�u������ԷX�����v������G(�n\�݇��C���k�ϓ��=J�.J�Z��2���d�.bS�b�'����춱��3���k{�v��}ԶY$�$EJc�K7/����N��I�Gu�?���#���R�%
edj�u���㪓��>��ڥmo`���[�ι�B�o����Fq\���T�z�p�t ���Ti�&�7o�u��䄅�9�\[��]���e�ˇ��o��q��nH2�ݎ��܅��f�b��I��C$:�6=!)z�9�s�d��?�܆�W�ܤh%�|����R�Ϳ�.%�R[ØU�����yf�0j������e��j�a�"؋{��}��,膂�` y3���n}m��<����{T�@K�ׯ�5�tb��r��yJ@B^f(1/���B?�Z
�w�V_{r$a׵״ԕ�i�|������a>���Vg�OKN.��G���=%���.>>���J~���ᡴ�Lkk�x0�_AU83�l�O���f���Y]�PXQ��^w~�|@#>^N��#l�����s����3���\L�T+�Hw��z���?���?
�!*���.V����z~d�Sc��9��oOM!�ܬL����vK�P�~Ů�4ZW2�H��jE[ß#虀��ݷ_�T��^H{�l`����k.��_-��"�����|�|y�����<1e�jz`Of�ɮ��,�ͻ	����zv0pߒ6E?��?�P�*���~����~xk����h0�0h ]�s�}��s��ޒ#W�cJ�I���#X��g���R���X�����2Q�
?3�;��pw�#}4&�&3>����sa33���}�"��������Ea2���Uo����l|�Ƃ.��jĊ�@�vG*Ed�os�9�څ�l����d�^p ���g��B���m%o���LZ"�R��u�W~!9�����=����v�Ff�1�So�i7��+�0��6��k����d�W�_*A�i0��O��Nv4羿'm�Ub-\D�Ծ����K�mZy��/ ,�_Td��bj�fxb ��B���^1���Q�h���-XL�%7�)�1��i�������8�l���OOh�\{ ��Sw���ysǀ����Q����gZ^�{��xMT<�<	�-6��'I�;X<��~��\�TY�Mg��Yͨ�J�%�l� �p���$�����)�o������]��D��eK(l���)�&���I���o�L�z}}���	1	��'*�;v��Cܾ��P&�,�9���8�8?}��+U��MF����H��3/�~��f|�&�X�lB@f{�;���;�G�A X��~A����m�).�Źs1:�_c����������ak�ɽ���[�r�\�H�O�}�8�k����ST�a�t�G/]���ĕX�~V�&@g&e��C,�Ȉ�{�Ģ+-Z�|��:W�SW�A?Y�w�J%u����r�G;>��{I�s&8j���jK��&q����ή@��6v�f6f���i|u�mykF�,<(ê�]�4��?�o� ��G�}���gW�Y�I����d.N��:7��:낈�%��`���Q��e%���Tt	.m�z0�Ƃ��ʸ��]旴��G�BJ�I^�����<�޲��mص2-	@?�+��� ���|�{2�|u�>)&
M�`���g�:L}k����-�#�f����k�O�r<�H-��7�Ğ� lU)������TQ
8%�z�x��t�gR���{��}r�4�+KĔ��k�7�$Q�/>�Қ��9W�告����~�UC�	{$��L�%=��ߙ��.��M��Գ���Q����U�@ݙ;:����a���T���B=���n�����.K���[{��nb��Ζ8�� /5�7�8g'��_Zc�L��.#X.6$��XV�Gɽ����?['U�
n:̫.1���q�(q�ynz���Tc�����!���R�ѯ4��	w��:�P�L�:w�(<�U��\!��/�R���P K�G���!an��C�XCJv�I���k���E~e9���B/uǸ��yM?��L�	pq�\Z�aJs�u-C��j�N�1�C��b�M�6K.�Ő�O���Zc�5l�)�T�œ;]��P�D{�y�y5�2w�W�Az��گ��pF/ʜ�X����@����E��u2X~�}ł���h7����IfM��7��<�/G��6$�
E����<y�~��%�׹g�<��/&���#���X�i�!Z�BJ �Ęť��߰�r)�-�뿅t>`Gↁֻ���1^ab�����K�	���|l,���7tŸb�k3؋�F����س4��G���=<�'�OK��ūR��Ox��rP���ǝr�g�{��;<m�k�����ȶg߾"jG29/Қ�I7a�r1b�ݜ����ZN�Ҫ��ޓ��\vm����),��nR�/q@qd��4H�	�f'�z�'F\���TX�q�2oy�����JZA!�
����ի�H���W����/��r�'J+���C��RcH(�u�K[<e!ca��e۞����ãǱFsΗ�-�Ce����q��+��p����5��u��u�8�w��l�����o:d�_�<��y����4�W5p%*3�\�7聍�w/�|�g�άύ��xq}}�����N@'Ͱ- �8zaƓ?�����~Hn,5���!XcY��aW˸H��-���b:15,wŭsE�}|?�),'�*v�w��	K�����Ǖ�l���T$��dq�2�~�VV��ONK_''��uz�X_�*:����a�m!?#�z�q3���5���G��q��k��6�Ć���I1��O��$��G�`Ii�?3P�����_mX��&���F�?�bG{����"u��N��@r��q�!h��������f�r��G,< �=�g��ma�3�a�B�;�J$�z�^������\��=Kr/x���>a ����xo�}��*^��٭'���ڔ(��G2���"����&0}�a�i���x�4�[�3�f���_�7w+�P�>x[S=y�
�7�گ<�!˃�i�n����F��$\0%�&%2����ª܂ZG���g�$��p%��cVI5{ ��+g�1m���#
�O3pYUFXW�Ͼ�=�X��4���{�чxZ�ƒ�hƭzh�I�es�&�l����ݠW���^�N�2J��)Lw�+��K��r������_�]�W�`�;O���-�3U��~4��X��b�M�f���bm��BR�<�[9g�L��r�/˂������MQ���r4�ť����J�}k���o/����õ�vi��?	�� �2C<t��a�j&��~Á��-�d�kݗ!E�<􄆪��d9m������+*�:��V>�����Y�Щ�Tϑ��9hd�7@q-��7Y/��_-�Xr�Z��]:,GFb��b��oS�\r�Vf��v��p�x(��c�r����JC�o��/9Efݻ�������yy��#���7������^o��L�w'�O��"�T���*�G����
�C�'��F��B�b,j�|:�#N]3#�ĵ����=��ψmӯ6��\��X�kt�I�9�~���(5�N7a?{9DuЗ�lX�TY0&��	~��Ux��ֽ7&�0C6�UY��Wܼ��6O[#dd�����	�rZ(_7k�ÝD�;n;���K)��B ��6�[=Eg�h��	��3Ew�o�o�Q$�d�#��v��g���/�����B��̀��z"���d*����5��r�O���Ar��>�h��n�����+znY��[LJ䕺x�*�/��HW�!M+;C��w��y"��@vl9�+�Z�]t���,��:�i�t�T��%hT�ц����<޻t�T0Y
�H�-��\�8�$I/��j�l1K�����'�.�8�8D1>���޳��~>�`hb��;�'�៉w*���Q�30:�#�P���
��p5�Θ�/]0��p�:C`M�����2���v	��ω}����)U��nR�Q�&����T}2Q�ր�X�%�� A����k:O9F�[�d��$�-�u������7x�a�O���l��t���	����E��'��}p>�+�SA�-Q	���:�Q��{���gn[�OD9e�4�@N�-��7����l�r&���݃��q�_�����Nm5���)QzR�z���q��v����%��Ǖkq�Ŗ���u�����Y�Ý���mW;8|�Uk�r?`J/����t�5�!��9�A��=R���jϾ�8�c�ӗ�;s~p:��V�M+;[�����Q�4�5�>�͑�d�ؘ�����BLOW�a�z����r�eѣ�a�����;�B���/�_Ƴ8���|��K�`�a�p+��C5�D�n,9ԋV�����6"E7� �� �|W�e8c��\�F��-�Q��T��&,4ڗ���F�n2׶�w���Dqd��cߺܟ��u�L��90S�w0_׮���e`ް?c>_�2��$��FL�ۺ���I4����a�/���{}UB���$�.\�B�B�vm.4b�nUd7�A�w����In^���p�c�4/#&����LLM�s�*��+m�0VQݡ�b�l�{�y#p�����U&kN���Z.[��+h�&��P�KK �Bհ|��[`�r_�[^>� ��13[\�G�����3�5�qB��������^�x�|���0��z�98�X:�RE�,0b0t�����+;<^ݞ������Q�%mW�A���=�a�+��&ey�T�pL��uj�m�t�]����`F �������ʠ-�_-AE����I���!��ꝫG��k���َ�%p5��9��6��'
��{8��{u�����)�^�TNӰ��Y�݋��:	1�ޚ*9~\��8�8)Ҹԓx*��ah&T20xv��o��l.�ײr�����`od8�����ug~75a5a�~��^5[�#h���Vk�C�p������8M����ұ���`c����z-"��-�)+b��Q��H�	py��A�ok�:6_B�8],>�l�<W���Z�5}��7n�u�(��**�Y�S
�̚��sܗ�G^B�}CVL��&@f:I�Š�#�� �w����Q_��P-�-�D�v>��Bι�h�vx��FZ´v��J���w��9����!q�N1����d�ɖm�6��{l���}������/����^n�Q}�4�����+�M���ye%^|8I��	[��.J˳C5����fdD|Ik���dTdJ�J�E��~c�g�$�rHZ|I=O�@%���ճ��`����d�u={���Õ���k:K���w<7G]��FK�Xx�L�b#w^iLJMH���G,�x�(�/��3���jLC`�Tv�ElAS=K,XA%me�۩w[�ɇ󉊮�/�Y�ŦG��%�yg��@�������vP��ᡗ"�i��Ɩ�f�Y�! �u�Yd;ē� �;�]py��~UN�]�F�n���MM"H$�@�C��|��L��
'�}4��V�������ʯmeQ�7,x$���kYٝ_�J�%,�(yI���|�Da��;�x�G���Y;�$~"�. \��7�#�=��J�'�]㧷���G�ͦ�q7��R�O�n��|j���C�ƣE�dq�\���'�������O.�rum�I���첞��T���"�Ăr��H�$rթ��Y�!����I��V$2
���G��T�YOʸE��w`��h�=X�-��հ��Ų7����ql��0�T(s��q%#���>����[\�M{����>��Q�6��<Ii	p��7&
��[nh\c
[nk�����^!�~��s��J�MN���� �!�&����R���u���	��T�_8=�:^�\����i�a�S�=�MG�N�����ݫ�w����Y�M��<�vO�x���}=�������!�*6*
��g'ڰ�����$�ʶ�sz�}���_��	���(�J�._�ז��~+vCn�z��_�D��Bj�2|+rA]�ƃ�Z�r�N@�>OaG��H����`F�'D�cV��zv\6T��E���t�ms~F�t�=DI9x�ۘ�Y;��1�l�vh���l���D�:�#su�D���,������Z�*�	���X�e�T��l����'����ԑnCp��U�~��WF�_��6ˌ->&�M��/[�,pi*--�U���Ը	L��\lm0=��t(�Դ>L�b�Ӹ��&){�O����6u�>X�SXޔ��������?�S8�tf�S<e��������@�3�ג?)�ѝ��o6	=y����x�'�����ϧk|���'���C"��##;��qSMyyy��1W��6�e�Sl�6�1|׬c.*���:����-�D,�t��> .�����S���'��5̜]���d��x���c�u5���+��Ë��EI��~n&k�X�k/~��Q9�6�3�F���M��T{���ԤGC�]�^Z�r�;~�Rܣ�ǐ���_7�aċ�X�j��S7na�Mvwy�w|�s�>�[�����Ebff�����őL�&)�շ5� ��f�<h	��,&`��Y9��=���x~y��-�y��^F�y!J�:���>(7<r*���H��������d0% ��,�pC���P�F/�f��+��a��z_��&pP��U�qY�I�/��������J����c4�93a~�}�Ō;8���;�p�/z�M�&�uч^�������>����{AsːG)�y��۷m��x*�**.{bZ::�#0����q�rL�] _^�_�6�_��ډ���T����ߊ��qb&��g��W��F2��k�#R�h����?��8�E��y�i^�L6�BlA�y�<�}�K�[�Z�ƨ2�'�pE�Y�^탆�	��y��J�?m��ף�OXG��^�F�6C��ֳzEEA!a ��>�J����9��i��PkO�AрU�UT���(#.#�Zw˙��%G4R��y#G01�"n�b�?h3�Jɰ�v;�ִ��=֍�.3�G������i=�x݋v�=>��ݶRv&�2`��g�}⫧]����F�8�J�u;J��$�.��2=-2)�g9V֩u�3����GI����L�o�\�8�u�I��.����\��m��M���g~w��d�E%d��dڀ)�M%����t> �S�l�������@,#
NdŸ���v<�d*�qQ��M#���-k��Wd\��O&�/���<.Z"RW�����F��� �W][��Wx���e$H'�T
�s����#�v%c�pct���=|��`�����Wƃ}'�y>t����,���n��b�o�ESc�d�|�M�z&�oii�Kw�=a%9�Û"~{(����K���(ْ��]{a�G^�ˌ��ͅGhC-��@��ˌ}Ï�`^��^���H�N�O�>���9�l�qC!��~'����"��;:Q�zW�r�ܼ�#�����E����K#b�`D�'Q�����Vx��Шk�Q�N�������H�;�r��4|�a�#pB�xE+�����o�*�<���_���⋷^�������XT�/�;{���R0��D����\�k�T�E,����s���:�L��YƯv���m�8������ѧ(���$+% ��;�CڹSr?��mo�G􄰲�6?�߭Ơʾea�'|���>��[�q#o�+���no�)R��O�~,� 7�A}���ea������o9���3����MO�����bPt��B����}�3�؉Ա��5ރ�9�$���u�CZ֒���e��q�t�=z���}�UQ��/�8j��G�|^�C������7�^d����I��JN7_P! RT���$����$�L��Ҹo��\)K�������6R�y9yK���֗��4�Y�3Q	ɹy�kV�T�eX�[�?L#!��(��t#��ݍt��t#  -�1RCH���R��!�0�������</x�u1{�����Z�0z����D�	0g��S��xTN/��sO���_���%��_mcJԑ���X�N�a��ٲ��HhX2��I��@�) �)}[�AFۭ��kvf.!���Cf��ٮ\��t���ɗޚ gL��&u��Z�q��,\�����mi�B�>��Ij�H-�(�<�rF�Z��aj[�Tڗ�D�S��;�F<F��I���Gp6a�A)NO~oV�����Z�t��Ѳ��>�vP���;!��)}���Ǡ�A��D�cǏ�;��0���%����WrC�����$��X�xM#P���ޑ��m��0�+Y��g�`M�}���-6���H�B��}A���.�)�.�1µ���$�>Z����%e���%���BA�丂^�T����
"�yo��YܢN�<���rÔ&�O��s��{�fS�}F8� �$-&ZD(���M��蝄j+%�w��N�#���I�l���0>���Z��=�(�_s��~ �d��2�C#��sh��?�T+b��_q���Bl�r�I))6�}7�K&��=AZ:	S|�!�6�" ؝lO����V���Nm*�F��P"�����D�xla�naI���Z_2��D��CJf�}�6�/M2={��h+���P��wgdA�jY��{tV������S�\_�ם$�[_Κ�]LⲆ�����ҫ{����Aǫ���Vm�R�{�%
�n��w�w4�������b��wM�L�h�8�g��"M�8�ӠT�	�*�v߹�UZ�<Cn�uy��wa��B�{���Il��т�q���6��Zoy~)������/:ӊ ��w��X���dX(�}�w>?
�Γ xq�����uH*�P$6�B��tR׹�v�*S_�����I�D�>�����R���3��r%�6Ɲ�@�KS���"������ə���-�k�P#<<>p���ycEVX�#>��pk2ʤ��L~�Qo4^�v��� �����ʬbt���²�`)��N�Cx�kvO�lcy��@�k0	�C��Vt�H=v\���CK=�0v�jJ0���k��+��	ӂ��2ؘ�~�D!�n4#��6��;&!\vĈd�!gp��#V(�h�5��0���Hz��'B3�+r�F_��>9������� ��-Δ�W�����ǅ	��N���������	�p�f[��&�T�;�_~�x��;���3j'�������Lac�U�ͼ�}N �+mϏu͖��A����Rm3�B܄*�Ǎe¹�e�o717?�>�_����c����C
@V�K��|D#S�̌��J���3��`��._�W폞-����nX��D���'���\�n��bͻ�?��5�?�[.*h�t��֖-odK�)�%-�:lJ�6��Ĵ���4�g�薪L�I<��}�B�A��s^�Zk�zE�C���0��/~�p�z�V�*��n�S��¬�J�Q�����Ќ��!�p����ö���5�4�%5~F�.ܧ��ݏ���ܰ/�+����ݜuRSU3hi��B�v���ym!~��Cu�X6���'n����6iPϽg,|�E+�WZy9C��f�<��x�0nQģ[;__��Kf�������&��Ć88��&��`�D�6����5�ܰ���Ү�������h�p+������1`��[ʡ��MwY�SK8�G�xKZ��J���	Ji��oC��Xp܀ ���#�2^�t��V��[3Z|m��NҠ�d�(T �z�;���;d����h����שWֵ	0:U�5��o�����KzLo[N/�5F�`棵����E���Gy��y���E�'&����0/�U�_�	���޿�:T���,a�L┽:-Ҷ�HIK#u�hE��8>Ͻ�@_� ��GT}P@ �2{**��b��'����/����&#�a��6�ؓ�:��tP�ն���U_�x�6N?f%���hXz�bL�\ŷk��bǁ���T�˷��f��������ߛ5�����pt�$�_J;l'_��%E⓾l|w�x�&z}+�;4�s�\ƿ��=ƛ_myR��P����T��?ko9�~
�ǎ�b{S���FE�Ђ�f�JKK�W���`���}]g(��'����A&�{��י�i؀��d����:�1��:V�2��S�Db�d�	��v�[(yg��J
�t-���'���wD���Z2��|":��>�����Qg��6*d[�'�Hg��PS��O�^Ćap��� Y��b�^K�䷟d�Eք������VA��e��G}��O%%��4y����?$�g5��Veى����gi���t>Q�cTQU;�Hb�� ��-'㐤���|*$B�/��<��e���d$RL!E�I=���pe6�wR@ޑ��a�p���[��
}�$��o����5k��@���_��Q�p���0{�*�Q"aH-{-�T�K�=K�#�����%z^uj}��u�����ЖE,���3dqc/)�^�Q�7�;��߉���������.���N:��^�f�G BO;X����]��./�v�h��soP����'�;��lo�d��:��$	qh�y��L�	����?H�o�ۑ6��x��Rc��ǃ���G>=gq	-��{��A����ނ�[jē� �T�ӣ6�����q�J�FX��ף��fU:���?��w�sr$��]��d�B���J9R�?�x�k����`+�������ǌW��`�j�Q��a�Ɣ�Y���[��8J�O�� ކ]��ԢR���7E����~2+�������I�Nr��O~u���O��ێS��IQ�[�E!fs��<�㎊���H3){��&�����L���x��܉��>�	$}�����O�1D�ͨ�IU���zW��{�����2u��]O3��u.I.Þ��+�KPH^͸�q������8�Je�9e�d�����j�[��Z]�ͯzS^��g�F-:���U�X�a����Sfp����
=AYٔ	7COp��W�d,JJ���r�T��8����:�WFc\���sr��oz�MY;?��L���{��u�7��+��L�3�C��G�<����寒򵎣�� ���w�Y������w{�)�GK���R�D� 8_`�c��Q�o[��r)8��M@�3�������»���� t� 7���1�������fB���Q�����@x�0�߳��|.�,hL�`���ME�B�	P��{w���V�j�t�X�j�c6�[�?|��֍\�H9�Vs=�	�	���BM/���큖�;h?`81VaTZW��M����T��.�ݒD(��0�盰�N���X�>R�Ѱ��-�6U3�b�@�*R=e�<���~]���05��wFvw\k��2�5k��V�L$��~@7����j�]�y������Y��������"�66X�&���MV+�u�L�2��k�Q��"�6vv�����@(�e?Q	��񉐭��J���fS2$�eÝU����p�����q��k0���	ц]�����<1E��{n�	��Z��AP�s{� �L=�b���rW�<��~����>/�u�3о;9���3.�:^�d�$��+�9��!*��4�Iԫa#�k<����7��j0��R�:C����7�}�X�FF�$���f���.a0?�Z�W��
Y&��3/���jQ�KR��'�Mq�~1�}Y�`'�OX��Py`������2��/EC���W#������@VG�5y{�j��[<��}4yQ,+�_��L�;˦*���{(7e�hODc�R	���P"�O�!�|+`�7h��o�w�!=���.s�4vǄ�!ò��(��OL��2Ѯ{.a���R}���fy;2ݴ��e��[��l_��b ������D)/�e6�e��zT���آe%���q@Q���I�f�WQ��?ߵǔ���r���$%���9�k��V�d�w !߻�)@�����~���U����m���o���fgz��7��3��Z���"qta�RR��I###t�H����~U����'!)����������{�)>&�᝹:c�FN|2y�3p�z06	����"����B1̒y|��*�H�}���o�X�d���6��Ï˥��Wo�zuT{we���<����d��gJ:Q��'�/�"^�kf�N�v�c�+~���|*����^<l����v���.���m����dz1��Oѳ�'���]V�,�\���U��J��$�W3��5��3E��dOP���x�sV)�Ϥ$0;�yn�(C!�Yp�WN�t��=
*8|u�<픤o� �y�:��Ȩwa_�!^,�׉kp� ������ry�8��%�5�
���\:t�����R)Ļ�~�&�bT�L�V�"��_^h]d袞�Iv�S��B��Z_�2��#�>א01�mX�k���g�=+�<�p,��E;��@��w�����¸�/����I�O����k:�H�!�xZɀ��|�@�\SQ �lmm%db-�������|��\X ���f[�Fyr������#��V?�Lv�@o��������݆��a�{JL�tFz� ��Lg[�'����NN���M/��k��2�b�7t�h����,�E��S6��Z]����<klP�>v{�8`��=��O�E}rp�n�_�S��{�j����J�/B�iUu5؇��p$@�m-���I�)+v�=�X��Z�'�0O2s8���D�K���ۓ�m$�*�����F��O_z�O��\�Q��DI �* "�4H ��qɳy?^���]!C����py�uǽ���%߰^!QɄ��[[�)��ɓ�I�����Z����~5��4G�j3,��t�t�Y��O�F+������㟭k��cSS����a�p[q?��D3����+��Zfe�+�Z�fD�w6�s�`�a�[z<#�:�����
o��G�_�����G��#�Q�a�m�b'����%#�F�1�]*�)����A��'�!����0�����`۹)�����������7�!����]���*\h�U�)A�ɻ/e����l/�׫�����@<?#EUE�9�jaar�yy2�� --X�P�Z__���.�.��Kk����{�臾��x(|A��6�B���e��{���Ĥ���-!���G&��m/�_E���u��;�c`q�LM=�j��	�L����� K�/�n����S�s�ڔ����O��7�*$�j�!d��	�w���aL��'��,����C���O��c	5eN�R��D+��-�3%u��WM�\�8�F:�)z�zwjy1<����U)�U��9�o�����~a�{���y#��y�=�~�'����s��w��d�2V�9Lw���^Q $L-T����]���L�j�vޭ9)��^�P�Y;R^=
���:l���z������I��ex^75���~�Jb���������<0�E��O��{��꥚���ib\������;*�g,��\���ed +X����.�5�r�W������G�6��������/�R�G��~ɮ_�sx����0���d��r�@�6g���0b�h9����c`*�],��0�����3t]��#{w�'Gb����;��-k[eb#�4����\�A���gE�x��%�j��N\�������RM!f��&@��7�<�$pK��b��-�@xM�`V�0���r���崸�R�SO�1���y+o{��)K�����O�%�Nm�+E�3\dW�kΖ�i�=���=�n
��9d��R�i�jJ�r��Na�4��U���"4�#DN��9�#�krr=Fee�#�9NAA�Q��`Gb��L��ш4;<$d��#@�	���b	�}�����e���1�g2�)T�L��HRRk;'��r�Zh�0��<<2���9﫩����㽰;\ � pѦzu7��{m8����w�I0��_Ow6�=ǎ�/�l��F��F2M��p��^�ojf�^����mc�� 	���ڈ��F ��Xr����!��Px�/^�m�;�r�ca ^�� �<a�,���f�m��+ٴ��b�yMW>�xM{��N��HĐ$Y�O+��ɜ5��T���	�.~��S<t�%퍤���}����6_xmooW��3�AX�Ɔ��V�i>[y����v��7<|<Ai����7�4�h���Oϲp��jK��@��u���!;+�/f�/9������=��oE���>��ND!66�c�`pYX�-����.©�T��[@G\�d��S:F���}]����U�%2�5��W�:�`+�w/[ـ_�
'��G2�I�����͕�V�F�%b�Svo�agD$!a�0l����ޗ�L�z�$
��<\�{���!mԩ�F�93��|����T8�V{��C�]/��?۰�T���Q��B�LYYa��+�B�jy����T����M�G�	�#��֝��Zm��p�9�#�>G�wn��a,r�bs�X!#�=>�)�m@��c����%��B�����a� ���>�����)7��3���n�潕�k<�6���]+ߦ��O�Z��55�8�)Ē�l2��P��m7mG7��Z�Q�ЅfGRIIɲ��ψ�'E\D;�,b7��F���u��5fTy�^ASJ[
���]cϢą����5�9 �׭[�ݲE�g�)>dgZO��V�s=s~��_L�T�����w�K��R1=^DMB�1` ա��:SZ���S%%�|ji�z'�ak�U��}}F��el��;�"�D�/SI�~�-�������,���KD�j�}���
�ʕ��5�x���qy�O&�	k �v���g#��ԯvK�0O߻g���x��(Tl�U.O��W��c<{�����ASzG;Q�8�Jdo�}}�=���3��W����>��� T7���f�&`Q�/�]��"���8T�* {�E���Gc�f�z�CO/�>xv��/��8�{�ZUt�Ҍ&{:4:�ibb�>�TY����|Y���6*���-O�p�wm+;;��EC.�����45[UU�< ��yx��%��Dd�\��" l��E˙oqs3��R�M�K�E��pB��qo����s<tr6gz*���=�{����Nm.��W�L
#�Ap�D�1��&�H������㚏�1�gQ�p���Y���W����ܾ�Tl<C5�}�
�ׯ�(ʍ��C}�GU�|v���ztG�]f���i\O0�"���6�`�KLW�Qn�βC�綌sn��M!O,\�JDWk��R�S&��-�7��>hu�=�[�Y��&�ޯt�ȷ��ҺNgf���X1�s[J=[j5/̆� a�0���� ;�Y<X��8��ώ����T��B�;+T�[�`�-â�&6Z�"gqf�>������a�������Y�p��� R"ù+5c����c8�&A.�C8��Y�_��+�<�M�!�����@�p?�d)��.��v���������"N����j"�]�⌊���;;���I��|��ݩ������h���SWG����5`��Ğ:/|���	�;�k��#�3�(_@��B�@�u�����Lx��nq,y?��ο=(��6��iJ4�0�dp�.��Gk��\Ȇ����,ߣ���ӗ�o�L�n�Ok_�/[��4$ y�0�NǃZ�xR�������ӊ�f�.'!�{V������Kl������W�+�3��T�;/�魥X(�s7�yl����������ؖ�ص���,���n�w~2��U�����cXHt���
���Bd]uף� ���p�h�D�_B�V��m3[����OԎ�Q��������X��{�7�r�����i$����=Q������D�Ǜ�+D�f���;�lV�L�
m�D:xV'2�V�W���WC�����{�w���eb�/�������,y�0O��1h�Dʟy�(o��C��M���S����p�0��nQU�!pR�3f�8$?S �Y���_+�nIlf�o��B�"|5c(���_'o�aJ嶚8�N�9ԏ:@>2���(�鷰�8�z�����[m�7}�cr%=��k����Ӣk|II)F]�!d,���w�+�at�M�s�.2��5���VN` <t�pi��soមk[0����߫���ҧ�_�/1Z�����K
�X�����!�@~zs;Y�]Jŝ�#G��������i��C ��TTT����WR�'
���D����k+|&��L��f���M�ϵ�8�ͯ�04�Z�����l�m�x�M�l�/��^fe������;�e�\ާ�;}���z���i��zB���?�O��z O��Wi!�i�}V�c�8V]九-�1�_'i�Lj}CA��!�;� �}]%ů�\�Y�=3��9��n�j����Q]�*�����G�}�F9C��q }���T.AF�'ȃyڃ�p�_�F'���O׮���Y�r-�vҠ|�3z��&,%������J[3�IVN�8��b�ޱHh}��n��dG�u�7�+}h'`&��հ���SA��c�R#������Z�@\�&�g��F�c�[;lv�Uƾ�_ 4(�B�oY&����F�:��ޖ6�ܖ7E�܇:�M=9�ȏ���`�GL���T�9tI)��M.����w&���F���nM�u����x���gAPWbA�e�3_�d[�t\��O�c0�y��ɬ��T���g�j�M���Z�P�������Y������X�`kW����Ŵ=��v�^�9�z���u�l�R�^ژ�����%�U҈��d�#�q���n,��oP��G��ƍ�����j���Eg�n�<aŕ� y����c� `���v,���2����&���{.K�E��q��'F���2��8L> �p'*8LqN���1�*5g_Î���<��}[���
����,��=x��1P�&eb���[y������`{H���ac#L7����'��饈>����.�XTi���Sצg96yz�ƓP���[Խ�>o֯{�`pi_�#
��j�����\ScRXt��6�s�=���$۾�f�8j��SƸľe3�F��Η�S�Ь���"q%�?�@yE��b�B5 4O���IBϥ�Y��刯`����{���U���� �F���t���/l�J�قf�^��s��2�L]��H����/o�t��|-���(L������дq�^��4�U�?J�gy*�μ�}`�W�|5zKmcbc�Ng�ĩ��) {���p�r�i^��:�=��9� ��IJ�ZQ=lԩ�<��>�pʯ1'�b���x1TSF�O�3��)��}�kОM�����R�?��'/t�r��7Ęo���S\�ש ��E{�ԯ~
{�����w�@���G�2��N8X�:X�"���'6vKO~���U�۝�d�^�����)�.�d4�o��/��ܖ��'�^0bE��e�[��fl�!H���7�ӏ�[���z:n5��7M��H�r�vk��;�����{��� 'Veoo�����a�_O%&|�9- ({�;��^�v<*��{�Z�
S=����ݓ)���n,������Y�ۻO|"���AE�WB!ɇ�h��#��w���c�ںl_Ӻ�m�R׶��@?�ig��%G�X��U�pG����ZK���#+?~Q��S.� ���AS q9.dH�����H���ݛ�o���|���@p�,I�{)O�?DN���8�I�ox_8�0�=w7G�eevoM���wM�x7>�W�<�=�Y�������b��'�grl�,2(�3��::����c"��:<�yF�C���o�0]�!ߟ�\��	=���!6G�/�rFq��Oh�Z���a��TG��g9sT���[��9��Ɍ��*�rm�tC&��z�[���a`����	�q�Q�P��)���|�k��{�p�6�tg�z�����+�`>pw}�
�z��gNO�z-A����>��HtTvR-�n�� �j���Ĥ���:���m�ٖH�~��8(���'Se
R��Fz�e(-ZR[$�YP��`T�I%�u3P>Uu�2,��xb�_P$��\���U�A�N}����&�/�>�a�Y	:*��Yy����kۛG���(�¼������۷��JY]�l�9��h�|f��&��Y6�2�wq�8���ĚK�"\&���ߩ�^�������=*�u��N�E]�E�@�����ͽ%>'�FVo|�U�{��o/m<ݲ�_�Ϩl@|�2#��yĊ�v�N��!���:���O�Nt�4���Z�\����wkFB�Н���=�;�t�C���E�C�����������:mtz�Ɖ{���mh'���C�\7��Aq��wؐ�������;5���y�\D�?G�kQ!�޻Ab�6���j, t4U5	�(h���_���	�pHߺ�1����	��Խj�b8r����+z2�GEA�p�H����s�Xs]��}�gR�mPG��m��s�n�B�������ϟ�m���9�op��$.�y����ָ坠L4�Fx�e9X�F�hq�ӈ��vɴL7%�v�/Ci�� �~>�-:t�^d�Q�HS��[ʑݧ������_��B�8��i����Ȍp�黿��^`���N�4�VR��U�#ď���8<�)+�vIe�O}=�q��8,���A��#�#��V`וM�xH+#����A�R��z����y��L�Ċ��]4x�9��ږ���uG�E�ތVg�7��8���$ r�螯?{'��6�|;[�cP.��(��h��/�j�oku��
d�T�}����m�����3���I/M�{Tz��)�?� ��3�Q�-�Ɵ�A2���i�
� z��)����PMOg��&I�a[/��_��g�|[,������p�.6!�Ch���x ���D�`����B��cߧ��'s!O�{[kʩ�:ɞ�=/	\���vJ�����M��}b����z���ug@?�NB�ރi!�ߖ�U���<g���v:���/�m�݌I&�u��充[|��0)�4��(�~LП%Ŏ5��F&?DxG
Lo������].{p���V���WٟxcX�j�ƝTQ��b� �П�X3%�V �3�8�&<Zk�D�,���l�uT�{rd�DY�� {V������2���|N]�k8�u�(*��[#�����zqj�&��a2�y����isr��W���Ϗ)P�1e�U�����g/w�?����LR��(���2d�����C��_2�Q��T0J	w�h¼������~�x�v=24�r��EC{�����w.��{�P��������+�$���Y���ӎgY�:>��ue��¶1՛1�"�^���%\~Ad"�7]#�ȭ(���	1��~ݴ;�
�ZI����5��]E� ��]'6_X�AY�=�|U0��d��:���݀��i5O2��O���[NE�ZY*8׎��/�:��a�
����WЀ������[�z�O�SLI�w�}B����c44vx닐r2/�Z	5�*�^R)~����~�����R�=�G)q���o����{���=*$��_5i"�7�-%goܗ����lr�KN�����Z ȗ����t6M&���) Dǰ�U8ER�-�`�ߠ��񫷟o�m�g�Q�2ӳ���8C@�AA�@
z��H(s�Q�W0Ц��	He�� ű��BU$�Z֚��U@���_<���p{�(���N�ޅ�CKwO3�G*�1W5���A�&E�������)�������kL>�D�,5&��z�{�-6�^�>YC2�w���,�×[eP�mfoǢ�
1Bd��:��?���~L�OKVnؤ�U�E]���܃m+s�0��L�<�����3&�7�i������Ͼ�x^����j�&k]���|��>$h�+y~мS�qp*����T�@�m0:JЇ��2���[��)�kM~���B���yG�M���M#�����B���(٭-�ɋb�e-U?�{%���V��\�.=;��m�����2~�T��~<��L$�g\8���Z^�69L�M��c�B�I�]#��!m#�σ��)3_����vE�lk����q8س��jV{�\ʱ2��+��x�.��������K{�Iar�ĝA��B��1���l�_H�+�ф�곲^=1b�`�c��_������6� ��/X>�V��Uv��-o�x"4����4���&)3n��(d��B�z5�>s�za-�n���&gq?<�yI ���ɳ�#W�H}v��p�V��i�W�_}���99��n������tϭ�I�{�~��t%+{P�u�V/M�t��4��w�������S�ᢹ��b�4,�S��^����n7�鵫�R!��?��M�|���Jm�Rf06���{C�s�4iD��=d�6�|�sص�T|f�Yh�ޒf��K�+ف��|�{�O5ܡ"�?uv.�߼>h7��p�Jr8�Q���<��$����i�7���_��J�E�ռ��c<�	Y��V�H?6��5� 4|�$s��X� U��#W
�)c_t��8I"vū� ��G�XM�쇮Qoh��\k	���;��Q�.���@��.d�2�߯l3���e�����UkM3*F˸����`��wΥ]@����G��;����o�Lw�������v�k�I!�1���;ˊ\�hS��j��<,�R�p�N�e��Ƈ��˖R�0��!��}��Q$��[���Z�y��ҭ�8�r}����0��mʤ�@y�Q�/Q� ���q��c;�)�9>b�gP����މq��
C�l~��d���d�i�6��W�=����m��c���Ο>|f��ܬ����_���7��kDav�)ᵅ���g��BBdzN���h�ke#�7����m�\c����F)��g��WU�(�'��:��+;@4��QK>�[^�d�Ur'�l,�N���mp9iߗ�c!�^lc���E:��D0u��@<eS!j�o�0L� h̀c��_91���	w\��  ��Y�H��z='�ZH��n��|Oh�`nr�yr��^�nHҐ����W��*^A`O�l�Ƕ,�pCyEMQ ���~��5�կ~�Q\��[� <!^��a�y��|y��)�b.�.-��"?���%�e���z��� 5���V;{~*8���
FBW[��S=@�3J'���U�	��}��YZ����0w��l$t�y�q�b�>�B�@��X��+�m��}]T��M)X��K���r���h��|���Q���{��g<�ʝ
�k��A�>7��)QN�V&�ט��>�N���C%%�)sn��wk+|чK|�jٔ��f.�J[�ЎUe0��a�������>n�q"���pws�Py;vwE;<2�-��ϟ�^_�ȩv�F���e�O,�~�������#�ͲX(4*����k�"�@���������f7Ə�K %�G��jumF�/���3��/;s�Hŝ:N����|,�/��E�s���~�?�����ō���L�4l4���L�Vq��t%��P�q��W:`�x[q��.�&~dY��yՔϚ/IL��5��T�x �"}��/^�����.y�%�fZ�s\�Hp %�	�>,��Z�yk���ׅ��2�4ǡ�|�?"({>  +a�=q��H������P��zJCf"�nj[�5;�;?�J(�m��ƫS������?1�#�
�#����`��+��G~��5|!2����x�r��Tɱ��tƍ
\8���lw��R�͢���є���m��DVN
G�;�kg��q�	�s��\/E'�(�q�RΦ=��7Mr~]+G���?J[T%�7n��{��$�3e͐>�k�q����7��b�2����iW�]�(�⠳\�m" ɗ����߹�7Z���F� �+j�(l��c��j��L0Nxt�4�`��o4q�ڦ>�¬�q)l@D@�FqM�zA֚���(�\��eG:�{վ��30��Tx�{_p���wE���X�*(q�kW󽅳cU�r���ٿ�
Mʞ��*��	NF��`������F������dd���n����eP����w�S��߁@GQ��:UW�����������)	�Z���x5%bfG4�5A�!8CeN�~��?�z���υ궊2P��;F՛�7��vN�����<�����L��I[^q��tKATv{���'[�iF�i�,YF���`Sח�ɏv&���rOt�X?��aLa�t]*d�l0Zv�W��A�A�L�L�`��:ڤ(P��~nE�v��1;�&6���J��r"
�`n�T.�u�}�k&Ch>�*�k��e�U;+EqS�Ǐ".B��2?d !BN?�;V����2y���W���U��>���q6�qy�1���<�\�0�n�aLaWgv�q����9�����.}]!����\}r��)ͣ���=��j����R��	�V(=f<�k�fA�n��Ι.�U�D]^C$)$��o��{_MlL�dwJ8h���F�jia�mu�j���Z�2��>����F��^`�9rPӇ]����*�
�1]B�a�������Lj��f�:AI��ON$��6}m�&d��
�u�*s������cb� Qo�t�����R��$�f(��Aa���o�j�+M5�*�oh�U�g6��jk��qZM�?�f�O���M�������'�F�s�Y7͵�8�_����jܶ�V�G���ݡQ@����������h�6���>���6�={�u}2�2�K�U&�����bE��F2�%�.�-W�I�Y��dDK[�֭��1u��r�u��Q��և�||:c��/py䵚�ij��=���+�A���]'	��2��#�krX������e�_���-����u�,!m���(���(�����!R�aYki�kly�'ü}bT�������c��7u�'��D��	�ix%��+�Sk��&� )�f�&�*(&%�F?k^�HD&�Y3B�qtys �e1���|n����®�����o�1��+��;ٗjj�{X�c�⟏0\���)^�T�̗/� ����rW����Q�D�$�n����}���m����D֋��O���k������X6�����(g���<�����l�]?���4��O�X�k˶
��0����E��q������?Ǫ��C^L�엔����FU-H���y��thp�?9�W���.��B�>o�qb��������j@�f�p�]A�� DC�����`���x���ync�z6������y�4��_.ڔ���{6��a�8"Q�L��#��/#��Q�I`
��g/��������<q�I������������^�a7~f/�g<�Pƽh�=��-������T/&����u��z}�C��J��'��?�+���#��o�JT>e������m�R�r�[�}U]MU�i7���U떕d�&S�����C|���~�T�]Џ�?	���)�r�7�4x1��������~QD�yB��i3+�fd)��C�;�	�݀E��,i` �s���{i��7��?[je$<S���cY�`U�׿��*׿��c��9��*{�aV�.!0J�g#�L�V��c:�G�**\��(^o��(�հ�US�J��I� uoE>�	�F� ��f����ui�h���o�q"ZחE�h��ZK�΢+��&�������T�-⫔�1k�K��S������>��78�lvll��'�ITܔ�u���}���TK�fvl�HE@Q5��d	5
o�d����5�kQ�֔�Rq&`)��mT������ݗ��u��w�{��J�q�7R��A����X�7%�� Zz�������2��8o�ɻ�]C}j Ǌߋa�hqF%$$Ե�+<
����i_�wIGU�\�!^ғ�M�
{�~0��uB��඗+����T��a����$L/g�3�a��X��� FھokZ�N�n�K�A���$J�v\�n�l�� ��KGf����{��2=�S6t4���u��Ń6>܈2��t���~�<IBdtt��،ŏ%;$|����a��'#{k�@JW�C���غ��?  � �a�Aʹ�R�1YEPX �����K�6|��A�f�\�G��J�����:<�.@��-^KpY�%oou�]ng�&�����w'v�ݿ�'�U�ї�CA��?�[�/%��.�f��^amc߯�oŋ�ABT����15%_>2	�3��`�h\x������/��;^͓������ZJ=#��\��8NK��`oio�h�F��y�+�8Ō2{��"5Z_�(%������}�d�;H �ʞQj�M�;�4���n�Q_����a7��~��|�3��Ia���\���ݻ��Y~�^��✻��W�UWa�ə#�\�ee {zz�V�n�>����G�)����i6P��	@���T~m�BP���ؾ�u���2+`#n Aw{��;���ш_�$2�W��+��X��!毷V/��uK�*q��jެ��費-���.5Yc�0JF��-{1B�
��=|EIIY�o������@�:Y�U�<�Ƣ�m0�2����CL�Cp�mlR����>௦!<�����y�=+Ǵ�QE���zd�� c���:�=��9_�������G*�H}���q��������L]��͹���l�|���z�k��~\���¯�uݒ>׏�;��S������M��ׅۢj�ޔZ5kojU�Q#j����U�gѢZ��,�v��{� �.�D����}�?�~����9��s�9J=_
��q^q!Gf���*Z�_~��W)�CѺ_�-�&$$+�ᨊ�<��i.��8Ǵ�����xs����E{���G�Ը�{,�Խ6y�T�D�W7d圣KA�/���[Q�@��P!��b�Dv�|��~Eyu5"����ۯP��ײ��~����K���Ŵ����觸$6��½(�5��pu-Wп;0<� ap����ϧ��e�Lbu�v���ͺ���e���v���X�#pBh�zlNWق,����O�|�G8
�G�9����Rc7����X�4���uz��Qg��8L�:��*��N����p��PG껕�3Û?ĎX�i��f�"K?���m�J��cLzx}�t��G���2�q��L�-��7�_�PG�����x���0�~-,Th������\���SSs�{'`w����b��aT��b>J*����0g̕�>�es�zaR��#�t'a3�j��N$i���T�mG��>�l�yZ.�� $��z�*�����s�2A�#˕){�X��9]��͘��d�[OHO������AU\�ԁ�I�e�v�<$����2?�����9G�A���R�:��+-$�^�X��������7t��N�v�./���!gڰG_>��>RF\�}�.Q�u��Ӣ�><�&�����a4��f�����KV�l}�TCBҶ"�la�.(�nڤ��%+�n,�~{
[�=^7a)D��L���%?���;}�s���yHQ{E�D"7.��lc�T劌����=4�E4����ަ��>m�F $�n-P� ��c��!�b���r�������)�g��d��~�������踮gl�Z�"h�iQ'R�Iԭ�Z�
H
�g�	��ҥ������7���_�/E��͊��\Fl1%�O�Uf���gS6I��[CZ��}je9.�S�����J-�P��ƛ.�(:L;��E��J:����*�X��^��x�5���Zb�e`U2�l)���T�봸����c����O���/`�:�z�I��������c=B橨����(����g�Wxڟ�$�/H�gK���ݘ�Urjm�L���#gu
��m_��[?��|��[!hZ=NNi1zq��|X72����"y�*���K|��@\�t��?T1��	�s0ӝ���3��'f/2�}g�ZI��K�2�/C�V�"r���d���#l�d����P홍��Y��lgL	���ψI1t^��z]�^zeQ��,!�j����(�k�a�,V|��˨����Q]
� �N��C���*����S�D�����	���s�Z��}��ɟD)jG������S�&�}qs����y��3�
�.���'�A4h����`�j[�k����±`�E��M$�d.�R�����x��B랉S��Fe|+z�����lڂ:E�`�X �qa��g�&�/;���~"/Y����P��{�w�8��fk��yB^N�z����������u��Ie����^���D�����?��66��L�sb꭭n�c�ЪZ�oEd#8+��oڭ��;(��&H̀�;��O�T��
`Ig�2�#J����H��Z� ܰ��:��%������[��z��L|�#��ϫ�N���%D��{�y��jIF����1����oEzb#�l��:�6q���>\�_��`���ߋLD���nC��uk��0�O��.J|�U)J;#n��:��8Զs
���r'ӑ'�/{To�iڐ|���������!���xGT�秠��)~o�DV[���}W��߈�k���1�����sttD1���E^��3��X��y��X�=Lc{�K	��Cvs����#�輻�3;���j2�>k�����`|h���Y2s����KT��+��ȂuJ�4-�[��$Ҍ\j�r��O]�]d�w���!�XVyZlEf���'\��L=��;�q���.cOg���������Oš���.�-��̜-`�"�b�8b�C���q���C�4�B���8;Z���;��f�烼WG)�+�ߋ��L�o�� �<h�{�Iԅ
����cS'w°t�:�N�tu�@j����xsj^<R����D?��� ���W��Y�c����o�'u��
b:ְ���C����۫ߥ�)̷Ǳ)���ψ<�޼���WYƔG��C|��:/�|���U1��[�������8G�z�����o���F���C �J܍�]�
r����F�����k�>��
���'�*��-�J���\&���<��OM?,�38u�e��]E�z�o<j���q�<cˤ��<{Y�]��y���������
l�<���#z�̼b�.�*�x�p�����,�|rK:���:r��]2�+ɓ���K�|@@������S��X���co��j�9�.s��r�)�-�ފ�12������6�a�>������ǫ�v����^֓���K5KtV�������}�pY��?��	���_��y �w�ܤ��.4��{�Zyؔ��ύ0�+��	�<���jĥ42�X����8e�$��ڕ�n�?�l�-%[���֗��I���g.aN�C�_Z��J�Ը;�b1�x<�O�j�e������(�]~ki���WQRz��[�)`��q$S)k)d��|���!gD�0o<]�dwߒ����f���&иf�ēBpڂ�{d���o��U������"���=@�}	��T���=
�s�a0.�)���Ϭ�E(�CNc	�2�ٵ�}���?���:t�DəC����nm�K�<F���0�Y�$ä4��#W?	;H��T$&Yi�_`���'<k/ŗo
"�_0�x��@��<`Y�e/�7G�B��;�/�̷#F���j.Y2h�������6�W͏���ql�k�3�"ޚ��*�)n=�hf�����mI�}ڷ�I ��~���t��������O���������b>N6�֮Yhz�9��vY��9�"�6���7S�'���b�K��C��Ta��魍��=�q����J��h��A�?�5��X�z�,�BH/�^�qD���q�c������C�^�U��Wm���|]�4PGl �hF8����n耒}�i�Lo���G�=4�6ؘ��I��lnT��oG�d��4�oE|LA��Ӵ���.�i��2��(M���ֺGQ4��Ҡ(�eyRo~5a�?˿���0^��\n�+HJwW��_R�Z9`"2ob/���$y
9,�,2~��OnO�m�X��PY����7��Xg�RR7-�n5|���-��_hp�"Y.������L��IQ	()�?s$
M+iL.�_]@���Z�֬Q��u�>%.��4-]���&:(��T�6��T��xY='�S���OP���{�7�ǥ��vV����j8���97t/�hyς*��8��5�m�h�����E4��d���c��h�ѹV|*����G
�w!�$�͗�Õ�{���YX�Vp��&�
�pe-�PDs0p������O6cIp D�R.�(dN��i� ����J�����*S�����!-��䬸1�x�f$��@�mP�<j����%`%(e3}so���������d��<^[�S�N�q�(�:�`N�E�� /�T���/Q#�Fd��G��vա�_K!��T}i�bџ���������ة�y'�
�~r����d5�%��e��F|z^&u����Y����@�ި������YKk�i�6?͙q�x�]�/^S�`��0[
L�/�����* SS�¡�����%^՛6�\F����͗�1�CÂ�(ɦ������%���O�\0�v�A�R�����ӿtc�S1U��P�o���&�r��(PF��*>i�շ��!ۘO���+
�9��ח����
:$�mM�̡���_&��-$`R�f��k]7j_�\�5Ñ1�g������R��[	�gۥ�q	V��ϡYq�!H�9؟P%��2y�Y���~ȺY��OW�vX�xBG��|-T�tY�;���G�l�q��O$�թ��l���Ӝ�l��C{���'�ԢeK�9���f�
x��OAa��Ѝ���)�/X ���4�?H�eJ�r��������� b�#�9��A�[mW>w+1E��u��;��g^�
�q�\��{9����������|���M�' ƛ̈́�u��񞰣Q�^Y���c�b)�Dě�p��E�9ju�GsE�=�B�S~��Wى\�l������m�Հ�HG�In��,!k�f�b�#�v�cӒ}�� m��ju {Vw]z�/qu�NN��&����ZE��O�?���� v��-�k�mC|Y����[�G儙�e
m�f�+��� ��X�N�$������I^A�ӊ76JJX���'�������~�`��G|+�DC�8n��8����Ֆܦ�,N��秒��M�Mw�(�������=�3��-��g{���{��ʞ��bhʤFj�y����r4��obAhf���/��ux]��(�����<Js�]}�2�WQ2r���`#�a�HK���-�^�Z\dpԽS��k�?1�
2ϫ���lu���a���v	6#�C�{���3w֚�Tª�}�j��4�.E5�u��y^� ~FjlĎh�L��n�ΞI" ��,�^�ǥ�]n��d-6�F�~�$����xX�=�^e�dI![4k�3�&(#���πIv�8�Q��:�)->��T�-�Z�h�d{ZFq��T�M����J���je--"��Kk�OB%l����u�N��`�s�$��YKy���Jz��j�R�S�WU���TQ�)��9�S�ߊ��H�3�����f�P��IS~����"	��h��@�o�|�u�_کljj�h)`=�Y�w�}���^��|
 	�^�|G�ȍ}�݌��m�z��]>�D$�����\�СN�ͪ����'_�q�?y�vE䓁DV�6���K��vYHk�ݗl�"'��+	���hgE<%H�F��p�a��}/���ɷY��7��-���������V�����e�����w�{����������M/��?z���j�{;���¯K���&ce����[����s���)�+T��G5�� ռ/<�8���u�T�a�U���g��5=�zWQ��s��Z�9�XH���΃�z�\	�=�\q#��it�^��=a�H��_H�j�1���n�s��(�2��O���B��i3���iT$n��G��л�hʟ8Dl�l�sq/���.���t�U!}ι/.�M�|���2��L�R1���6$b]��vN��Aǅ��S|�4�� ���
�� �=���H���v���[���b̕���1����~^Q���N> p��F6!�x���җ�:�L�r��ԟGȽ�ԩ�R3�� �`��8 �0�nz��;��6@�Z)��NR�m;QNf��~,�ޖ��ھ�dY_x��B���sDD=��W�5�t��D`�u=��I���;_�E	�,���ܚHk�8���ӗ�/�4Z�ih���齌'G�.��PH-.���M~���]hl*z�_s�]kR����O�ݞ�>�L�#�I�k&�-+#b
�}�����Cٔp�5eZ?k����5�׆{��[C{���i-�ʶ���as׷���V����kYJBε(��g�J�DFPo  G/=<jꙋ[��=a�.!���H���;E+��=�WKL��٣����Bo���Vu"��nq)�4t,)L�#Q]W(��ks�8��Ӹ���z���i�2��&�4 �e�E"@�ϝ^T��y�#7���D�<;���ˮ�Q�`;���K�`3l�^��<��̉Y^�s�w���A��k��%_�=�a +��o��%<��Wh/���LE�����
>�o�xE{4�t'h��1/��Z����R!���LY�
<��_4&����2{O�y���x���+��Wl���G[�d����kA����$�]UX�+�%���^��H&��D_��E�Ć9��2�E��qHcu�]��xT�"hY�i���s�ՀvL�It����f`jʟ�r��5|�uN.[�����.!0���Gy�ܡ+вE���A�����;,�!�^�7e�b
yI0em�]5����qU���E/��Iy�R�t|�{̣A��pW8Q~tt� 3�{+!�T�0Ǚ-ݯ	W^�G���<�0\A1_���/��1��})��eNqFb��9���jo��
���p���#:oKO-}���>��76�-8G��͹� ������w�$�
by��L�]݆��g<M����A��o�4E�)S�q�&2bx9	�y����w���0&0�3`X�r�u���H�V L������U�֔�9��)$�6��qSKKIL ¯���C�ʵꯛ������� �@^Ycy^��9��F���Nq}@�_�ܹ,�	ڽ�x�����K}�r��;���qdFF�Ѽ�����( �*�aYZ�$�|�G���%��j����#��'�(�<�O������yq���N*�%hմ�[`�n�番���|�y����G��¡�ЕX�omr��������OH�=WH��v�d������aA��aQ<l�Op�N^zn����n<1����2�?.���|�!�C��N�gi.�m�XF2O�
���+��Z�xA/H��s��҇������v��Q�^��=�5���r�g;c�*���o�	���X����~+���P���C0�-x�@"�籶�͟WD�	^hu0�^w�kV�M*!0c@k� Z���������S�(�q9>�UͿg�Q��O�M��(��cm���.�wy������F5?��`���|�f� �,<�� 6՚:�=�'�2hn��'B��[9�$tRy�NW!��t���8�:�|B����` �^,Qߐ�;����ѣ�F����3��]��ʡ��C��D��c䈙�[�톿u��xA�#ALK�;��Ñu:�à\�Q�N�����j��U�P�g��a��;crON�d��K,+^�,���p�b����.n�z
f��I��E�y����a�U;8!�N�H�o9�����X��ёF�w1��Å^c�Pe�Cg��G���R�^�����n`�L{��!3Z��P����K��lT?HU��^Z-�Z�E(���wg�Y��@Ҝf+�����A���0OBQ�
`RI��2G�����n<��R��G[Ӵ��6��>�c���
3���R)�%�
��C��J݇�R�3����'o\S����0�-?:fw{�q�ס6s�ς[A�,~�K�����NN�!鎓7�L=p�4�"Z�j�A&�˟A�/���fW1�4�v�O��]�d�<���ݧ���xm:���9��^o~�X����*l����,K��v�z�`4������H�j_��`��\����#���m��Z����r����@�,[�PD�S������G�O�/�.+�䀤{��@�j�^�iW�N��n�MY�UN�Eƣ��'����|�m;9�A�c���q��d�ۆ������^mx�V���4b��'��O/��O<�������x��<�n>�]t�L���<�Z��G��-��j���S��_m�x����W�^��E�t<�'���ł4Bz�z�-Ɗ���~Pы��}�P�!1sO��-h����վ�WA����wz�xk9ˋ5����-��
��=���2#�r:�H� ��C�SȎΘ]w��c�$�T�����-����2b�#�O�_I�d�Ҡ,�O0Ζ��;/סLb�ō~���~Do7��x�R�ٸ4	�ͩ�0	И�!k/xD�Rb{��Ίm 3U�E>۶H5�Gm~����9@i��G���� u�͋�� �����侂
�_ BA��ohƜ��.�9P�v���B���a!���h��E4-w<	6�����F�V/�r:�?{x�Z>�a�t4��Bs�c�%e�*ww}����y�*>�C���YsJ��?�\9�5��"���ʺ���姀�]���7T��w���?�s��`2���U���V7Hhf��<�VΘ�:�����!�n:��^��n�Np��9c.���Ϸ1 �2�X0�7�7�Ь�XJ�}�Q�Y5�χ��[�T�jܥ����U����_�ks��k�?C��pDGWF�5�T�*���[�!eF�0T��{����� L�����ހHDkd��u�s���s�o�PbQ%C�2�}��O�����/��,.XHc�+��������_�p�z����70rR>�W��I��p��p�/�C�3ه�)2Qv�f~�9�ɭ��#���83�2�
��3~��D/N�*s��e
�����a�/h��@T���mg���wڄ%X߹������(@��L��`�5B�z�%	���KG�E�|�$q[F,vZFCdF&H����l߅ �;7=�l�\/T ��PЎQ	�{m��@JV�w��"G�p�ۮ��]Z��j|�W��ъ'��m (��]�G;H��2����D$hj�>����Eܗ=����+�/L<f�ct��T�D�GlW�ѕA����ס���Ն��!��E�&_lKF�u|G��8j�|˖X�Zt��&yGE�Q�G���yB�n���l�@�nބ��O�[v�hP+�E��)�I�D���a�g譂G�=S�xE�}�&�H3��J%�O��*���]��\k�Y�o��6np&͟@�\?*L�&�)8���E�RG����a�2X�>/(��2:�	)��|G>o3;	z���8�KlvF?�A�T�k���/���jI܏�]���x��p�׼Z3����U��<�M|#�~�mV�.��	{`�쮊�iӇh!K9�����y�X���%�Ϛ��+�1g�5!%2�,S��s�Kd�_c_��>OHK�:6����`v����|�h�F�e}�����}�횙88�"q����zw���Gd����g��	!�p�"��w��"��@k�(��p�m�=::�=j�'"�^�M<M��\\�����&i�"v�K�̌g�`x6��l���*+2+ƾ�͘ʵ����l���^W[݈/#+z^��dN*�/�1.�M����?(����l��DD�i9��I��j~r��.D���!n�#�N>�����P�o�nTC�n��1�k���WPU�OI�z��x�F����U/�c��/��	<ÍT��ւN`��{���2�=_�������^���<(G缈s\.wN�zw����L/5�i��5:����V/dΙ(�ƈXo?�1q�o�=;�����6��=���j��������r[',���-�c��'w��9��_05
m4�'�D�է��6��6v�U:�!���K��Пջ
*[��q,�3��0��*D�q~����V�QU`� ��\z5sD�0i���t�ș��������M��uj<d�Z�d���]rL>>�:j���0��(V�/,��ܥJ�yc#BM*�MA�#'��+�;0�6���[��l$`u1Jdz��2���d'��T����3��~�3�9Ӻ�޲M{��;y������:�C��%����6y0US�H}P��9S����m�����������L��c�贛���n�r��~�j���u7d_(�Τuq8R�c�[J7�#����+0���S�K�ĒtG��@7��K;k��Θ�Kjxc2�sQ�^=^3��q �4���e�-�>����/{�<��H��<�؊��q<Czg�H��9�2?��m�E#�R)�V=qN����T�4#���|�m�M���2�׳f��u�Xr�ַ�F��Q�Ƥٺ%�?^N���[�鄓�^��"�w��^���{R��P�mi?b���"f��+W,TR�M�-Iyko��#8�q�ܓ�{X,�g2�cE�O��ԥ�����hl�,$���*8l�[����~�B+��h�����ᖖh�#�Ass��Åjd9Z���\�VyTN����Ok$�ǎ�?��hd@��6�c%��%�K��cKS4g��M���_��x�AM�������y%%U
o��~yw����'בy���p�jF�����-b����毗=1��%ԟ��4�k����sJg�X��i������ͷ��@\���e�����Eh{(��/�X�9%�#a�a��i5Aɗ{.�M[���U����4���gB�O>[	�t���\�
�4��r ԑb}ހd��o�2����g�Ś�u1��ؗ��$B̜WI��.��
�u�2�<��E�tw�������XonX���Pe��a?vB��k��2����\��ꡃѪ]���<-�6]�8e߿�-ʺ	6&N�[��q
ۃS�b 鋅~K��bޢ�=�> �ݵ�Z���~JD�KjjAG��{��6�|�d�i�*p{���g��
h�E�_�a頬�/�2�(vl��������߾��X�:�W�r���ү�^k)���H(��bu��k��5je�Z�\e�zsX�,e�O�nѣz�}dݼ����4�1|��t�ǩ��~B�&u|���/��_��J��,��~W�6�՘�M	*TP�W��Hw~��%T�FDw�#gt�� =F�כ*�>��2�l�_o�F� ���~��ʏX���w�I�����SA�
���u\�����}��hB���˶�sh/�	������kF,CpT���9���xB��� e��X-��r3�go*z�nN�Kq�)�ѧ�}� �?Oܳ�Nu�`d����u��J?��!�eaz=VnPQ0(������i7?@�!���%noJ�܌��e�yk(:��`\���9�d���r��-�����i�.eޘ���	THS��qx�kX�����2�im$�LƦLý!��ݙ
hm4�G�r�X�>��TJ�k�.�l^���D������Q�2W����nN1�wj��ё�]�>2-^1|�l��W���$Z��6RP�8戮��Y�
��2���Zǉ_�I��8�b�s�|�yj�~.�	<wH�SڱϞxd_�9we�A�9@�9�$찑�ʤ ~uA�:��V�����.[��Ꞔ������Q�4u���gXt��`�uE�|�v�sy�>��l��NNaBT9훾Xf]j�h���dߛ�J�%W�LoYq�QL��6����M��V��7��O/܇�R�9�6�B��#�)`ErL~B�ґ^8rێ:�̿e�5���Gͤ��u�h�*.�6
y�V_t�P�TG��Y73w�����hM5���2|H��$�Q��W 56���t��ڀ�jȔ�,RY�J_q�����1�즿�����l�ighZ��H139�`�����ԈVQ'SYq�h��5Nn����k���e��Aj��ҳ���)�����p���[Z_��p:��Sų�a?�w�@!xѯ�~x@�xA'vw[��f}�Z�W��6�2��=��5*����TIpn/��_8I���ZI��LiPJ[y-�����x��|W��\���\�H|�KD�9��yc�+g�t�� J��Zv�V؆qW��y����-�{N��5���B����N�{Y����a��>��=�����l�^�R�� WS�����Z��a'�"Y�U�����Un"G����5V(\��0*"��{h���[�^�ֳ`ꜫ��'S�/PCy)<W�9�O��
��p���!z �8<�A.�q%>�D	2U�H�{_/ �������1��uU|7�H���W������][CD��������_X�~ӽ(���VL���hڹo;��t��%bs��ْɚ/��{�8��?�y�׷��2=�`��r����, ���M�'R姹�;����O*�2�K�5�����T����bSM����o#��[5����3qɌΉ��j�-�-�9��ֹ9P�Ef�BMҧ5�����hfJ�?&�p��ï0j@_�&�=�˺z�\	�U�����i�b���)=͍��<�a����ӆ�&fyw��<�������:�j[�8��%
�W�aJi�}�]W"S�/�#I{�1�w
���H��i�#X�36(Q��5�g��;��MS��S�.��[�i��^�17>�*�W�q�pz��'���2����O�J��򴴟��9���߯��W��1Rp�_~�e��Y�/����b�/UUq�<V[r��~�J�]|�A�7�����r��s��x��w W2v�N�OZ�������"H�#c��9^����'ph{��`�u�2pk��s����v��*[L�|h����C?��S�.��
���Jf�L����L�w����1��_�\e�t���Y�XU&�pkA�O��;))8��)(i�LBg>ǟ��*v(CE�Ӈ�P%��i�F��⁁�v0Bvyy��� V(/"@���v6����q��;"3�J椗�F>,�M�SغQ�c��3�dӈ��a��9��x�}!�0�镣��C�"9%/L�n@�+�!Z�s�È�Ǿĭ4n�}R�c���Q��ĥ���ޗp�R���Αډ��J����X�P�N
��B������m��<�>��:ZZDttt2}ԟ��nz�2��Ne�|��'Wn$�%�勑%'ߋȫvg��,c�'�!�n:�,^���X����r�)�I(,q����b꩏ÞT���������[_)"�":ucߣP��E����B�دǐ�6G��ˇ��N-�l�*�I�E8;;OJ�S��8����������y�?�����)�Y02�P�]�
�����u���1B^��m��}��k�NWz.E�:j�~m��@^>+s[uS�oii���D�z��p�̈V��r��VY������w6��i-:F.�"���@ծ04��!�@e�W��%������*��6��M����3�?���~�z��rC�|�<zws˖.���N�]�}$���X�sCt@�n�@�y��� �����ku���_��]q@�E����!Q��6�k��s¤|�B�*y����~^�R�'�/OmΘK���
u��*�z�I��J��r���F#���>K�|8�b�/�����f�����C>~�dSW�8�ع���N������5�9�:j�_L�l6��RB����k,������[�x͚ۏ��`��9\'ؿ�jT@���ԴM�D�rʄ����^��mM�\�VL�w˖:�59s�'�C,���U\��7�?������ZX��\(��{b�DYT	�^�6��5�=���Xu,���%�ԉ�2)(������ɥ��*�i\4df���'��<<�(4$y,E	O��Ж�@�7A����z>���M��ү�*ӷ�aG31o��z����� �u>P�gh�0A)?�P��<:�'.���'��˻_�vf�� MG?`r�%�ٲ�ܔ�ebL���I�rJz����!�g�_$}M�s$� S�:�u>3��ψ	���<�qo���+�5m��4�{c$,��861��|���)򠸵�g���p����C���Tܾ"��1Q�J��B݋���R�+��װ��C<?�_C� 3���%���է�:�v��I��ݻ��0&���R)_����@�I~3�pN�r��2�n��Q����VR�#B,2�������WZ:M`���g�+j�NtT���p�3??����ۿ�Y�Ͳ�S������(�Rso�h�2��}��x���\��B�%���~�o8ѿ�s�F�o�o0p�8��DP�K�;'ocJ��lҶD�p#à1ݱ����s����5��\tt0a2�hȄ�8��y���eT2�,����A�P.�C8�I&J����j9:j�{�@g[8�����Wg�a��֛@-"gg��.�T��H��a��s�h����,+�,w=i��>��v����� �`�w��{aCn�|�>��!X$��j�R�^_�e~inn>�f?�0�=�Z1���$�[ɸh[6
��jP��@�����S4��):^,��5������T�[�(8f�:&�4:o��ɜ�G�������8��l���������\�j������󆝰�A�L�?U'bu�!�>��H���)-�7J^mo�S�0�n;��8����F������׏�������3���S@�����HS����b���2�r'�V���69�����ʯ����խ��4��,�lI��0�q;����e��,#��v��z�ؚ���U=���VH�1��>�JBӨ�E9"�1���O�1uj��ɛ�^��ĉn:� `v�|di���(|�������'_�o͔� �T�|e�@{�LY)oI=����B͹NN�u���ޒ�������4��w<���������������2�@�I�+!T�������C�w���=���ze�h2#�X��,�F�݅�-���Q�.��D��H�ׯ7��m���7�/��eS�L�,����]��/(��� �|�|�E���+�w�J��������v������P�<���_�]�~�/��s��5��x�7m:i�P�P��\Z~s`�#`��F�N6��c9<�nn0�%�ܑ?�{ak��Q{��_�*:�9���m�X4$e̚�H5��fHf��g�ΘŲ`�U�-�.`�!�v�ɓ�Ց=�����������޵���AB��E������������_�ޟll���)jhh,,����bL�b�X�:����8�u���@�^�e>�-sj_�g�.��cR��:���Z_?��,i|Y:{��?�������6��6~�`P�7W'j��hGZ��
�����;ao����B�_bW�����������v+���������k�p�,fo&��aї9�����%. ?����c[�-m��Fc�;��_�[މ��X;�R�����"�R�~���K���������}mov��v`s�@�J��9��oo��.����9��ʜ�>�"u�B���+�J6!u�+�w+����W�Sȷp>�<�JP��x
[��;�jK���Z���2(���}�$V��S���)��f~��^�n����ɸ���3�=��bQ�^��>�qb�� �bjF۫P D�k�6��kZ�<
ٕ.D�5cvC=�����d�/"�}Y�����[Qɔ8͆88�r�XI���U|&�2�1,�RP�����
�>��i>�#E.��؀���z�ʧM�U�~.��K;)RJ���1����b�ڏ,���qνec\�c���n���P3&�1�Ҝ���\�2�j�%pJb_�u�{M@�ʔ*�������4Y=�<�?��4���y	b��5�������H�<�p�|H�s�|��v��D�wvt��� �j�ϴ�f�� ?�_ҲI`��U,q����﬌R�UN����?�o�s�|"T�C�i�\Y�w	��V�81�n&Bٔ2��5�6��	R��9��Ÿ@����`��G��5��ŵ1`#�d��h�K{Z�fA����V�Dr`ܙ��c�T����OJc����a4�Xm�fƽ�r9��y�*>́+����g�&�g�uǳ���#+i&&YǃqcUs�@��S�\�"U�s���7���&[r�o���@� � p�2�/�ӛZ��������h��/�"��վ�M�ٍ�@�r0y|D�۽r[2Lv-rQP��#G.YQ�������ߺ� "�s���o5c6��~�"A�O��Ȧ�qQ�������tqU�_SJg���PsF]C��I>�k=�2L�D��0��K�'�b+3׃�\�nT������P��-n�7�b����E"[�(2�Rc�K/w�?K���c8L��@�����}4�8�e����3Hz}�+�֭!�� ��Ds�����©;z;��SĠ(f�`�]+WlƎ��H��G0�
T;Rm�hr� �g薉d����0����K0�蘧�$J�:�@4o�bnC��?K0U�FoV���M��@����~�9#M�?��̄Eβ����'|l��M����	w�9����{� ̰���OJN�����$1]�THg�)U
�?7�6p;W6�F����`�+b�g�r�ǭ-aeUȏ����KWg�!Xh*�fy+�&���|���{3ڹ�zΥ�*B6����4*ս���k��'����	�˅��/�BeN�fҿ�ɣ�3�4H�D�Y�| u����$M� �������wk��]����$G`g�����0�(F��Px��p���@n�>TaÖ3�P/��ɡ�d�^���6�����_ƕ�_y���G�3��� r�C��,|ϛ��w	��b8YI�Z
$"Q��'^7�X�s��Cy�	.�,��)ۭ�m�Y�$ޤ���'�(��]v��=��\��?�x�h���b�osSKwR�[z��$�������������Q]��sZ�^�E&�<��=c3E���ʟ�&��~��o+�ZZ�39�[�6r
�tDD�>���oֵvE:�y+bf5����}^}�a������/7g9�ƕA��n|O�|90����r3ʈ"��ϝ�CP�՘��q�3��w�y�F�՗�x9M?��v�6H�O��N���Z^�Ϙ0��*+%�Z�`*��K���P<�C�:�7.�;��lĤ�Y�Om��1�O���ED0�N{=�m,��u��k�7�ρ;��__���
p�#!�t�����Q#�2㖘�C��"{����_���JO�u{�9x�ɤ�a�����W ��5����Cp�Cp������ݗ���K�]���	�o7��^=��������眾�}�)���<-V���C�p�R�0��`3����g@��g�,"��/�H8�����$�J������(���He�Y�nv�"\�8e��,{e�5d{����7�I���
4�n��@�����Z���w�sҺ���_�؄���I�һa��I���5�l@:������?�6����I6�߄O�����.R���7��fbS~-�f`C���do����k%t�DR�0y�f�r���@\H}�N�KB|�rv`n3N.)��gf�q�˰S"�;��?�.Z���#��r?gB��:�.��_���w~�*!Ŗ+^r���l4B�{��0�Q�Bݞ�Ľ��m����gƯ��b��w�|̇3W�Rm�9n�lW>�F�!*�w�&~��}�ڨX����f� ���h�q��?T`�LOǇ�e<[����o7�LW.�����������nñ�*lL�Ӳ�˽��Ł�/	�p6��p`��z&�7����y��k	�E� �A�<�FƟ$�Hї ��(��+��B��B{�!�ş�33A�ӵN/���)���%Z9 � �5���iݘ����R��kU��I!��Uӳ 27-Y�����5��KO���ޚ��\�UV���׋�#�3����J<��3w��Y�+2p�#��%Pr�5�چ!��vKO|�8��֧�6l�;�ZlF�Tr���fI�	[�B&g��!^FW{��d��罐R\s@噬C��뗆Dga�:I)�,j��)	��;'������rw~��+d��g:�(�1�����7l�|?���jo����cc�ǹ/�J����r=�w5�%�N�DW�nȺ�������PY�7(7SGkʡ�l�c���K	a;�!�`S1hw��m�*c�0ºI�J:\i�u$g�x�E�Z� �r2�#^]HwUgQ|:���!e�Z�p�3��q`Rc
�3pV���)^X�рb����f��?f
z���ڎ�5��w��*����8q��u���m��Ib$�niiD; p�]՗���|t� Ff[-ߖ�lX��4����?���CY['���>:��ӵa�@Q�_.�35y���B���g�L�(log���oJ��{�w̨w�$*��ʐ�n�PW4)IV�f�V����_'w[�����m,��V�>�p�l����D���J:R���W���7�B<$v�/b;�>���~���Х}��W���o#���5j�/��N��Q�2\�`Zx�����r �'Ț��AN)4> S۰����YfYa��MRc��t�ZbTV�S�}�h}�a(�e�~ȡ���)����ř?�CU��!a�8��H�,�]��2�֨�����qa�9���K2�D�m�:�t/R3ݛe����"��:m`����
��_-�g���Y$�����Α��bv��R7;>uc��� �7@����U\k�>��ў8���Z�;ߴIh�r�%���A������-?L���;j,/,�V�E�'��ӕܨ2=~��h'+��g�Nl�?l��>�7�ܱ��W�P�DCC��;B�<��r�����4��hDJ���>1_~�5hM�]k`-H�m�΁�	��VS��cI(���	�� ��I�f��W^���)��G�_J���g�ڽy|������� t�z"I���{�����p�����I��t%D+���ҡ����O�}�7�o8���A#iK�6�C���*�\��&���吖����Ď$�����OeC�O���|au��sc�\)�a,OGL����m4_W	9�,�ޥQ����Bj�r}��e�"Q��;(��o-���|+��Z�c�����%��O��YX�Z|?97X�t�a�}�>1u���R�xk~�4�ޔ��)t`�Y}JCy���X4#�k���i��_�Y��0R��e�״�4��Z�!J$/���6�L+��n�:�o6 VB��!�(J�P�Ł��)ѿ�:��ąg�`���Q�"�0��G+Ni�h�zl�S�!�%Ov���5,��ŊC��P*��uo��]�<���!�Ǘ8�V�����6#��]]K����c ���Ku�^�'��ٙ�n������^�R�ꏇ���3�%��E�tv�B�Yr>��Q�Br��
x�`��9ܪd=��JTdHj�/��c�������v��t�P��ׁ�u�۱���!o��eN��--5��V�[zMw��QS����K�w,���I�O�IO��_�W1XN�K��t�^�U�Ώֽ���*�]������L����b#c�����v�fyb��ٟ�2�:�4���f����X�=Z�������@
�,������(#�]��c�^`�zR��`����7���QL8�U\PŷN��!n���O*��Y�>�}H��z�I*��=< �����-?k��$��x�/����]���O���s6�J���L?E���8��
���? ����wƺ�cO�5��gLNB0��,(���	�ׯJ9H'�i�w��0�#�>.�#�%Hn�n����|Oօ����#��啿�/�����~�k�X�>����z�����h�<:r5��ǩ����~�h���+N��+��ǘ�!�qcI�:܉䤏�a�4	����V�4c���C�;�G����y�!���X��y��{g��<���|k�U����A���,����ȞVD��s#��A~�,������>�j/�\��Y���2��OtG�ዧ&�>Gse�{Y�NGe?��e���@	�����Uu���i�LF��v�9.�B +sVY�lR䉅N9����h�!�G?�7H�P�=L8:Y>�^-�ZW�,v��е�8S�I����깛��[�����'Bt���Fi4��כ�U92���f���Rdu�7@!Ô\ta�?�q��G��w8��<9I8ć�ꑰ�l?:IB
�=��΂QX��0�����N)t�����j����27R�-͛0�I�c��;�M����,���s�#y#�R�.�C��&��r����&������c�?]����mѽ&twE)Z�"�(�g�9mCT4P`^��h�5�/����ZM�Z��-��E?'Ӥ�^��%��dt�M��N(�|i�q&=�i�$V�fd8����_��:]�ȉ�},!��hf0Q�	�|/��S�w�ǡ%m� �@	���qxtr�ޝs�J �+Bvu�rc�*����q��[c���6$��EMY���@0�����0����/w[j�y!j�|d�r�2∌�Ƅ��F"K�DQ��_��+S����V�pF\A`��	���D���ջI�T������<`s�ͷ3�B$��w�:*#��O[҉/>�ŪYf)`֏�j�\�T~�1QQ�G�����f��o/�W��+
�p>��[��m�<k����x�L� ���)��␠�^e��C�V�u?��\�k�D��t�pe+�\�����*y0�W�c��3�������"���i�d�R�~�������+�1!ŗ�grY�K�:�BU�Q�Ws��2��G4c�N~S�L5��[��($���+��N��Q��R���m ��x��f/s�;�O\<���h���n����#��� ?���eտ�`�JPs��ԗ�tp~X?�ܰ��,c0��K0��!�� zˀK]��+JĎW�|�b�ss�2o 2ڧ/C^�](.]��Ѭ޹ɢ��ӂW���u�0=��l[��Og��wv^�8���`�Qv�؟���\`��UCzP�Ҍ��r���r�#�k��H3���9����2E��'~k�@W%�SLS�}ZᦑV"`��6ZS�u!��ߠ��*�f=�������~'�
�A�@)�k�F�}��k�{���؋f�}�H^~v��U$�ѺN��D#[A5��5�Q3��C��q��wgt�v��o9u��>��=-E�/Hg9�u���.�bش�fE.�K�!��ŀ|8-b�7�X�9�j}�˖�������"���*�EG�؅�������2L���ˆ���߆"U?�%�����ᬥ4�Q��/��rPR�qq1-�W��I�y��TxY�p�����6⚧#���l�k?��T|�nk����P`�]D�2u{���Y8D�d+a�i&k���F3D��T��'����	��.w���FB0gJ���j�
��2��.��*E��G�\��(o4�*U�z^o�>�Q�����
����O��K��6}�ڳ��9�Dl� �2��󅩹U���0½�4�Vces�5NgY����T�Z�ttML51%\�Q�nRe�KXbᛤD��x�s��'��q7G�,���t��3�ճ� ɋ�=��PB̩Z��Ω]��=՝|��ԭ��T�������Iq���!4ԙ��2d�0c�-'H�w_�M��Kc�wsh��cZA�E3(
�J�)�0J�h}����5�`#8ӑ�M��"�^�|����t�x�ǋ}��b��Qk_?������055�}��}���=��^)��y~�1�jYQ��U�P�r{����KKu:]%>���n"S��ݤ�HN�-|����1ٟB�����ܵ	��gXHG���i�|�<4
�~��u��iA�o׿�2�#���ޞDy)��t���Y��!���62D��?l��o��)�� �Ռl�ܔ�Z9!s �qZY܉�V�|��eL�u���EIw�v���姵�m���� �F�-���X`�ky��+��]UK�_��/} ����o��/��8�gEo�'�vP8��sGt�!�?�I٭^�?>!w�co�ih\v�.������9�����$��#��f�Њ�0 ��%�1'a+�*��]��"��W
����IyM]�I	9���c^�y����EE�J���������33"������~��@R,�,�۝��`��U�jD懗�h֘��9�v(�Ҽ}#?
Ӽ��#�7Uţۥq���z1�5��ֶ|��o@�	���X�ZZF���I�Y�Ʈa3ӈ�غ��o�#� �����J���n|K�O���?m/�X�����y�|��s?�x���;�aҌ8��d�S�ݭ>��Jt���,F8%p�
��=ɟK�aխ�Z����jT��`�n��r�pn��/�κG�΋���qޅ�г���3eBV,��ֻ� ѺWɝ������0c���3�����ď3|���鯛�v�W���Ъ���GCN<X���k��{q�##�4;������}�e9@T-SGI��;��?�V�Q�|���|��og�G �Q����ew���~�=/���X�hx�o�O�lT��N��ۅB��`fј�0��Pղ�Y�=�Z����^9C��t�LߙZA+
k+Ԥ��`�yY�B��[��-.<+`��D>l�e��N�<Rl7ٴ$7�<[�"�O���t�Djc)`$/�'���4I!�%,>~]�Ce;���6�QU���(X��(7��T�\!N`�U_~Q��������3c��W9��!��6���*fI�4�7�>��n��X�����>.�:|��)��������.��W���.n�w�z�|\���`�i
�|ҫ�dA�����0t	^$���_N��l�d����@^ir<�װS�E�(��4�4��9�w����s�_��:(��b"
b6/�_uUF�^\z�珮���[���A��]b	gH�.4}po��ܪ���n�}�k��m������0�5�����s"�:=�N1�6,�Ҿ�`�v�g4�y��yl�N����_!�,�s
���3͖��S�	X�۳�����5�����ι�uo��[���ƥ�՜[�Nn2��.����EV��_��C9�Ɨ��H�D�Z�LL�'o�d��nd��O�_p�w��bS�r��}R�4�7FE�e�{��Sb��ik��6�\k�.��*oC�������
�&�g��������.���N"6�G߃��jy��qk
-��fw�?(��P�� 0(�u5�k��iw�,��D�꯰Q��5<e��I,�Y��6��<z�@�A�LUM-��j{�đņ��൘e�Q^�</��\2�a-E�a_
u�&��0�B_ߏ�@x	*���3ysSy,	#RM����/�`���BKl��+\�t��
��{1�&5[$�z��ye�l�:]���2�vp$�Q�O��0�}��'��б���6Gǽ���~���ʇ����qM�o>P��F-!p�Y�W�H��`�n��'����ΐ�1���6����A0�~�H�I!N�uҨ����
�YQ�򡘜V++���UV�k��շ
�&+����� ��$�[������&��(X���U���Eu��B�IL�O�d���j�PC\XQ�j�I9|��&�l�*L��Z���n��ZN�j������
�rՖ+iH���w�6Y�a��ly�ȹr��A�8*����]���E��h:��K�H$����u��Ch���(-�]��R������D�N:��*QN��s)Rݻ���%�l(x�ߟ)��wvB��A?c�2d�do��u�::��qs�0����Ǭ�~����&�Ƅ�3�n���[0�^�:�_�IN�X/aw���y�#���Wn����f�S.�Jެ�'5�������\f���wG�'��y��q�X��oOM���Q�����,�����N=pE�Br�~�n
]b>b8�i����s~糷G�'o��b��o���^��Ja�&Y�=�k]^̾�{�@�("'��˭z"ڭ��ߚH�Ρ��ɥ�sQV�i�����q'��}�$��[���ף���TD���c�z���}p7�Y4 {BԜ��o�v��~���g�����VJ��W%��jߠg\e�Mx��)�����"�RA��< m���@J�f�A��h ��W�ZXV��(�"|F��F��B�H�9r-AD��
꓁A� �����R�>�vb ��b�(j-=����޴���}yFp��N��d��s��M[%v�ַ72DjPbON��)k�DT����,E�H��=�8^�t���?�R��� eQ.��/�eN��N"f�����2��+���E1��#���'�H轤ω,�*uJ��Y�*b��p��vu�3���Y��Gfꉽw���n�0�[#�8'vs�����}�ý�H�` ��m
l�:�S�W�.o�	ѷg"c^��4�H�D�T�d��ѕ��$��ͷ$��H;�A��������M8�4zH�K��g�m��1 _�u�{�)y$ǜP��q(k�5����l#�V����y����H�́1����V�����@��@�|�&��m�w� �����6�;��m2[0���B�5@nln&~�Ɣt!=:�-�`M�H5��16���ףF�2����]#�hƑ�iu����588���XJ�WN�w�gνʉe{���E���@ �9
�&�\MC	����PCn��r��J�j�B��j���zL�����[�(Ur���)3Wp��R���u;>Q&c(U�(�w�.F"(�{
��.SSTt�9��������^�e��P�O��Ӹs������ޞI<��#B���QZH*�j����$�
8�,öe#L�R�9�%KKP��	|?rJ̈� '�ٮxgN~��p�]�X|O\e�ǹ�p}�j�W�}���:T�QZ�%��uQ�}�(��!-Qq{/����eMǰ&�z�-]�e������8�X�ˌ�|��`�<��(�jf���^$i��#!�����Ʀ7��^�ˮ)���e�:��bBPwwt�	��7�Qv����*0��"0n�&#(L����N1]CbL����bTV�}�f�I0�}�R�0�3܊�P~�EG%��R�:x$UT�G+��ܞ�ɪ%�l�i'X���U+�,�21�Ƒw�ߖ�T�X��L��3��%I���aq�"Վ��UR������͐>:��:�t1��~���k<l�&��.h.0h��,i~��#��N�4�Ir�ΖZy�671J��A6j����H���n�4���և��}���Yjp0t�^:�i�K��&��L㧬��i���Ox̪Rh�Q �.�.|6(> W�p��hG���=C��#����@mx�5'I��>ё���9�a����ݟz���q����Y@$��p����چԣ$5��1�z�z�}#n>��i�@UC&W�RQJ`� ��#�E8�����&!���	��������	�.Q�qr
�z�{�������L7�}�?�ǂ�@@�9X
�����s�h��JgՏV��X�����M�'�#�'�9{��ju֚C�!I,,[�{s2P������Ć�U�X�̉��+���
���Oϕ/wRP�����Q�_��*8S�BS�U��b���P86��� w���$��'Ȍ{�c7����⪨XQHu��7�o����C,������J8�ǔ��?���VG5ے����0�LM���}D�?#R[k�A�'�-ނ��E�����G��72ӥQ�̇�?���Jl
cj�i�ƨ��m=����8�q��@'�[���~v��	6��n����C��p���$�ؔ��|���ӣ�����] -��ڊĞ;ؖ��l���.�HtCҸ<R�4Wa=4@*_P��Fm�Q��v&��SK�I$�zg�P^�n"����m��r <�h�"v���/�`KwBũ�ՌTfw-��wҊ)�~�߼��W+���$�+cq��ޑ|������;~����g�{��}]3۬�#h�'��w��s{���)�����8 #�R�
�t�WW��vQ9�x�¤)`��$v�mL8�{g�$![��{� X墲)�QTS�9�~��צ�`����T�lgDϏ���AF�0��
ط���k��c6�{���`�����������/���.|9J�4�r���Fb�I�Me�%:���0����r#�])��������F�{V�����âGӭ�5�V��;hk9Y��hnۦ��E��!�g�,��>�o�2��Fʯ�G�>k�:�t��Nnմ�L�[P�]��3ɸ���a�p��߮Tօ�$�q� ճh?��+i8ڟ(����$PL��G�_{�^�i2~���(��G��Hw1��S��ف�M��6�G$T����b��#$ 0�n>�+͒Z�c�:aݺߚZ�+�{�(D�u��|U��YF$HO��TEQGR�.kE*�+n�f
ڟ�t�;]��h���,ڡG!�3�\�.����dn���;�<�֫	�:�'��}q��߼<a	�Ka AQq}5|�&ܰ)M��H��DݻS[A� �:���Y塕&�/���̀�o�������?�Z#�W�ۍ���|�����eO���?�$r�M:m���"R[;I���0Y�\�B'��$9Am"Q�m�'h",fԥLA�:��D�δ
e�/��� ٌ���.g;�T�q%W�OU'�O}�8��.�c�yn�����/�13y6B��CU�Xi5��#m ^�@� ��㶄����O(����J|�iWL�c�ۦ������������p����w��Nz���1�K�����E=��}jJ�ǳI+�f�P=F��ix{j�n��
��*��~V�KFІ���Z��뿺�c 7����^"(y�0�r}g�UGz`�����Nvu%�x.��a�����p{���6�>8:2>�~����8n԰��ķ�����g�5��! p���������v��Sk�z�/_AӦ�(znQ�� ��t,؄Mx�ݧV]��p��K����p�_��qҍUT�7��Fj��0XF7 lߓo]��r(�3Y_ޝ¹�n�l�(�o��چ��]�@�2Z���({rf`�2ع�[^|�'����O�וE�a7�c�K��k���@NzX�6Y��9_Z��!ߛ�:�ڙ��W�hy�$Í�y<�5������Q,������k�H��}I����DD��b������k�u�'_%$�S��P-!�G�] �WJ��~I�c�/���1=T�C���8�J�s�dℭԞҠ�v,W��<����Ϫ��e�����w���:��ᄢM�˗����s�rKI��C��Q����'	C�C�s[Z��AUϡp�Sx�S��Vh���!�.�:΃��:���-�8+�o����#�Je|�P���dl��ZH��m��� 3/�0�����m͏��y`�G�`�iz�!�KA����P�����<��"qC
��q�تP�6�'�8O.6+�t����]S��UI��XX�Γ�ڛLd.,'
j�j���E�R�t|���xN��kB7Fq������MQJ���dI�Cgc����~��k����o[5���AA��sZ�u��)���O�9�$J��P���A;��1��Tp��B&���0ݳݤ4��"�k��2�+(�&�2��Pc=�����A�	�wn������F�U��O���.YƳi��#�r(��/j�o/��r�6Y}6�Iμ�	�n����a�U�Sл��B��╨�&:�`�	 ��<kF�?ooo� (��d�J�<�lo`B�6���󆤽����g��"4<>ٰ���7���B�ͯ�v_�[-�F�|��u11s�Y�6N���B_�ⲇ������Kl&v��ˏO��F�/+0#����a�/��M��]�.6πgK1�`f�+������t��0f?�)��W���Ĝ��~+T���}k�ة��8�jB�`��2���9�N�Є<d��z�s��}�Q~+:u�5J�d���5�����-��r/�ۅJ1�\�[��0�*{>�_�M�������5�=|�i����~1���af�Br�(kX��̍��E��oѦO 8��Å���P�����Bm��(�������X�1�����������b�Ht��9�iE�\���:|�T6L-7R��_��^�,ry ��*��Y�����b���u�Щ4`n+���6j|�t5�ͦ>�6;���bz����������{m��Q&��H�z�7
8��bed������u��ԁ��l¥Kܥ^Tҷ�5�����(���	bB%�$�
�,j�3�z%v��Ln��:@���??�б��ڡ
�yP��)�ev{REG�T��a�]l`�`4�7�PzƋ�#��ԏ:�~h���df��w��~��S=	x��#�g�"ؘȖuH(#�c�P�q/�����@��3�	�c3� �q���gX|���%�6kZ�����Q��0������&	�����<dt�}t���y}�~ˆe�uy�Y�C�8]
�SΤ���_R���w8v�?!�(^�]Z5S�8V$�������[��q����!�@��Awjv9�(񕏦>R\r�P%��\�[8�mA��I*��У��K�A^_��+3�^����W���|쭟-��&x����z>��)�ŀ2�@���v!0 N����5�������C�[��J�Ou�:�o���H5���X8�Y2�'��]�L��~�{����j�Q�T)	�7����:�jXQe�K���YF�����m�+�kV�z~���tQ"2o��?�M5w��Z�.���~̞�{�H����ݎ^p�	�͇�>�$z߃���f�̓������<�@)s�/ vv�����B��8V]7������Vԯ<��D%�CA���%���X1�9�c(�՘����e�o��eLI�AnV �oʫ;4�G�.�?�Mn;�9�*�R��#�=何=<#�"�?>qpSȰ˫�j��(� &lr橡v#^�RW�]�����b�����Vح�Q��� 9d�A�����R���)6`m����Z��%kب��,
T	š��LT�(�KaCp�|�Ҵw�)t��;1�J:U�8�0<�S�R_��J�aD��o���q���:��U���)��#�4�Л#�E����E�x.��,%8u�S��7K��|�N�6fS��u\}�Ex��K�2h�ҳ��<܍%�=v�p���lli<W��u�p�
[h�"���+-a�;[%�������G�:�8
�~�n2R݋���T�Aq6�=���ȃ�?�I�|��믏�	�Y�:��%��!�fk����c�?�֐&�cf�-�5�-U%��1�d�iF�����fW�k��(�������\Y<���N(/g�[������'��W��; ����ּX����v��W��o%���<�yo��]g�V����R�Po��att��M;8 ��qEW��>h؆���r�����2m3w���C�zg9k�$U��.��6�R�f�`���~1c�E9ǌ��F��V��qKt�#j��iK�N&��Al�h��(��,��Bʝ'��^@��#�B�&&�o�?��W��jQ;D-]���8 ��N�iZԢ�w���Q�`�Fq�^Ծ����]<��3�S�����r
l�(����4f�i)��&+w���@��
2&5 m����)Rp�k+Lc|��(q�O���-B0�$����F��D�p��~^E	������x��|z��(�$db����r�F��AL�Zh������`E�v�`��.l�=*�ָ�ᐠcg�c�4��z�E4#/y�[��e��1�0cӲ}oH
�'g������N$a�p7Ζc.!�P0y��D:nѷ�SI�*j��-�G���n���|SbZ�iV�8a��P����9�CS��*rH]�~N'�>e��Nc���)�$� �`A��05��w��3�*+a�@�+̣e9�Tޓ����ͷ��8|Z�pc� ���6~�W�(�0����U碩Gg��[�875�G�c���d�8�d4��{�>���܀N�\z��a%dd�Z���~���U��$���M�_@�u�~9So]oS��7�xXS�9�8�+��~���&���zp�w����Q�TK�����Y"HN����jI=��0�e�$�P�5��U�⽙�d숾R3`'�.k��~ �����d�b�����隍-���)	{R1S��D�x��^�%&�vf3���QBN�mHD��f�HB�߲�f����b�~�1^ �abbG��@x��l��r8xAB'
k+�?{�jR��<4�R�]�zR�i������0r��F�r�ǡL�f2h.�c�A�e{HF���o�F�ϥ�=7�q�g`���H#X�hG~��0D0qC(�f_x���Cu�H����-��*D�w�D`�ٰ&���,$�@d)�7m�j�5�l�kE�4f?������Jx���{?��Sw�y{����G��s/:��2�FDA�
U�9O�}�ĩQed�~"60n���IB��cq�'o��i	SR�S���'C~������/��� '"��� O��}�CIP�Ƃg}������p�5�=ݝ:���ה��%$�H	H�=��>+�����鉌<�i���A'8�0xi��A*TT��H�g�gl��i٩������D����}�ȯ2�o��{A��+Z$0K��� <�N`����;�hӷ�K�i�Q%�)�X�v?�O�D����6�k�	�����#��w��js�
�����ӆ���a��;#=��8u�r�Ʀ��7���ɸ��5	�%�X)�	ײ��`Z��;q�RI@j�.Z����,�����y��t��}E�����|"�u(��39�>.�����&��0�X~�IX��:^����\E���E���_nnn�
rK��h��Y7�&�3f�c�����DLcV.��!�`�h6�>��h�4����?���\���v�����Y�.(hv��3	Y�0�)M,g��L�_�Z3��B��8��Uܷ<�3�+(�3^^��������:�}%�~#�n� �K|�a�gэ�@I:�T��vgSֳ���t�D����w=J���R�'X\1v��l����_�u�Ng��Cʮ�̏��}z��;(���o���7�vҶZ�� ��9���h�S�z���/p���	�gfʯvZ �f
��뻦&������=�ôQ�·��-킟y�	-N���'��}�1_����z�/��}�_�'�w0�Z��b86GGF������0��n�d���4�?��4k����k=�;XY���������8bm��0l":�ݭ���X�)�ל��-��22];�z7Fw3I�������PͬϨ
����B��G�Ui�ǩ��Y��	��F�%�K��0>�M�Z�`/�?ru���y�����Z�z����N?�f�.r��܅!J�-�5�{�Xx�[��,�G36"�|��	~~�/��6��_�xx?��W##��sarS�������$D�����2�-�]6k"P(#�f�m��[�����0�=0��{���$����R�t��&&�>���։�H ���bu���i{?ʫ�Ӥ����l�3:ZI9鵠;�z�C4����~���Qs��.�&���@��Q�l�H.�yHC��%��& D/���	��P�?���:9 ����\Y�+˜6}oɡ�j�hZ@5	���m����J�# �{��?��wJ��%2,��#(��"\.��?�>��!��]�Gт2�f
M4���%q�H£�1qˤv�U,�&d�oiP�B���Z�Y���㛀�� �����>���tY��Of��q���>55���b�� 0�P|Yh|>�@?��\�j#R�_�L�7k��W>�J�8޴R+�w����+�{xNi�xB�JaL/>|�Io5��H2vz)U����MO�P�/6�7?g�Z��� �p��p�j���)V!	Rd fFp��?����w�����2v9�mD��D`EgǚP�^|�`''�+�\�N�x�٤���~H��n�C�*���q|_sy����VFFO���v������ب%.�rFLө莽]P`z��+��M:�Ɋ�˱�P���٬������]m����6���YN,nU*X�x�ؽ��]+�(�C΀���/��~��̂�k�ݣ1���cvn��!�FQ�e���`P]��C����5A�䈓�OӦ��(���(֧VcJ�>�
��nm�esA�Q�͍rt�ŵ��	�{ew�ljW�s�<��E�G��O������EyF27���j�v�b����
���	�EL���z^_��0vG3�������~�)Dk�T*�i1FF|�K����`�01��3�Z-��4�$4�3��x���W,�l�� �V����a�g�'g;RhE�5V���뫒 y�&������*���J�g��W�y=*����X(��Oo��G���X{a!J�ƹ�F������-0�Pnl�]p�9G�r�qc���&Q�[�������p�/vHG��@ο:��zN;`s\�R$��`f&(������U��	G�|������A�����sk�dH�T�Yѳ��h����l�B'R��͖�im`2��`_\'��ʊ1��˭䀱�fŠY�>l�����ߔ���F�����(�˔1������S�#H��ͤ*T�Ȼ ����d�j~N�����S ZkX�!?'t� �[U14Lh�]413�������7z��B�X�;����X?7�����&��z��Bm.2�Wr�[�.ΒV���zz��>�@W*�G��w��g"6M�r�a�i� �e�����7e��L�Bn��D���ʩֱ|��P��:q%���щ�N1�T���q���E�)~9/��o5�pm�p�Ϟ@�%���"N�+��8�a_��^���~u���Ѻ�S.kE�x��経� �h��Q�[W���U��ce$���m#*}��ߗ����`�-��%�"m��[s=���!<�b�[�OY9�E�R�!� ,s��  bH܀��!2�1��g�������jx��a��5r�1D_5��S���j��ìL\\܍x���m������әx�7��>_����][54����gE�o�7I�5�ꉢ�Z� /k
�a=Ůڰ$?J�{�(]��&� Hz���t�Ő��*ä�KC?�'B�����(b�DjL��'��!"iS��Ϥ�'*��3�2��X�U�@�Pbc�%t�u�)�Kw#�`N���IM�ZX]���˫|y�8��9[Qx�Ho�<\���P�sڐ�1C���������f���Q��Kp��� =�/r�v�A��,�Sڑ�!w�������|Y3v�f[ږ
��rX�\�h-�S8ևs�rD:9 ;����([]����hl3��̡�����nM�p�x�zo�v>����j#�R�W]�)m9��Db��	�sN��蕚��Q<�0.&6�GN�Ȳ�Ϥ�����Y*�
fh��DkcK�y	GG6�]�999�2�1X����G�~��L��+��Zt�������щ ���I.GGG� �f�7bC�t���*D�xޤ��L���/*���dѴ���<=���BCa"8|�ӂJ��YHt����5��x���O�e>w����lcp����)b�Fp�DKf�~D|db�4P�쓍�?7��4A���P�B&�~�#a�^�q�,@��䢊�f8 \`nn���ڽ��@ӎ�U;Y�E��6׫�b���h��%�hj��Gg0��__�X9-�Z�����kT8=_����I<�j��n[�a�����>E����lQ2��h���lV��H�=���Ÿ�]	\F�p0���G��=\;�Tت^T Y����r���ݯ���&�1@�K�����}���#��]�6��&|3�]4��2q�l�k`�FE���s�yH�&\��,��:�hli�l���m��!�-���ڮa��-!��Hw�� ��t#���ҍ�]��i��Mw~��z��C��Pֹ��sE���5�F�33��R�^�&�!�ٜ���o]��*B����I���V�B�u)��d^A%z���f���Jk�D��ν�SY��B�Td�r k��쎑Q�bx*��2��`��Z��v��8��_��BY�Թ���Z�p�2_K�=���{����G���d�o+��\����a*HK��zg˾VYLѴ�nD��3�
���'��=9����oo�oDJ��y�ϳ��}Lҳ���s�YAMB��[W���4l��ݶ�(�0?����W��%f�W �"''��X�����`<4d�勥ا�Թ@��Wʋ�s�����	ּmq��Q���*�G���ŶE9�[�{0�V���_�E!�y�YD�R�A���*�J;��m��rm^)5���H��ތXd*���]}Z�ԑ�9�/}ߗ��a==33���p��Mt6�Xaަ��6��?3�U6� ����$�-Sհ�*��KE����'撴�#N!Kb�gL��j����M���0�đ�m�ȋ��Ig���#W�@��nP�'��A��q�ۙSd�;݀Á5y�X��R�f����~���|I����=��$C���_9qJ����hMԼ���d�Ywi���84$�x��'6��I~{��"M���)��d3RR�ْF���%�����Ȗr���@���a�g�?�LP^|�%����K2�����K*#ww���Q���xm���U��p��p$;��Sp�z?|c�K�|_�^�d}}Q�Y��F��2���nw���R�Pa���a�/�K"ڽ'�]�5[_����>���uCT%[F�F�ݿ���f���3�i�|���F�����&?ur(HduY���2-��X&���(,����'�C'���Hl���O��W��I�-���(E=<��AUm\BWxF+,5\��b�
�[��)�FL����uk�͇�����9Q�2������5�s5��5�:5&��'�ĒVlT9��l�/p6\0��ب�Ă���(j-�1�-��c`��Ы��y�V��;&O`���[Q�r6��M�NQh�������*���@]����j�)�J�J\�����fx�_-(�Ωm���:p��[��Nn֮��e�^ł��;�}E���]�ll5�pr�`Mm�Q�Ɲ4K����vO�Q��a��=����Op��}tq�\��%R�?4-�2��f�7�*�����b[!zhhG%�7\�8�62ߓ���L����q��:OA�����ֱ֮2�v��훹�P��(��r`�}	5�7���<I��BC�l���9�Ρ
�e��zS�E{H�\^K�Ͳ+٣��!3��aһ{Y �s��QQW���mK���9*֨���)Tb��0�{���!NsɆG�T�?��Y���$êx�-N�
��À�NHKcH�j+VN?R=�o���B�Z���ұ�鸿�\~6{#vP�o��4B�#~�+ڽ�/�ʔ�T�?-��*#����{��?b/����+%����Mvӌc`Sly�Dh���xr~>��p�gY4VvX�l������A����D��"�O����������s����
CKY�|":4�N)k5���aq�ט�v�0�R���i�_�p��z{(����°������T*��h�C���:�ۿ-Ҹ�9�x]�ǂ�1�,��_�w�{�:(�Jٯ���W1�TC��AE�܉��l��!VA���0��yo�����SR<k�����P}��d�o/!��u�H +=��r�5�Hݤj���V�|c�j��dD=Z��{��^�����K��G���S�~f馾,#LG��G�|CCJZ�1�"]�G����h=�W�����(����?�����Wl�����Y��q��8����%���$4u&��eml�>��^z��G��|��$W},���:}���ձ�9�zODA���>R��'��x��&�a�� y�0���-��}W�+�p��x��Y
�Yq�ڙ�	k��8�2{s�'�T�P;/�����ϖ<����7bF���5�Ι�fPU�wQ�g-��0���1$�u�gR(�-v���F���{sYD��U��6�hʓ�Uu9!��6lE�䲚 7�H�O�2�����[x�k�jDP����'f�������r�
�mw`�y5C�:�9�R��'K����L���
c=�\��R�O��n��N���^�&z�����7J�t�Г`�A�"�dq)|�o�Y�\M��Yt	XM�A����1ٜi��Q'otDvw�P��ʈ_Ζu#�y�.l�A���?t��!-�	d����"����KP*����w)�㜬��0�����``@�Z���5��_҅���S��Ư��ğ�\LX��H����+HR�b��
	�yA=V�XAH��pz���'������h���2�C �������L[���$*�Ac��B�Tє��J����ug4�l�(v}���y�D����1�T{����{�)��W+�����(����v�o�9j�ϖ;�����ch�`T\���.����Q�y��e~$'eP�Z���瞺�����w�bY�Q:S���
\�v%�T�sRW��g�^��GO�
 �3��Ⱦ�/��^��{dU4�#���g�z�ՈL|"qB[�7�^u�'17x�ј�dC�(]���c�cX���Th�R^���nF�v�rN)��6�q�����͝���Y�$|ߒ*o�`L����>���
X�~����j�5�	u��i�N���HY]p8�I9��?.��®�AA����k��H�P1��
��Ȁ���m˛����o��!�����h��)��tI�Ĳ"��E�6x����W��0�����G��EF����Ʌ�����s��%RQ�)!vW�&���:��-R��I�K*\�)��b�leM���sz�B�f(��,/�ײ� &�z���]��b����n؁/�l����մ|0��ڴϚ;�j�C��:����:���|�
#5�nh�������gZ�E��bU��$,��%�q4�+��F�/^�Ew ��|�B��4���uW��(�ę�ۧ��u���F�3dK|���oc7�/[$]�w���Fg�w!�v(D/�'�o�嵇��(۪+	[��$-CD�W��4]X>Y�h"v*♓;|uV�<�%��-�,�W�iJvv�5�)*��V��7�Q��'"� e) ӱn���tt���t(��ө� rc�Yϥ�����1�D7�ĉz k��v0�w{89�d������2����	+�$%�co��w1��WW,|=�����#�a�kL	
�Z�͉��@�._"xd{e�y��G߾)2�|��􇨼��Ak�c�gA~Hg0�nXs3?PjGBBB��%ةz������p�f�K������a������E>�z���\���Ѥ3�������G�)���3{nͥk��Hz{��TipDD���èV�o�l�x�`�&�M:�e�F6�u����)��Ed7��0����\#9E�X̔L�Gm�)Z]�N��3n=<*���m�1^|�U>�I��f�G�0��V�����~�}gTI6ߩ���}��ۚ��\61��<�=|=�H�0r�I��p5�2�6#FD�k���R�'͍ĵ��ROBBH������g��P��T��{?������%�GW��G�@�%/����8~�'�'ˣ0^��C����~����D���*��I��1q2��(ގ`�:��r���|i�LD��쫃���n͉V=GA>ը]~T�p�͖�dȸ47�E���� ��2�2�!8����!q������Kt�J�Ԁ�mKo�Y�*��|�O+E�`9W��yҊ@o����\䊍	���?2TeO�ДU��b��I�<���Qu�r�`
�]w��i�$��g���F|���ϔ��>E���WF���	��~�DQΤWXlPN�5
Y�A`�N�������Sa�� d��!��kj|�=n��ӻ1�|>l*�t;��H�9�1�pg#�4�r��'���ZHb�ecTmЭ�-�����M�,Z��ap\E���>�$K�~+Y��ѫ��'>(�񉶥�������I��r��L�.���$m��+��{��cΠ��ǝ6�J�����}��F�������v�N#�wz��/*%"���Y��1XIOOҬK�X��`�C�ݧ2�i4���:!���[n����h�	�؃ϒW�N��r�M�B�0ޣ�]%չ��p�`�|����8q<c�/[�P�_��ưP��~��7�u�A�#���q߃&ei�^�%?�@i��FN���������F8-�!uXS��<o_�#�>�]�cQ�E�r��������aHL�~���>_�
<������ W/��pԨ�h˴y� i�lon������꾫�Vv%�IҸR9i>�bF��G,�eפ����XE�S�������MJM[��6��%�����ֵ�X���>&sO���������3wJ������Z
����K����O��0�/TG��	Жؕ�R�D!�1+?M� M�QP}-�����,{���;<�f6�1�|Ԣ�2��C5���s���ۓ��÷�K�Bi�(*wͼ>2�_�����&8p�ս���ۨ��r��~�) svv�Ȫv뱔S㨫��΅6~�=l1�C��2��cͩ��`�vr����4��I[�Nx%���=@m�df�T�nhP��u�]��g�@z9ɵC�Rbe\��w�>�ٶ�?C)�m>X:H<�o�5c��ÌW�����ۂ��c�7���F����Gd	{�:� ��qy`x\�Ƈ�����yf�l��}s�x�{�lڥ}�}�}su�Q��KE��;�����+��������Du���f4�B�ѣ)��_M:ϩSK�2��F6s����p�dd۠Ў!��v���o�7~�H@��Gr�^�O/k��W�%L�~s��ߞ���WE�;��}_��ƴ �[W����+0�:K%4B�X6^�f�{�����#Ô	6nV%�W|}@�o�;Ψe��/#/�a���l�VE5����\���j�i��3OG�;���\6��S���j.2��u�_�/�����w��@�i�n�*Wc;��S�B��[E�X�����vwBlvw)��#&�Q�%��l���{��3{~��;�vE��۟УRNm��l��t���τ�~6,�~]c�{yA�5���؝�3���}3�՝���>����d��|�G�-
�! ��']sܪ�&��@!Ш*+��V�8����e��7vk�A�+$��F��&�H��<�mݠ�hE�W'��P	�n��ݻ˔�}UX�"�t����8�E�-���B5�M����O���g�@O_N�(P6��C�CyʥDX�y�^���
���v��!"u ����9��MOOM߷7�/7?P��G27f�F �p��Up@�sj��b���FB�h��.kEhܹ���dx;�t7<�4�����w6˞��Q��{.��Ĉ19����|\�:��E&��DL����>�=�S�p9�X3�+���8�1�ڍ���<ߞ�	~C��+D��֗�pz�$���x����ߎz�[��ټ�A:k�� pg{#��(o��6�E�CPUd��,�i`�u
zS*W��4v��_���˂���MT�&gf�ّ��X�9�3j�d�>�ܝ��l����%��	�Gy���x�6xG���혁O�q�u�ȫ[84�	�rrJ:q��Q��x@f��d�����	�$Wn����%ڎ)����S�^'�n��L��-+���:�)3�idE�!)˺n}Xn�4cM��4��di���)�	����.��� �-�ק��lv���^)�ڰ�_��$ �/�)]ۚ���VP ՐׅT�}���n0~ty5?�a�F�vye)��A&�o����N0Eq?�omoǡ| q�M��jXv!�fi�Aɟ��/��z7��&�~p����V5L���-�Fa}	�o���bɋ��18��S'�P�������k�׬��d`��*��I,�u$��<έ�]����e+��J���7�3k��J<��%r��X���p����$�e�⽢Z�6!ɉn9쬶��4]P�b�������7�h\V��q|��·=�D������x��y�ײ���;J@%�С�᭠�,ٸ���ڄN�c����9���țm�/��������N�i&w�i���`���gՖ�y��@��ƛ��á��?8��(�o5V�\5ҩI;%#㳇!��3���GF���}L<�a�q�G!��pE�'������,�D�%�I�z3Zw�hE���X�c#������0���l���#�D�:��BK3L|��!�DR��*|i*����71|��� i�VZ?�'S�Ղ�/V���� t��Y��E�ƚ��#���j$��$�V��2G��~�(g�����-�hU���Ig��������إ�C���_�)6G������o���+�-��p0��xYUx	�x�����XZk�U4@i�ڙvd�6z1�4Q�Y�����#ƐI�~���)9����o!ʭ���.)K�#4��%�_��
�w�H�/�P�,��@n�*���9������,�q������4\ ���S�©����k<x9+IˀґC���3jk���� ����pr�7��g��y�a���ݥ�o�g0�q Gd���u[Kl��*��8�,�q蔑�Q�T��ˍ\"��I;$�H���s���-A����@Ә�!��j�&��5`E���E�D�����_�)%ipp�F�!"0}"E|�3. �V����rp~_3p�C��TE%26e;[��7K����y�ڛw7IocW������C ��~v��J#V���_�W������YBV6~r�k������+����(�&K$#��-R��jNY[�pb)�r(� *�e���C^�zݲB��.�O��-T�::$ ��:������>�3�eYx�6xW��eV�������^�M:��MD��1Mp��e�7�;o/�@S�na74v%D��9����D��x*�P�L�S���l���S�~u3^M�1��Q���Կ)Q���v������sO��-��w��
�t�U[}�5�������:�kX�z#���s�{�&yj$����4b��b��ܴz�%��4�K�B�@�-Eķ���Zr�@KQ���҆��RD����N� U�y�e����z��]������}q�K=�DZ.?/9�VV�z��X&�~9�vۋ����@���0����-��^ �D��P������ɷ@O::Y��~b� �Έ<���oH�\M��HYk�� E�>w�z�"w�·k���LG.�LDL�Z>飦Me����,��|�~�!�5�a��2�- ^�o�ݿ)������������L�t�p-]�m�v��!�Bs*~x���O�PQl��CG�J(Mm�&�\��\�[���`}īt{C��	�;&�0R|�bWO����c0�htwk�PZ�T�\��P�P4��L���ח{q��'��z�њD�{��9hEXI���d��a�ex;��WM�5�`�̖�6�t�_so�j�[����H`T����ͺX�F����k)w�e>����tpѤ΄�(O�����+��]��ȴS�s$v��{�^�q+��uw�x�F�M:2R�"���S���k9x���Ǡ�z�c���%���5E�s�M����}D�n34������`$^U�4��1�(�P_��k�M/��b���!-���w'Xˢ���1�3Y�aĨf�<�p�d���c2Ǝ���"�e�`F�eI�i;��~��h7s$~��ar����e	2��I �55��v�^ <:5�:K�갔-��'AC��--r��D���
 51$� � �{�F˝��ů���s�z���t)Vn]\�����}fk��o��/pm3��VV�i܊��t;3\r��JP�W��u�dϧ���@C�԰�5r9�QNi��Z}r�k�r2��9����[���i�ZH���Ϻ�9~�n�c���c3	azϓ��B�-3og�������+�j�����>�}��g3�(�n�KoC=���ݴ�kn�a�z���V��%�w���5��|;�&����僋�$c��z�!��e�TOc�����7���G.�_Omu~���mm���B����"\�����T����-�WF`5ޤ��Q�=.���D2�~C{c�.�;���:��b�PJ�iE�g�C.�.��;�J�K<�|A��Sf|�To ��!9
r���S�A/��tI<&s�V���&���ӱ��B6]���="�g�J��<�@�iL6�iy`��M��
~m�"<,�V��f��Ygm ������M�����z`&g:
��$�����?�C����rc��ܓl���y��y�V�4�C��x^��m�|��h��1�sR���*!Uo��I5�kj" ����W_zy�	�
���v7�b�>�=�/�Du���+����T���ۿ���Ҭ��)���]����,���i�[)�_dQ�+� Z�T��ifό���ܖ�XE�����T��k,�c�ǿ�������?,k���F��C��_�5 K*���4�ˌ�RG�3.b�H2�S& X������o��
G���`a�*����0@��x˿���!�����������-�2���?�M�7S,Ny���#��춏�R��r<O���ߕ䬚���p���n�g�PR�j?"�d��v�z����HcŽ�QAR�[<�}x[�|��: Q��ܻ��x[9�Y
p%e��(�%�l�8.�G�9�0b���MQ�N�r�o�>{��D�JmLczY1��'�> ��+�7:�>��4�v˰�B���x��N7X:�I(�q���`�K�\0֏�I'�绺bخ�#���?���%n+vǏ4a�.��fS��U���?�mT�iE�$a�8�47�������N����F��;����ᴯL����Y2���߸#`��
�w_p�>>�?+���x1!��������u�l�n�3!�"46#�x*jWFW�~����X�Ku��k�1��qͿ�k��LhQ��nN6ޡ����z����a��k����P�Yo�$�I�ysZ8>8	;��o���e�ܤ�ږs�)�s�W)M�`3n��^!��	�Zi��sc���3�av}�r�k*��+H�wk[,�b[?x�6��p6�*��
E/4�����:D#�A�K������q��[-��P�n�����"P��G�����,��(Dͫ��Ȟ�i_��R�W�i֦�2���E�XD}Ʋ~��D�F6�\h���2�n<f�ޞ�9MSɪ[idj�yE�+1�N����!I��>�x��G�e��*�;���k����gQii�(�j4~�|��Ag_Q�?[.fs���a��ĳ&28�U�f�ኛOK�5?��Io�vv��R�E��o^�h)��/��d�{�k冚>�U�����63@#�1�}>J�4�/?�WS���ͮ]+�/��\���x{t�S�s�$�yB��s��"ݯau�s@��l�W6NN��n��m�⾛_�«r1H*QLp0��ba��;�z�?-�o���ƯO�f���-���?���ډ�5�hoy�9%����V{w�#"O۫�q��A*2($�c�1I�rWv�w�x�������{3V$��k�H_���_�T��?z��=ݘ�I�@2
��;�����>���&�LSSfo��i���Jo1j�#����P��S�Y�w*�����|x�'�h�+�/�+�R��~�[f_�;-��-Ҏ���������ƕ2I]��~~#m�i��v�nk%�د�m�����e����g ���fY��d�Ļپ>2����r��5K�����[.������~�%	#
)zZ�fZ{5�b�T^��V֖b��pH ���oȼ��D�X�oF�T��jxЉ!p2�^��k9ra3E���^�4Y�~2��`��{p���إ%mm�e���?��	�f������#h��f��g�~d5�Ȗ�LϏ�r՗L�����)2�N�)��񜭞�E`aD����m~�c�;�z�?�v��jf�ǝԩP�G��cW}��JƬs���dt��7*�7��`���w�J\���x�)���~N��ӓ�����M箉������˩E���GZ�>FFT �6Z�ݮ��_y�GGz�2I��f���!��� %w�b�Q�P��7pU����d��&Q�&n���`2��O@f��p�e����DC��D�5���OD�g�1�����+��SV�GG��.����8�A,��	�ۋ��[��zӫ#�:NF�RQGGGe8����:n������}�ߜ��?����e�����H���mhÜ@�[�N�_�n%�ޝ?X��NtS��D*�ȸ��o T\����� �o�Ji;�R'VUS3u��l��Wb?
b�OJ3��&~���z�L%���/f'-�0�_F��!_^7n��!�t����R.?�/�$y�fȹ=�~]�.M��U�G�SD!�أ��M;v%?��*��J �Q�QS� ��5\d��H$��]�}�:�%�?�y��-�<@x��s���c�؁��B��3j͏m���\���Z	ږʟ���l⵬k��H|�L�%�c��x�5A��}h�������ʉ:]�J��s
z�p�D~<ͺ��e��M[��:��BEaC_��Q@���P)�&���w��y���%��1��DKS��,E(��h�&���_X�{:�-y�!A����tkcD��b*��"plL~��c��Z�7�.+0���.���Bb<�Wyu��7�A�qAI?���_?���|�c$H�h�x�]��~���l�xX�Q�����B��~��Y�,� V��6�#͏^Sc��%���/�ZC���J˅��j���=��TE�(ޑ"-��z*H��,b�����y���Mz�����e�b6.H�ңdcL�^HKj²F�L�5��ƃ�]/��[M���o�O⪿7�K��9���f�X|������t)Ywi�^"}S��,��"d�uq���t��a!�Ґ�b�\i��&�M�?i��B�ܼ�m	z�Y��ۼe����!�:4�ϴ���^�d+wji�Hf����.���x:�.�tE|���-9����l^������{�v����� �����?5H~~z�^�+���?��k/��`��y��vC<�s������C�6KWVQi�1������G���J�&��h�L:ބK����-�-��I�zL�w2=��D7�/��� mtnW3��P�P3�	���7hhhvw����:ff� Uv�LP��"�25bb�q*jQˀ��V�jОF�k=���4w��~a�~���;$��+�W�aN�\�)��Ĝ|~�&�m��7Vz=���I���K;v�W�o��
7qi��Ŀ�{�͙qE��>/D���af�j�l��Z.��_����T^Pm��37`�P{C��}�������FI%T�L�m�����l�䵶v���Ա��Bc�hĎ�~`����*��@L����6�QQ��!��3H��\���5��S�P�԰l�spx��v�� ��Ll�X"���p�Im�&��������8e�	7t����v�ł�e�:�"��@������́� ���P�.��!�*�q�`yc/�Γߩ� z��A���K�B��t]��7/O���n��O��2�)�%uL��V���.R:���F"ΐ̿���|'KqS9C_�H��6Oϑz����C�J�㢉���:�o�[=������\N����a���n��k�%ԊB�r��ףݐ���o�f�v`]�$�u��Y��$�F���I� �#��H���XG��<�)5��y�@�v?�mҹ��D
�N����3���B�*�����dϧ�-�-�1ҧ3�z��9~VV��mQTU5.��q�R3Z�ˢ��UK�Q9qqT���Γ�y��V�>�k�-3k�[��1�;��n��f�g=/p��[�^m��TM
��,YO�����0k-�uE{�Q'+���@F1���ɬ]�'s�����Q(�F��`�^},���f,�V�Y�z���&ƳŌRm3�Ums��Q��,;�bn����m+N
X�f8O���8ӌ�ͳ�!Ɗ�/�:�W�ג�w��<��P�jߖ+\ﵟX��U�l%�J��n �������7���G�[��~T�\(�&�N>�u��\��S��^�Iq�£4�_#6Ȉk�W� �=ڌ��ǒ��ya�h��>��B9"��J�PL��<�	 ��2[o���^M���GCn�ċ_5
	�ksRg~U-K��_\�W	�dȶX $�y\�&h����N���Y ��n�v;o�%ux\[G ��I�瓤��N,Z�m�� A��|{_��jC��ZG�^T
���D��e.�`q%��
���h'Tk�_�"?�0�rդ�=Bd��9�m�1|}�'9jU*d����8@.��qW����?�B�kGN���u1���Px�?ؔ��0YI�{)koan^`���o�e�3ۡwW��-�~��߀� ��AG&����V`��I�.8If@��I��<���s(�◣��X��]��a�����7���P�w?~�XK�j��t�����Ω�n��93W��6ǾQ�.�۵W	���.��-V�K�-9�00����"��s��x�C���]2>�[��ͼ��)I����Q#��-A�^]������
��J�Y��ۼ�Y1�٠x_��X�,BrUDU���!�p���k���i%�H$,��=��,n'	1+�������PQCp��I]]���W3@� a��>���0n�D��ʉ,1���-��qCj�wu�^X��5�^����,��~C.��7��ú�o�A`9�g����1�}�F�%���ˏ�tZv{�$�TUy��g��?Е��7�	��E���gy�v��'�տ7��_q�AI�G11��>�͙c5�4�5������)�u��l,�"�D������b�{	�]v����Y�;�y&��{d����^�	��{��j6��*��.'9kxɊ��
8Zơ��h�`S{�m{�;
�E;��Xx�4�F���>G�Ӣh��{?p������n�^�G׾�W̯�/���p�ll��Y��'�:� ���gT���,��e+iW����f�w43��|b8�^'��N|��9!X(����Ծ[��Ӎ��܏T�yC��Z}�`���R�Gw��x�q&'YD*9�d�̥����opc�{�����ٝA��ʭs�.z��Y�r�<U�\�럇�xxF��g��n���k���o'�L�b���`��y�Z#�P���E;R��Z����aP�c�W�B��Ph}�m��>�ڝ{�!��Ɔ����6������	�޽�򪫕onli|w�⏫~g�1�3,�#FW�L�{r��tnuAr�lXʏ�M���u#���3F��~f����f��`���7��K���;�ߚ]���C����O+�z������� �8u�xc���Uc��R	�l���hW]���l��;��j_�I;<��a���I�`ʠ-�y����pں�%�q��ļ}��{�g�:;����9熪�Կ|1�A�&8_k�@�Bh\��P�V�:��{Mۯt2�iU��v�w���,��(��\Ri+��~v	�SG4�J��-`R��	�����]ն旝r��;Ocj�2W�ObG�z�Z�lh��.ɯ�P@2���׿学ԧ$M�����ۺ#s����C�F��I���NZ��6(h���6x���s�i]X��~�2Z�`U�+�,0y��5��m�l�|<�6���"N)U��H�?4����șc��u�������R�l���]�ź��ރ��б|���7��:vk��m��0�T�Q��y���&C���� (:���-K�j%�PW(�v���ۣ�jܝ�o�;�.�>	��L(�4z�x�[#�J&4�G�����ɜ��}���Pu���\��M�.�����e\K��
�Kxy��8�Ɉ]�!��q��RB�#��x�]�������s]A��'m@��`�� ����p���̿�ڭ}������(�(gk^PSg��7]~������5^e��h�(�.���JY�ݹY�zo��	q���y�s��-D� 2�R4�!K܄jz�|B�W����W>222vP"��r1ֽ�}u8��Y��Aj�������% 7�51���*毴�׶�U*�+�-_#B�eׯ#l4V4�4�_Q�s?ּ����j��g��s-����Y��=�p n�3� ��Y�I�Vz�%�Z�������^���|#A<ߩ)l�>�s��g)j�P�ܰ�����&��4?��?�r�/#S��>[�����
���5I�Z���t��������;�<r��w��#@yꎳ��w�I�K�}�T��k��>w�m7��'}�:� ���hXhYk1�כ-st�V�ش�K�XJ��ҭH��S�u��E�ZL-ϐ�=�5E�q�$�#��Kc�["|�Y�p��F+u���)���)�q]��w�x�̧J,��,>s[q�*�z�m����yI�j���r���s4詄��p�� 6*iߋ��V\R.�����0aj�	䥠�#S�Ma�(Ĥ�'���0u�h�i�i����u`1�5�ԍ9�s�.���v�C�t��v���g��t}Dd]?�T�w��]��{��@u����ZJ��}ȶ�<�Y/S��0���@[�!2�˧�7�<=��"���1�P,�%f�rHL�.���'囗�>���q��u�O$RPV��c�T����t/eQ��"�Ъ�Ҕ��ɂ�_	ǩz��1+w��,(R��L�G��,�Q��7�2���)�Mv��� ��!�'����w��O�Џ#�b�(t�r_<~��s���3Z�j���z�M�8�ֲ����.?
>�nSԫ�ok�ds	I�{���s�8���WM}���q�L�r��*�G�ƀ�"N�w����WN�M�F�JP5V��V�̃s�v�^^$�aʒ�˓�p��@�0�QL/�,�������ː�h"�[Zm��hN�ۭ7
w�{���i���թ��	�O�!�_2Վ�y����B^Z����[LٯI���W�(�]?J�ɕ�^g�v�EG�v��i>sC��[�R�Wr0Vs�ʞQD�*a�0�ı.f�a�UB����\�A(B�m�вݠ��b��|h��q��s	]QJ��HΩ�e�t���t!<�����f���`CO!��,9���oH��>�-;�[��
�eEٚ��3��5�ب��Tux��k����?`"�ݨe�.����Mb1�L#j"B��7�+?�����q2���My�w� 0����/<�4;u��>;�d�a߬x���Q>���걞fY���������J�)#ݣ�A�x�'��0�a�t�V���G����'n�����w�x�q
�ە��d#O������ߝ�m��<�"�8/�_�@��u�x��],D�����coF�=�����Le�"+^�?oD���m}C�z�W�1�K���!�@Ϻ+6l+����P(���I`?���K�ͬ��u���,q����1o��]��' ����@��3��%�U~!��B����\{`0
BW8��[o8���QmQww����a|�;PfZ�W��8�@A1������h $<���DC��<+2}���kh�N�<5����4
��d�P���H�T�]�Zq����C k�J�� ����f9��z���w�JU�t��-�~ �ӕ		�z�5(&�K�[����BP޴C�#9�L2�z�xx��BQ�{�Hg�X��� ޢ��8O��7V�d/����:���Q`g�`^�����=��A#�T��0���mՃ�!]�'b'}���U]�fީIO�s���Q�KRc����s2�U�Aʯ��}�'"��<���"#���z_o��WEb��C3�pť��M���J,)��P��XK;��Sl3f�6�J�PH+p�<�cp����{�Y�7$�u4@=ojյ��h�҂�N9!�k����ݡqzӕ�T�]�-��3��튲�T�3-j�����a�,�K�������t������KG6���X�� k���p�b6ƀ�sR�ˬ���z�V]��K��6#��ф���x�M�Y�����
�3m������Y��=�TH]���y�څ�d�2=�4�ғ��6�fD�~hWⓉ+�%�(k'�4^m�%M��D6�\a���0��	d�N�J��k͑$g�X5
�ݞ=���-�T>t��ǩ�����4��_-@�ɇ��
�Ƌ<��6� �n����G��G�B�PP���W�ܞw[�S<����q<+<5FX�H�����E|w���9��ef��!>������-Zޗǋ��n���GZ�5_�� �Ʀy��:�!�����C>�X^	�;Zx�%u	pB@��D�yi6�X.ő� 1�s�Pr~������0�?�v��-�p�c?��=����^4"#�`�0�<ã+�:����k��_���])�qb�5�O�䕆��0����hj�{iT
�{�n�1�o�;��G~�`���C���p�~����P-v|��jQ�҃�DM���@�=�1F�~�q����fw�Zw�i�[z��5)]�7��y��3N��)��E���#ꭣ����q@:�� "�ҍ�tJ��tץ�A�����N�KHww�����~�\ֺ뜽��<�̳g>��!zz8.RZFw
ؚ���=l�S�=~�ؤ���ViU�o�(��[����Z�g���65���ھ�?c����֨i�$;���K�����WDxڷ�]`�<W!i��[��o�o��9S�q;�P�0)�Wz�#��j�#���YA��$a��0b���M�{E"6���&K��Y��t/��1W�tɗ�FbU%�����)�C�,u`���
=>������o�)F��cKz�ڰ�ȶ��d�	�g \��� _�]�n��X:��J�����_�)+tc����S�ɪ����Ah�x���dg���]`��R�1�� �B�G�F�������T��0�w/U��g�|p���,
��b������`� 益��\��7S5TK��QȂ$�>����D�Z�ϻ�Q�a	>�ɳ���E�i�}��'����%fWa��,{����`w�(kDv���	�K7�Ph���޽���A�^�%��,3���6UA��Q����^p��ڞ����L�iJ�j���Ep�@~�A�%q�~�Ulls�7��u��t�T�(^���@x�Ӏ�3�:�nz��`�o�@���٩�����P�(�NM��3�\���L UpvfE�A�i�5����sVK�@��e����0��;�I���g���=We9�U ���8S�Y	��X�/5�'�V_q�p�v�L�|Z5:��s�¾;0��8x��~K�����y���Y�����]���V������?u�\����@���������6Q��w>R��\�x��\O��J�iڻz��k[���0����E��?E����W7�T�2K�F��cN"Y�C�%�\2�Y/�^����Q��UH��1s��i�?�~-z��E�{���w��*`�l�W�_����.7Kl��B��J=Ijj����|���Ǝ�ǖ�������ɘJ��@�U���N�p���d�ˉu
z-F)d�v�{��c���F?U"5�c�wZ��1~^nL��#B����(�V�T��:bOp�fdg�-�[� �0>Y��ip�l�������
���$���}P~M���*��d>��C� ��K9Vi$��\kS��6c��q�A{���&��ǜ��<�e6�މ�ы.�ĥwgV�t銲��GaFҭ��=$�i-	�+�+1��p��R�>ެ�oɟ:�8מ���F����l~t��?�}7I�����kv��p����x�4��a�|�c���{FOI��h�����%,��S�gKGr|�x�m�me���W����h��?=+��j�t�&�{f�}��B���0Qz���'*�EuI8i�f
C����0���%���j���L�>lĈ+��@�xS�'�
&|;���5Cy�9�+:>.�2z���w�=Na	�K��;PDv�9��_�E��z'������E�O!����.y)�`��B�~� R����E��ܠ���D�\�3�e��}a
l}�$��C��f �]�R����=�����ԯF0cv3R	�_&7u�]���Ven��Wp�찒�<�W��:stKR՜���C}Z��$��Wz����v?��E���_��?u�}�|9Ϛ�!��O�׶��Mnz=E�;u6���ֱ�;컨ٳB )3�S1���|�Z��ˣc8K�2i�e�k�o�&�'����ir��oS�}�lF���`�ɀ�a�2w�`�}�VR������jة�w�W�m.��a�>�o�R �;;>!�d��+Y�_$""�����F��_�P�x���P�L�-���kQQQ�k����c6²b���jf� �V�/��ퟛ}8z�j;OF��b�7�cX����������%�1���;���ВXO�A�1�mZ�������׼�1b�6�}�M�|��9��6�I��0`�>��W�BYNm�p���HE��l����i댒�Q�O��*"i�Ob��|��k�����������Pii��ь�
l��e|f��	�J�Ji
7"���|��(~(����UC����܈��������E�����e`��
��^Pцr��	�{�q| mp���m)����a>�U�t�~ӱ)�
|7VPLd���K�E�������CV�(.$w���>�U�@s��H)e���$�a*;$���N�	�%��^
�rh)Ƒ�g(�����@�����z��i?��ؘqѡ���1����֙3F_+�n�lti���]�=DCMm��I< v0}�R)�\{|���?5�4�C�qؒ.���'S<��ܘJ�N�]���cE���2F�]�s<���^W��H
FTL�\k�	���,�|��+��$� K���mi1B�ii~>�Pr�뺂�$pf��G6���A�iȬ�FJ
�T+��`�n��vzMU&")���/�\���L��#�Jd���o���<�ҷ;�!y�<D"ya�'��T�qC�&����C�bF3�����&+����S�G���~�!�/�h�H�,�$����Z��|�kz_����iX;��b��&�ƪ'E�=��x�4��eV	U.��mQ��̗�u3��K����=9m��ߔ1�Z�p
�4(��f�Y[s��`�X�h��-/\�Ea�jq�� ���4�]`�S�k�M�?f�Y#Ѵ���i<g=��%1z��|,>Vk��X�P�>�@��hAj� ���b�G�U�������ƒ�9��ׯW��.��γ�w�������Ҫ��hR���P�\BBB�����o��&&Vu����`X H���z[�]���^���}5j^��8����|��U����M�ý���8&���5�Cw�Y�8#F?7I�7.�1DXIQښn��Gy�4�]���~ge�S둌����(��"����U?��b�����9�4��&j!��nu�[V}4	�$J���_H�H́���es��8�l��<�17	TI���[[[�}PN�䢟A,�MU �K��$>��D�׳���)@��~��d��R��VY��*S��͠��2ER��Ҽ����9��\�D�u��n�̎�?A5�k+%+�/G_���K���a�/�L�c���⠳R���GU�;�ýB9I� HUW�����<'� @F�����*�������Px¥�ځ:�՗wW�<3�A'k�o3���c�̜���ol.pjFC�oC?GT�.��L��z���^�=86\�a�W�{uE&"n�X#�8��9�H߄q�5�=F��ڳ�~���]�a]�E���z����)$	��X���7P�����g6Rw(�x�\,�av���xR]�� �o��
D� ����+@�*�H�3�_��kp�˜x]�G��RӬQ��s�p�hr�{UC����AU��~��d�wKk�����m�K2��s;�o�>��|�#��6|�nUg�iv���@�'C�<���Gg���d��j�n���]M*��iϼ�apĮ��f��}�t�
Q�ZA%��b#������}��0��׹�kc��>�V]x����*�������ժ�m�ݖ^S[�K����丫� ڲ!k+8=|��*�Ę�:�9��3����H1e��$C��8�8�q��f����?��*F��پ/������ջ~��]C�����c��S}���2\Ҡ"�bSF3�5���DE���>�-��	;n4�ݭa�eV��^�n��5�V%D�9��� r�|�M��Zfw�Y�N��']�:)�+���y�Ar1���;I���E���9+ƛ��(�z�
����!a��e����n���=u���cg���jwd�ò�_�n7YЃms�{PG��G�qs��Gr�ˎW�<�ʏ�����£*�_r��Լ�ڻ���2 ��Q��Cp���!�&$H�g*���
9jW!���Լ�b��+Y�
zuU.F Lk:�<4���&����e�6��g�	�}^O�j��`*)Cc��.YQo�����2����}�OoKqh)�����۸n(�;�ջ@�~v�\gE6����Z�\��us� �����q|D[���?��Y��o��r��<ρ:��fqG����e,� �	LH�q�g��-B$����k�o�<J4:ƨ̡�nʴ5�b�!�m��ݝ,�}���e+ßBY�1�\T>)	�n�5bj�;!r�/-���t��:�^�|�����e
,g)k�{2ތ !q%�L`ECA�	y�#-�Ul��®M��̈E�V�x��
�{��u���\��jW�4ݤ4��l,>a	b�DP�j�?��v`��i�����a�^L%�;	b���Q�ӚX:��Z� �D��/�Ò�Ҷ��99��U�L���D�eK��g��܆�!��!Pk1�mX<���p7�k%jj\\0Ĳ��
�������������Y��*)Q�;�\�� ��旰�*�9�q� v}̢o��y�6l�Xv����jF������]g,��U~��V��bcq��9�iz��]�]�Tn��N�wȼ�
M�R�i�9V�s�dΦ�\/ߗ�u6��허���+��Vt� �,��%��вM�]⎻���G�[�ʹe�Iܖ`r�+�A�
?��'��[��y�<�]�B�[�ފmD�IX�-o�-����~�4���2fFO�3NOWf�5�lU/�N-*����?/�Ő��A,$H�Qp7��10���I�c�}�GQ=�Pʬ����][W�z��!��PM.������ʙXx������9ˌ���Ē�V�!妖h�nY;}��>:�â�;����d����fd���QӤgͳO��Y&GlY�-'�C��$���7�8\6�N��<WB���݀)���&&�`�l�.�D��Qf�Ƣ��OWB�d�o0*��3k�K��A:��`8Q��n��^ ǭ�� x���O%a+uZ[�*�z1.#�]{/"@�G�hĀog��n���G�OJ�������R�>F����A:_C���<o�"y��5D��5N��7M�0����c �po+��8d�����,e��X��A�yϩn�@"U��F�� ������:_���z�������<�De')����f�=�>֬�e��W�#��#i��.��Q�ߤ�Q�tϚ�l�O���T*̏L��\S�ԉ�~\�Fh;-	Iօ�c�qp��G<Ǩ����"�g��52�蝖nF��w.>�li��U�
��������9��wn�	zm\?��H������ߜ�`����O�m���|^3-��L��Fh����{��'�(6D�r��� T���s��4'��<{v��q��)�6_�e��<<_�pE�Z��7xm�z�[�m/Zq��\i�/�Z���:��ۚ���g߽�$f����F�4�1��Wթ�'��w�?��0���r�/�ǡ�b
/���ql����=�%X�ݐ����j ��|Ps�Je�#��;�Ɛ9�`2���R[�)�tm;Qo����~]�4�K�K��eA�E��F�-_���3�{ktؓ�����/W<���	g������an�De� a�n�fJ�v:����3�,�	�
��;�e�����~\p��K�a1�cyL1$& 7E��ވ��b�@/"��&Wg�D*�����t�k�}{E|]��*ŷ,r�l�\W�H��Yq��s����q#N<<<�s�~�7g[`9��tcp���B�b���氤�9ܖ/��	�TH���a+W��*��I,�a�Y���텣�KY�֣~��"���&�9��(h��#W�R�+�.��Q^c�b�H1�8��tAf2!%L���9���R���"�Y�;��+2�r�4Y<0�Wʜ�߷xP	�h����T8�����D��U���>�^��<�
>�� FTe9���*\����7	��%~���`�A��jwߨ皵gQ�tP����m��fq�,�Z��xA5X��UX���[���+�����c��>�90R�,��,�D<��u9&���ѣ!ٜ�H{Y���A�����>yzt����p��^� �c�J��� W���+�?���Y�1}���s��Ou*�����CG�y��y(\����[q����
���⦛�,��)�Ex�����I�F����x�q+Nu*L�jX	��4.��ٱ�Q��U`k_~��{��u �J�,,]��p ������ϯ|q����>�y)�k�����m�s�"ˤ}M�"�,&�;�
��,%($��y��g��,�?[NMz��3OM�8kE*�a�NI�Q'I��8�P���אE��
�&�tm��(L�
&Bg쯹�V���		6z�#��T���ޯ�")�_p����	%Ѩ��u��N�����|8��h�ݛ+��*aN�j�/wB���5Н"�r��ؤA*�O$��)�`����(` ���
*@6���}ç��y3ב�}��%is2���Y���s�����5m��9��F ���᲻�u�xj���o�EHct0���!�
�U�ڌ�
e�NL�P�r���D��=J,Q1ҳ�2P3���XA� �/�03��֗�E��!$e�9��[?w�p�0w�
 �z(Id3�� �uX_������w���3�M�nG*�d
{�Lu%ŷ�%ă�|��!��:-&�R6�/������5����LÍDF$�߬�d��k��N8���\a2��HW�m��H1��㕮_Q��j|{)��KPC�f��k6�Z'k�`�7Z�Æ-��P,�݂���#�t��$!��G˔ �_�[qo<���I�_�΀�h����;fl��Qi�&F`�PW_�ih֘�+��]����Aٽ��2ϒ#�$�F�P4�w�g\�R7�z�K[�)�8����Fv�"6Y�o&W�s-Q�l$�
��-����>o�GT��ſ���趤��L����u�N�%�S�u�~��]���N��L �V?[��:��R��s�$R����'�2�y���)�d2Э��#�'����`�N����E�*x� J����6�aར�U�s$���|8a��G
o�G3��nFS+4P�"�(Y.���Ė�C|�u��vGW*�rGS�C�ً���F�v5NY�=����t�=��
,f�R��� ���Nxv27`+�y��"��o�P�
���HǤz&�f!]'S��>ajv�$�4/��#�	,�y��[���hVP�7
>�iV�q<]�R'0e��K�$��f���w��_��FV��x��r�(Lj%����!E�/?=,�9PhY�S����;0P��������1s�=�Lv�T2�o^��h�I>p��ٲ���7��-��
Lm�h��S,�9��=��s�Iɖv�� ���jͪ��M�:s���*�B6�'y��W��o�K���p�
���$�`\i�ؗ�����A���t�>���$�v�m���������*�y?�A0��	�do	�J�>�|[���� ����}!�{���&��'�z;�$*��~֋-��hn���&��y�����>8ѻMC@� n����� ��ӁLL冞7�y���@J��3�T�ߔy��O�S��
Y���Ʈ05�J�ɀ�n�:e��qH�����:w�zp��G��w~�҄����|Gf��] {�<�U�7�45	,Fӣ��#N���2���������"g�R�ru��n��E6��m 5Q��%;h�9n,6H��fƩ�j�ۑ��v�Uճ�#�v�+�Hݓ`$�	�Ǚ7P।���vw\�Xr�-�)�=59���Ȼ9�Id�	����Z�˺�����^ as �nMIkkSrVx�x��(�y}QFo�j<ﶽA&���Ju�$S�����7����۰��A��2�/��pw_S�@=Mk^���5���2eT�}��@����:,��,�zc}��	�f�f�T/ܿ^a���r4I��|s��T��?]8~��el��S���p\hp���;�r��߰*�r6F��,e��7-�v�ڤ~�ԃ�����2�WݴZ���\_�l�/�p��-m�a��)�5�7��ؼ����F��w��j�d�U=�*��Ab���;��Z�	b�ύxÜ�~<B"�sRs_
�T�����}пhjj��3�?W^ic1��wu�^��&��S�����O���ah��ە�:��U;h�x����nFnU�e������߾�$�|��4	#���!��M.�����i���Z%�
��>O\�D޸#K�&3��t�%P���k�=M�Q�����Zѱ_܄�Bg�CC}��|��|�T ���,�F�������X��)Yn��f���`j��a���v�_غ�� lJ�� �WG_�,���� ���Y��3�TDn�t	6|ߙ�l�mْeҶ��x��G���WU/���<Q���������2@F�(��y���r�ߢ�Ҏ˳�o(4�g��!����¢%]�Ȱ�1^��1��⧟�p��)m@]�����ѵNlQ�����\=X� �8ؒ ���<R=T;��"�ˬĘHXM����5R�3��¡��@Y�i�NM޳�SZ����D��j��S��I���(��1<��C��[��v�+��"tL���
�u���F�(�m̻_z�Qc�a�^m�L.ΰԶN�~u/��,^bĂ*�4Ψ��oI�RG,�����{���Hr�dhr��u'$��p)+4�P�%��jz��9�&�S�!���XA�Ʃ��D�|��}E(#�{*e�}B�^�e)wE��ƺ9DS����)-:�/��6Q(+&��i�'"ۍ	/��
�F6
Q ̟M�a���C'T�F,�q�Igp����~�S�[��M�@x��{~�Ł�mrs��J@�g#h�CW8�O{��j��&��r��*�����ޢCó�/߀Y�{ȼd�J�qc�Oc���w�4��u*J�����n�a��!�A~�z�Qt}"Yf��;Q�PD���j��c�	��p�:z�vW��)��J�|a�=r����,���tm�E��?X�ykO��*u0ʡ�F^�<2�}bAw`�#�E�Y;5����сQ���R��g�9�}{�U4`��$��������Kv�|�:�s�$s�Χ�ۤ��Y�֣��:�ڰ+�_��gX�Q� ��T�J���I}D��᯶�9���H\�ѵƄ[�N�^+@�V3�&���ƙ���*ճܫT�f8� V�i���Ov�Z�z�t9�B�`����.LW�>'�
Ŧ|N�M��W�Ķ��>�4~ɝ�=@>��Fi'*$���c���:�w�p�%�7&j��8�(Oh���/�:18�!z�:��a<��0>�;�a�#!�WU��P�?2������r�i]���n��`��K���"������>�<5q���#x��L��f�y��A(�=���"�������P0�	��\\\�}�ƚ�p7��$�)2�r�[Ը���~a;M���B�� 9����S-��Wu�ce�s;�O��o0���kM���/l��Z��G�_Ù�K0����X̥�i��[H0��Cg�H�AN�q۷U�n\)0@ ΄�7řs��k��өw�6�9�c ���lpն�`�_�W�b�G��	��;����
�*ݑ�����Y��?'�a��Q��-��J����	?vLC+�-�_mb;a����JD|������S�a����c����ή��M{���������oiM~�H�%���"Q�Q�Y�(s��.�G�G>�)��ڶ9"�4;�>FCX�i]���2[��A�5�@�~����v�2z�2��Zc \�	+)�E�����C��of��A�b��f��)c%@��S�1+הoy̶�RrYe�������V��5����{PO&���Ʃ�E�C x�W�G-T핧��f��c�� 6z�qb��9IG��yR[�Gx&�@���<ׯ쬬�.��/)�����3�2C���������, �����	)�������\�Ww��>��Ԋ$�u��Fc���P��������u�V.�e7.��.�-����u-c�42��H��k���X�:�;� @g$R\����L�����ӭ��C����W�a��N�j^�^!Qv�V8�G���L��e�����m�x9��9��Ф�0뇆�d�P�ƈ�F��8��!V)__apѯ��)����mo�W"߸#4�(�>���]�f�����ݚZ����Y>E�
/��xӇo�� ��y���2��\�^����_�8��	���C���qK�%j�*0��P�U^f�`��n��5z��4�_}�snఞd�����乆ŢW�)�q�c���AN���33`C�X��/=.]t���.����y�����f?��LB��x�c#ݧ�z�#��������R?;�N4���Y��'��EO���%�+\wt~8���JD��~ʢRw�4F#9U��C�Vֿ=�����s����5،߆Vz0P���R1T�n1!v�6Xʈ����}فkL[�bCE �ρZ��Fvph��`����1���9(`UJ��"��W
8b�:o}���%����W6��?�H�`f�b)	&t�ϟ����P�j�&,�Y	|���+q��S*zp�kʟ��6G�Z	fA��y���+�4F	f��ψϚ+�j��|���Ls��IV,Sk��e�͎S�ڠ��s+ͣ�v��ب������Z���2�h�-- 惫dV���#�fdv�b��X��y��i�VW�J�ѯ^��c�N�p�c�2���ee4�լz(^�va�D��ED�i��Ӵt�/B�:]{V���y�eo��z8T�-�L��=G��B�@>��s3�>�љ���-�[�7�(^zv��G�x��h��,:�pg�Ý��/7�Fo�;l<�@��B��E��tw� ��Q`�7�~��l�4�4 8y:�i����2C[��V.Wٚˋǣ���o�!�� C���=6�u��#��ы������֒�)�J�]��ޘf\��"F�Q.�v�.w�2w�:�9�:[yMg5O��k�- ������L�.��B'�Ee�h �2ddc�	F�g��������z1�Ü�]��5N:����`c$��"	Wp2�k�}&�I�.&칺���6U���T�w�"�w�`y�AI:�t�[y��� H��ҽ��m�=���e�Ne�v̿����j��)�,�B6�(��&i�5���$�k̦g}�)�>�Z�%��������.��!�'�Z۹�$#?��s��do��'0p�%���;��c">EfJHs��̏�>LYJ�~�d�h�ńjIA�s���� ʬ��\�*l��3�_�K�mc�<ۤ��D��o?g�cr)m�[�!XM��\2�	d�DH�jR?'�
'i4�=`q�Ͷ�
�s�}�4��`D|��x�����}���'z�H�(���C /HĽz�q��g�¬w�~ܧh�N�k ���]��
O1�`�Ʀ����IզQ�L�c�=��X��'�{��v8�O@8��S�5�\j��Lį����!_�������'+�C[�Ow��a�'yu���Rqu���u�4D�Y� � �c
� ������1c�L��6��u���sjk	떼�K�/߃�j�Zn����|eq^�;i08bƀm��#TUT�\�����*�O�\�'I�	ͺ����c��1��r!0,���!�N���� � mD�����|�����M�g������E�������`S��v�Ě�x����E�8X�)8��łEٹU.����� c(w�RۇXYY�M�譕* �JIS����XB��k4�T'd8h��`���o~�?̸��CJ��W�_Z(E�E	���Xc���e޺yI���r�B*�?G�J���^�t�*יY�R��Z�F�V=���r�d/j-p�]��{\S���1�1�+�xNo�Mw*�"#��.H��C\\��>4T%MR��YF���R�s�Yp�:��VU�Ȓp[dVT�i�t0�56C��m�
������������y�ݻ�Vm��FmI�.ڷr~<3��d��ъ�X���B^|w/����#~��]6�U���>��qܗ��KZx2��@����c�jw���޵���{�YX̝��%b��x�i�p1?�-��^��3�Q_*��)������CJ��\.���`�w�@
������Z/�An"z���qhA�|�7Yk<�Y���q�k�|�S�ԔyUl�J��l ��M�ܲ~�ᯡ�~ĕ�����_ ��
��p @������x�Wǉ`�L ��y����(cɣ�&�+kmބݰE�8D�@ԀLƾ�o<H���pꇅ�b����$�M4����|�ڛ��3F_�I�YY�{�%�66��Η���s���opr�~�]���1�<���#�� ;"Xx������H�R�:�����F$��c�/���..z_�D���`펃(7\���VWCEL*3B88$��!~�_&� ��_�c�� ���!܄�KRYY]�g?X�����)u�p�/sZ���a�������9_E$��PL$di�K�`��é�R��U�\Cq� ���^��śƯ�5��{�F$|u�5Ҍ�NL����ӝ�:愎�%�I�DYݔ_��p�<�lŌY�������\�u;�`
ͥ��(۷��&�|�)��]f�{c9�{oBB�Z���f�:��_�٤~}�����d�F��;[a�t��
���P���r� ��	�-�9�?����=c�W:��(L͗n���մ�3�\���tG���ś`3�E,~VL �'�;gg���d<żԵv�JT4���+��u����R�>���!��#_���;;��&0���5a�����\p$���̀����<`�9�^�D��s��z�:A=��,�e�������%64�V�)S��|/�Q��x�b��`���9��5�Yi'\m�-:���U������1��］n�	l�	Zb��&�du��������dfE5��+x�Ӆ[�H�g��������(��La�u�:��=�噧����4ع�׻�����C(
6�O#Y�����bu����HD1���>=�Y���`-�������!~S����:�S�%�@��&��2E"6��Y1���5�5�ru����v$z�u7�[�rMCAa�-��2��R[Gmt튞+�z��4q��	�E$q�HM�L�O���Z���#�����T�T�~��]��;����`"x$��z��1�nُp@��ݘ��%��444���9����F��� �ɮ!����n��8���0�Uɰ�]��������h��}������U!����K6��~k�9����S�2B��e��P��£�����:U<��N������Jy�����|��-"��F*�|��"YΊ�t!���t�������*M>X�\�i�g��"�����/ɴFs����0�9��n�'+a���L	��v�t������j���񜷝���s����{6v6��oz��L0wW�^u[����S>��c��h��Y�s�����~P��Yu����9%���6�Y�l�<�g�膳.F)��i-j�Z1��eyL� ���@M*Y� �~:S丠�Q%����]
�J�R�Cӧ�0�N�l����ޡW�����E�CBB��'��g#BG�Tu_���W)��ފ���%i��
/V�^�ޅiW8οw�&'}h�"ߖ��Н�2��?n��GC�y��Jl��*�`W���v��#��ga� �C=��ټ�/H]��P����|�����^���B�W�g/�D�G}Ԩ�H^͊��L`Xg˹@��T����z)� r00��a��J|��%i�2�lx�j��E`�^{l1��}����ډ1�ܜ����YS>]�������d�z�Cp̥ d�RD;	6�a`eE��>��xF4��]=�$Ur �z���v���#��H �Y	j����^�?%��)����;����?L�K�Z�5��Ϯ��d��	����G��� i���$����WR�	:�3cp%b!}K簅��!2�g�Æ�/y�_�P��8R!?'O���F�k�����}�h�&n�������*Ҡ"���`��PJ�|y�E������ŝ="BB�'�]|%�# ���3����o���-��D�\���a��/�)�[)�كM0>hu�O_*V�ǻ�Jt�����_m!�f�Q�u���:J��NR�����\�1K��	Y���Zz�A��:��9޿`�Ͷ;� V�U5�Q�U���¤!��ώL&)�]�6��=}�X'��=m��qpWtr��4Nk=+�0�N�C+�iŬ3��AX�3��ҹ��og*DQ�h�;�=�������C C�A-�`4��*>'ܿ�p#�;�$	�M����+b��lJP#�N�������sC[�\�xv5�([K^f��%����9�Yx�F��븂_���܇Wh^T,������ld��`�3^�,%,��sٰa�����UI��pX������S���t,����H��B�H˽/���P���) ��N!���LW��0���O����i��Ɯ�>L,w�-�ʈ�p?�<EQr$nG���{ɘ�;��^mŮQ
(�X/�����+' ���M��Q�������لs�>��憎���tn��:k]�4��/���>�YEƮWI�^C�\�R��Jv$[�4�A��ݥ	�=�J��R��S���ڷ�t9$^9����c����B��G[CF3� v�T��l(.ao}4��P�G)�����J�8�u�]�����F��,�aL�<��>�{@yy-0�:%�@�P<�B������agAb�V��$*����C&�9q�YrY2W�Ϛ?^y�s����x�(@�ܑ�]���?r2��B̥3�`WOs�goD5���bs��<&�>��R�pP�2Pe�G����pG�純���.=�_kZ�^�D�@/S�Ⱦ���g�{��o��s��B���ÒBh�������֒Ȗ���@̂_:}�: -�$�A)�o�VE/E'`��Di(T��2��ϯw`KhUmm*O�������ꛜU�D�g�ӈ�t3�(<�P��r���+�D �y��b�Z �7�z2�K�+l4�@���i�+���%�+Z'��EG�f���P��o�h =��&��Y�'�ޓ��$�q��fv���2��,�	�39�ً˨�
���ٚ=�,:{a���������:�����
x9 =u�+����D�"�X"e������[ߩ���t�����n�+�p:x�wA�dy��ј��e[S�M"���8>s�Iz�&���ύq�ɳ�2�3�!�g����[+	�yN�+���xů�#�������ƻ[�(�{�^�.$��/^�_�xE��pN�f�U����+��{�z�)�M���u���S��V<�*|I
;������H���'hmO�=�r�����$�޷�ς��qO�t��J{Ӎg?x�����9����s1��0�LT}��R���~7ˍ�~��������	N��8x�2=N����<�<�p>k�)�S(-!q9#�<�׺��m�hB�c���g��*Kt�,�?��ͳ�E�Me�뤧H�M�3,�hͭ�=ؘ�,(�}�[ׄ�ܪdD���oKן��r
D��5��
5=H��Q�ӋN�[�d��N��@�����d�y�ls1v�����|��b��ڢ>�
s7�q�|�;�3Ɠ��'��i-5�$>��j����=���$t�_���l���Nͥ���b��}�1f��4/�*	��ċ��\=7_*�GXf8�bd�~9��Do����^��a�yL�����d�'�MH6�j��H;8g U&���BZ������L�O�D�zZE��{������q�G��$R�2u���Z\��Ŧ* �"!$)9ހ--8�|�z��({��b9����Ho���̍G�箳�
��)��~��fs��_[��@�t%ɷv�рQ)����	��h$WJ<+=K�C_�x�0[�j�%��<\�<�z�?�-Rͺ��]R��
�?���]��*�2�繽���m��*�)2z����+8���`=N���3�!�*�A�1l��\��8)|2ff�pвяK%u[���E�R��g���%nˡN�e6��勌��X���ݕ�8%JP�!s�|k��}���78��Y�=f�4>CI�	J��&�7э�J��P��<������4�D�Nn^5�Ҁ$�fK����"A�{�lM�/H��Ӟ�.����;;�`�*�QSX�8|��W���1�%0Yzrj�`�����"�B"�fS蟃�5�J��!r���53"}�4FV.M˅�%�`�fJ	�L1zP'�V�Sa��wVdUy.���7�0�'�Qؔo�\�bM�i'_��we���8��;two�T{�����5:�z\^=�#��=�Qs�S떔��
]#�>U~"��o��P?�]��Ib=�������m�X6���pa~�c[`#��h�&�t4_����ؐ�#)>�C/>�,r�?��/�	24Kw��� �0�d��Ƞ�
��.�&�^ҕ�PY�(�����Md�%��%y�eލ3FM#9{������ub�ux�%�!����ӹ�0��_�T������A������ظQ�Ŝfm��jv?^���f�,�^X��I,~ej��:��f]0�l�����>��-�}螝�ǒ��V�f����`e����E�Z��ʢ�k�#���b��F?q����@x��j���Wc��,]�ćüۼ�>�d���`IWt5�Ftn�y2%���[0�_�}g��h�-r��V�F�8�e){2H����*��.j�9z؂~�K�̞�����rd]�oo�"��qNξ=ݑ��I�v��~c��p���?��I)��πW��������:1�����A��5�A����������yoC��UTk�".��x�X�uf>�;#[F�k�g�v �ԕ7�?���ɰ$��t�EJ�����R�R�0B�� D	�1�Fb��ݽь�{������������u]��,r�c�-to�r`�-�+��%K��������׆nC��[ ��3JKKw�^0�e�>8	����tIC��U.iI�)0w�W�y%as����L�#O�,�,��H)6��R�sϫR*�G��;Wcuԅ��u/,�E�ȴ����Y&�;}���I��_w
w��g}u{/t�c�I�Ȁ�(���>&|`x:h�.f��Y�~w����?"l�v�qMj���.�s���R=.��p��U� �Ŝ�r*�(����;�Hoz�9�O��z_FkT�*Ro4�ғ���"�����P%��D{�l�E�A��E��" =i(o��&�ZN<`}Z���Ģ�&�����\�L遆&œ�<GE%W�e����%V�t׷o��t�/	�N�H~z�*�=�c�;��#������MлW�5{��7�����4��d�"g�O��� �3�*�t�h�+����Xzϖ����1���37�U?Z!7���.Z\H�{x�-�d����Qū��/`0���isoo�L��&��aMq�E�`uN‏����Մ��H�5ت�ŹʞF�l�h���[	�NC�(�d��P�%�~��o�$��ݽ�z���6������}��ʸ�n�\Oi�1U�5��/D���Q}X�B��2d2�E�΅��0+��.����j�������ܥ���v���q����X�����Ǜ|$qM- �'q܇�s�ta�u�'2p�Wz#7�Le��RUh���]Y)�(D��v���c[.aI��w���}f��`�7�z3p	����0�g�oD�&�0?��[J*BI
��IL�Tz5y�qC.s�颤�_�R�y��.��%��W�am�Gv��ҵ���~c��X�&G���+�{Q���c���ez8�ˎ�^[��+���1�!ɪ��h����Î� j�G�g��su�n74x���ޭ�!����l��/3fbǇ���J�tc�#-����t{ܟU�#���ٿ$e�\#���mk����rǙgEz��qD��;�OOBW�쭣7X+��dUg9��f&%�SX_�A�`���8 ;�)K���ȁ�<Wuou}O��H�z�.
5�a;o�̳�����BĦ5^S&K��nv$��h\��3�2.�NZ띒�("d��U�_/Y�����8ռ=���8�,�L�kE��&������N����t��kGG��P�W�D<o<��s�Vrk�[1^{���w~���>'�]����C�벨5�o#+��Sb�]�8�MCzl��	��i�V�k�����'+���K������9��3������WP|�&��/�땝gr]���`�[;�$;gfԸ�_���`�lR��=�FG����d�5�|9��֑ˇ� �ѹL�(�����#^k�߀�L��|$se"A0�$��=c\C~�uuą��1��ٙS�Z�/�M����rs"?�K�h���%��I��s�I�S�%��B��<j��N�AIV�E�[z�����Z�������"�;B�	dweq�|w�D��9پ�ЋYX��ż%]�۬x�y)���ꢤƷJL7w��`��{Į��`�� �,�+Y4��YY�gZ�@�T��Zaa!n��~��O����T-����|xX�7���=b�;�ڥ�h�`#�Z*�m��(��`�����N���17p�m!��Q)�q�g� R�㯏,£�ƀ�φ.�!8N0U��	���^(�m��\'�?�P���]c�h�����?\�|B����	g��ͭ�Ƨ��G��b�Ճ�y�Mw�O���y=��0"N�̫��Hk=�~]ҩ������I�;t,�cҫ�M���JiB&��H;�̕����`�a���"y�ƣg#g�k��1}�

�W�7�;ӎ��Y�͕�~0 �;��Yd��&⻯p�R��5�pq0Ѕ#^			��IW���L%��{E��z}B�.<B���cPd"C����������sq�@�9� �?T淰��b����Vt�+>K i��ȧT^���?�*+�/s�ژ��L�e)Yb9�苣�aH���ȣ��|��Pa��s��颣�J�;:v�$���t�DDg0���j;z�L�p͵��p��[���33��
@��Ą^��A�&u�������I�<ݻ����{x�g���I5�B��e��$��Ջ�<�Q���6]iR��`NH��$�J�x�����$����xjtַW��d����|���g��*ǂ4H�5E�Ip�k���ja+��&�k�G��W��`�¿�9��c�ůCD�_@��)�@���m�/ӟ�ݙA�VW�����>fD�����	<��.i퇹-ގ�P�`0X��Lq��K�g�?��R�Q��ǝK����lY�+�R{5v�aL���GHr^>7iP��L)Gb	 .�C�1��="]���:(涓o�>�I~GT���HҶb<�"J����o�:吨�����eP4$*��D��$8��R�<R@^iy�55t8��྅����$	ô7���Y���5�޼y��+nxb"�����p!΃323[��:�+�����M)�<�n�	��v\��R<���^��OK���h���j�:��Vt&��nI�b9���s�ŝ�נ�$�N�i�ެ�<��^����.�}�j:I˾^'N����z/�q0vM��y�(ztgG���$�3��n.;��2�~�vI3��	���C���ԗ%	�W����.�}o���#'�fz9�0Ш��-�ƥ��h[��;k�L���q(z2��8Z�����(u�!@ѵ�`�čj�ێ�6.?�50��b��,��uu�JD���<&��}�=��ZP���mm/z�i�����O�3N�H�`�L�݁�����	 4А���>�䥆�a�m9-P�M�+�oo�#���ԯ�)�m9b$Z��hgq���]�&)��܍g��y�O*���%s"�6�2u�a[ �a�.ۏ�e�Ɉ�������7!��s�Dh��N{��?1�[�YK��ޙ��$]dX'\�U��>�t����ר}���&tf�S�<�{�|Ձi4�L�����j9Qa�x���bp���YJ#��[�28;u��ݩ�� j����ׇ]��eŅoޜ�p͆m]c�N�'ai1I[ާRcK��� �^�����0V�L�{IZ>�q:jq]W�q�}�����N]��>�q�]
��fQ��M)ymM����.�CW��xYK�{k��^,��Y��K�}��`�����QʂH�D�����x�e	�����Prֻ�qI" S.)��>9.�Uۍe�����2�\��>p�P~\z?P4 ���t���� ��u#3�9��7�prb�G��AZ�_������H�?�?�4f��Ru�"��f��Y���￞���%$K/'���3�N3�/P�]�{�s���涤')�q��x	^��c����'}Ώ i�m�N.�,��@��A�Z�Ό35�m�[�]H�$G�r�X�0���TyE�����#1^��z$�~�ߣZT�٘�O�����G��ЯJ	0�@;�K��dK����#�&�Y�M�F��.j7n�_��P�PI�
O}{m��h<	�>�n<u����
zg�@C0}���Ks�(z����ZѪ�.&�߷�4�����3]��hd�h�k?��@�{_���ge���(�Q~��`�ԗ:s�e�C���@�
�6�_��J�i��񙮁4�������M�<�B��Q���#�p@�Їyܔ
 �Ē3Jb����H�ƞ%�5<<<��"���Pk��8J�^mRz��0"e?�J$ć��$�MEM��LD^��V�lv)�f3��V��fj�K�#p�����i}�jG��.��t�=
D�
���K���������)sF&��ϳh��^���~q�	���3����q�}�p�@[�UPPPf����\������D���o200�ʔ-3�"'�������P���p>�%M///�7TUU}��0j���e��N'|ϡ��d��¿�[�1}���@��v	����o2�=ԕ$g�ţ����gᄑ�R;���o^{�$�v%��T�DJ���6�}h8����:��7�<��؈�8�v Pꅖ�FP��钮*E>�:ύ��k��8���~��pV�Wӵ��ܱ��S�Ò��ܚ����S_�p�|[��2��/�Y����G��{���y2kx��xb����)���iӢ�������L��4�͑ۖ�7�~h�l�"�///ŝ�_d��>q�	��]����jҙ��j[Z�#X��-w�T�ۀ�&��s��"{�Do���m�Je����JU������օ|%��/r����WC^;�.�J K(��+���%����Jl��)1��������_q|zKy�Z��'nó�jl2w|w��<�,���-ǋ�b���&� �}�u��}y���c#���<��av������� �.v���ϴ�~�W~q0S>���=����k'c��߿_c�D��`Z<�Ԙ5�#q?��\snn�n`	s��n`svrx|���G�D"u��%lmm���ɳb
׃xĪ�	��u����(%��=�5�H�7U͒��˃�rv:����4Kpp(�$�����	��A�@3յ����O��@`ӕn� ��w;/�d�O�v��B�N���"�@��>~��bꍓ�#K���]K�=�w�b��}~V�ꥡ���^&4�pt�殕�nx�a��OW��:ʯ�:�$��2������i��g�d�,�>�e�b}���;���̶iY�J�^�-�
oy�!���e>�ܫ�v�9߳<��$�`k�V�?8�w��s�,���џ�'l�Q����?[���s�����{yM�	jW��d��R� �'���f�.����_��W���Z�5�\��OZ�����L�,�{�\�$y>0z��+x�ɪ���v��������`��`Y������S�5�ĚKK�(��R��{�G���3�v�:��`��7وSb��e!w�Z�V���O�{�lư[�沣���+d5��t�����/8H4v��T�E�	�+����/<rv騛D��mq����$8������ۑ􂝋�C33�11�m{��S���Z-�%j���⚛5�_�{xT���<�Y4ܫC�(P� YH6c��{�~k�.�����`#"���w�x�zw&�**�lS�o &�Iy�[�?���%{]u�r�j7j����q���-��y�񍏖�������%�&o16��Ck}@^�O;3���>��/@q�$	iA;�k����������4�ާ q��n3T¦��ۋ��$S��b�K����̪W�TGB�2�v,��oz��-�S�.=�?������H0j������O��Ĭ��s�]�㝹�o�W�n�R�؄� ǈ�zp� ���Q.����3��E����rvB��/-�����M��)©Ԇ����}r�>�'8��t%GI@�2ܒ�V��CR���ٷ��A�+�6�"�(1@|����|�����O��� q�ж���iFpI���0(�9=�?�  ���!�j�`�,R^4��``b��?Qe�^ڙ�}������]�
��(���744�y��TUW;��R%x�O������d���PܒK�^RcP?��6��h�Dk���Vdb~�q��է6��6a�h��K(dٲP�x��A?����r�OS���(]_޸8�����K��DoT����l�E*���gu>�7Rڝ!�b��X����~�䄿tO>X3=����f)��v��ɹA��˙��=�t�b�c���[�c��D��D}m��V ;�r����iX�e�g؍���##�DXn,9������D���c7ww�Ǝ��[�����C��(z����/Y{�8�=m7��f�%��wܧ�@OϚvy_,貾���릲�J�RZ�{��W�KE/�뿲����G�P<etv��$��fb�V1}(���m�R �:�L	kF9[ x5�b��psE��0��.�ʍ1�ض1Qx��!�w���܋�����q/�-1�c���9{�"��������2�&qO)f�=��S�\�<�"��m��	B�pw��XYYu�l�V���t��j$��)��cr��~Lf�s��-ҕ7����K3�Þi�!h��RE�Q��H��l7:��-���Zk
_�/�����>�Ը���A������y#���Y=�}���1��B$��鄹�L��lI �'#`�ORMԍ�
J�a�ʂ���vn��vJ�F���$��J�K��/3n��֦!��J�ɣA��$�~g��㿍@y��<��Q�7�p�5!RL��7��X�Tp�׫�|�Q�n`��ϧ�[����Ɲ��P�����v�8��W9�T(3-����m\0�OT$����r�����K.'��$?����%8�����/��Tˤ��R8�-�4�9&���o�6��A{�U�S}���T��W�0�2��N����r�O�s�_���P����^!G�?�݈�t��iQ��,�Ey�
jx0�2\i�"F!���l���/]��`��#&-��`ebaA����'��q�yW���qW,�Z�Y GFn�-��Fσ��!�`���ũ����vv|	�z55O_}n7�Y�5ITΘٹ��,�y���@�l;ۧ7�o�h��l�Ȓh9�啙k��څ�q����7�7m:#Ѻ���3��Aj�H�����uC�b!'Atx}xQ���؎�]΅��eex�MG���`�38]�iv#"u�~㾔�4_�m�X���w��[���3'V�u�O��D�3�eƿ�9$sM4kx2 4F�\�>"�pF9�x�������<j��[Y��<�Fb'��Y�4�P�#����{�cc: ��a�Y�ō@2�����w	���Qs��xx��)4��aܠP���`܍'��^-f)F�9-�YI��2 ���!�s����A��98&^�j�v�3��T,�\�vy�f�[��o@��_�y�$�(��з�]k�rB���G�g�dսl�z�an��;���x�4� Z��Ms��x*�V|�썄W�/�ˌ[�5���<�{��%j�fP�?MG�v���N�bbGǗ���^p������PiR�--�)�>LKKK��c���N����)�� j�����wB}q~I�K8\R��`���9d}=#n��ή���`hr�g;9cn`� ���pD�� ��)�J�,u������S�V�Y�VR(~gu'���W%���@K��$�y����M*�?W"�g�+�*�\"6^�Y��{.m���ʟ���fLN��b<*���o��d~M�3�p�9�����o�]��L��]p=|��K�ϴ*N�~϶�<Y���7~�$�:�~V�R?;?�j`Pbrx}!�E�&��oT��s�1���0������UT/��N�x������ַ����Xs''ʶ�6V֎�Aʐ��<EvI(555�G
4�������H���4�'aU
�RK �����ݖ���=�}�N4ų~��Na6�q#v1�v�[�zҜ�u�����S�')XR����z���r��3ukx8Ť�o(��Փ8Y#zH�ɝ��wz p.���[�1��B~+A���A�Y��3����zw㿽5H�,���������cL��fmW+�{VP�8Vvv�BQ=N5O���\��֖��߿I�ɭ��4�]]��{{�m����o��wW�_;N�7���������L��C��agg^O�<� �ITT��h[;;܏FGG�lRG�g6}e��I[t�=���S��u��|�� �A<|�4&`�nM~^>�Nà)�v�/j��04u��\:!�t����Wo�6���9����!xyZW@7���֍���b��RC�&ҹ�V4���3av�� ��s/��1~���Pwd"RT�_�u�Ay�q_���,Z�����rb�9�R����w~���n���X�	uf'��f��.��/��U�����l��{�����}a`g�g���5��͍&;;����p	?y��9a�|�㮤��p>|4!�XvNNμTMUUFv���������I�0k����W�2{Bb���5�C�w��\�C����Ip#�dP�)��������27��I���Q����i8a���%�,�Ʃ�dt���B��`|{o����ob9��>����Ǔj�I*��A�M�J��� ��Y��Z�}�j�2�_�6A�w�5/A�Z��.�`����������{��k� |��1�������T����x.�e���=3�}�n�ck������^����6�mn���S� ��/3\�q�>L[v�ل61���5��ÏO���y��B����&I4����o�����Mݐs�M�`�_�:�B��~����eT�;^�%W�}-x���0������L~�N���rCc���L���b�.Z���^��b��M?j�L}�M� }l�p����F	�c���)�|��H�Ph�8Qm���	��{��g�R���L7�O���̓;u�� ����[  �����(���v��	���\�4I����V��%t[�z�Rzy�൜��ȝp ���L}|� �V��)�231��T����K�|O��n����2X�gb�R�hV��*�1ڦЃ���TZ[k��ϖ�f���b].�Y��$���I�D���'�4%r��:OF�����GY�UR�����(7��#Z���xCf�[i2�D�^!Dhy]祊2�q�@R�0���ev��v�M��x�� "4ѧ_�wc߽�"XV��Q>�9؉Vg�Y��K�r��օȿ=�+䙠n��3���h�g z<"����-Ƈ��ڰ)�*�1b��{�6bNuk2h�ޥĜ��1�I.�.@�2[�/�17�eB���S"Ω�Z�n�;�H�آ+����W��X�U��eF����+.Z�*ff��6̍T�ۅ�$�)��cܑS{��r�i�;)��y�3�Ky����BwG�����#�i�2�Cp�i� ^�\oU�r�q(�K3E{�n�?�����"�G#s��.
�g��;�
�� S�h�mV��5�ev/v�)�eP����hR���ڃ��Q��-��gRN���G��M8��Y/qGrWGYڋ����Q���iVaֱ4����^C2ˎ��A�*��"�Ww�2��-up����,L�u0+!!x�z��B��-z�^o�*4�r�R'�9o����D�g�怯�*�}�i&��[�ۄ�\�o��������3�z	ѭ_U�M�Tl���Op��F��^Z�����LU�u�5\��_,H\,St\2�d��t8�Y!�<���3����/�������~<�?���D^�Er�d0�C�h���}��o86-_SJ(W3�0������z2�f�
�R�L��c�� KjJ�w�C�EWz^g��-K�t`k���X�N�����d G����}��"��ڦT ��?]��#�+s]��Ƥ8L��#6
��'��p{)�ݎ�j�v�]��b
3)�V�O6G���O��ud8�<���gb���fa)kM���R;�mq����-�Q8�Ӕc�>d���f��a�(�I�Zv�c�^�<`���큺�W��N�Y�2Vo#��V���뭊�3��
=	?�O����a���:ϢP��y�E�.Õ�8t�>�;��1�{�-k����-6�cAq����򞎕m�*����l��Z�Ɯf�Ŷ��!x݃G�UA(��;n�"AC�����Ût��u�"3%İ�����/�'+��j[^���&��%�]��4�����^Dl�r~Uo�r�-d��)Q�����bgI��I�1�چq�g�i/���E+nK��W_ �@ɢ�̴�z� Y�}��	��n(��=��E�%rn4L�������Փ��f�.�0�G_�8���?��O>}~1Fr9v���~��A<w#=�<�l̲�݂
�9�ŐQ�a	�tzAE�x�6G�u7L	�<��o�4N�z�9k�� �Bf+k� uիUk��z�Ս��瘸��׫eKH̦?��Y>�O��c�/BpGŠIak�w>)������8b��Χ�?��ç��� ���6	a��;4YZ���ְ�ٴ������}n��EpT��R����8(u�
���<���,��Z��`����Tʇ���9��nJ��I�C>��x.�{�*�,��8�W��X$��ίmV�#Pv��c�C��z\M�5�@f�{��\ʓdr.r?�%�U��#O�����-�6�OzRT]�&�-�i�+��O�(w���vA��z�K����[����碌��I�'�Y��Fr�-�W��[1ϳ�SM�GjȦ<��̈́s�A�"�l
4K�1���S�֒�fFj[�+l���I��R��Ty6���{e��|��3�e3��-��T%�������7<3��Ŗ&o�������>'2;���
ӱ��n#Kg*���3*�kv6��E�RyWy)G]�Rj6K�Fސxh?0���?{�JҰ%�`r|�2~�lNX��G�Z��$R�i���g��ih�0d�ȓ���IOy���0M�q�F�����eȆ\&� {ɗ�ٷ�j#��p6���0w�Mn�#�z�&!�:����,
�G�;�T��_� X��i�톇QϚ�.�@p� �8|���,�Z�v=���C�St]��. ݀]�|7F(�ܣ<�2�/ ���2���w���6�Q�܉{��Ơ��g�=ρe�<d�f�,�Na�.�\J\��4�s�|I&p2��]_EQC���1E�*�����]��EIt���I�QB���i�M�O#��eRj���}
s��>���Z;DJ���0K�(K�E�L��O���\��7�`��\��
I���8�E�=0��	G�w��|kQ����i�y���ʗ
h(��h��İ[�N�@�t	�/XH��.�����h��g�z�`��U��u�$��T�q��3BK��#g�I�`��ƩǂV�)�!q@��ئ���kN��=N�x}�sr)r��K+!���&[/�p�?��6�D�)с�,�M�f�͍U%�( �`�E���+:����`4���B���������%�zUʷW�i��in��D#)N��x�h#�uFk����x8��*ulIg���/�?���� _$�L���w�d�8����S��f&F>'�|>��ǃ;$���?��N&�
drS��~,�i�٩4j�i��o(�������	��*���/�FR����k��0��-Q\Z9+�2��q����!��3];ǵ���pD��U
�7��3�T���E�����X��|��V�W����3����{�H��-�+��tڑ�EfhB���1�D�eW�ƭ'e=gH�qI�?4���>}�}>�n�Uƛ�[�����e����]��/�M�~�����fu��׾h���Y�a���jՇ O��<f�<( X�`�zs��8N!D�,�]��>c���c�����#�b�I!�(��~�C��Q��������$<dUgV�|Wʓ�qH�%��u��GX���}�ϲP�Y�>Gꃝ8����g�4�z_L뼲H���^�x�7`V�o�*Q�!�ؘB/���8 -�nXq�Eg���c�ok/�nSu2ɸ���QC��Ee����&t�&���T%;���>8$�@gAV�=o�Gj��L��g4R*(���=���Q��k��s���u����+�<WǷ캢�袿u��:/��w�A�Ѿw&���s��nCL��޷��L�m���*��P�l�^�����(�)���%����ͬ��e9LT�4ʇpH�}x�'O�u}�e�I��S��Sy�HO��d ߬,���븡j)�}�-&�V7.(�'\�x�N�>٢{8t������k��u�>��X����La�y�RZ��TQ:�A����լ��b�l�r������Ѥҵ��I-���@���K� tAAE������'��M�@ �T��ؚt�R{�9Lk���U8�j��E6G�ף�S�Ҙsa|��C���D���P{��򩓬A�-g�-'���=u�a���}�%y�XϢC��,��s)	d&ݝ\fwYD��c�a2=��Œ#x��%�c<����g����no��ӮE����;ʻ�78���W �Y��a��}�yZ���.Y�^��7A�B�HٱST+�A�QT�1v��{��
��f_�t�Y�M�P�������.S��	yF��D�LH���޷C=��\��:��0M@�f�]ǌ�XD�p��O�@B�I7�r��<u$u��[ʾ���=�>�K���)'w<�#���6�^�cΟ��������Z��?	���F��
�&l�J�ަ��<o��i�aW�Y$�a�Iԍ�%���W[wI�;��j�D��e��V�o�o��C�7+��/��R=�~P)�����^�Za�{����KE�QY�~���l%R�P�H]X�W|�88 �4K�}{}JF�Pʭ�����p}��-6�pm�[s|�e��*j�4"��� �Ir��Ii���	9�)׈�y�M`B.��gq�z&�{����f�;uP�8�=-��"W%�}I��ӛ��s��p!�hST��5�M��Y�w�3�f9D�%�z���{<������'}Hf��|Bغ��=>��R�MN��ǡ�y2�#���+�A� k�	߄`T�)��ל�?���Gi��2\b�^��{l.�S�W{�y���ԑ�Ng��Tz+�,������ץ�Iн3/Rxޠ�q�A����=�����[֕%
|\��ꤝ&N�	7�ڦ�X2�u�o+��U�/�re5����n�i-���v=<�-��j@�Z��$�&�W�4B)�����MtȹG;�e�1���3Zyo��#��$�>�^���<v~pj�&�����_�f
�**�����6�ŭ�W��lF��^<�[z�~�xU��\�c�8=��hz������͒~�p�����&�����7�]�i��zA�l��7S�`g�U��k��,���J�Z��w�	�E[I�|M��[���S
�2WiWg�d5�Z��P���۪���[Sz*�U��l�Sޣ5�$����9P����+��,�2�}�;|���wb�AdIш��S,�m��w��N��-���\���ue<���+w�I�Q{Q�%+]W���A��Qe�w�}�@�8zv=�qjG}���w��V;j���(屖uQ)������������~�"s�ș1�6���"2�Q�{�z�$�[x�I���Gg�3�����+(�l�9i���'�s���xNɎ%�3 }��{�Ǘ�RҬ��5]W�����Yz��Ӽ�q9�=����^"JwE�-�(k�%M��#in��O��!q����q�G_��E7�CXJ��6�f��ϳ�F������vG�L�wţ��Wo�xwPՈu����G�6��p������;y�*��O׽
E!�y fl��و8cN��������N�F�����>}i�WR�JZ��@4��`��xp�C==�`u��g��E�U�Q��N�|�ƅ3ޫ�xl�+`c����x8S/�UEc��9.����� ��H�fg��L�z�!��bh.kBݡQ�/⎣{����;�L<Dm.\�X�XP�#KIZz&| ���9:c����A���&G훫�2^,+X��]f���E���ހξ�N��<Ҷ���^�
�����V_��%�<��^R� 5$�,�O&D>�m�st���Y�%�`t��W�S�P{�cC�|^�Ig���k���?8
���~z�`)���J��W��R ��^l�<����)�5c����M�;fN���/�ܧ"Dw[-�?r@/*|�It@�~G��T_��v�J�4�瞗3c|�1J4�NS�[N��W��hz���_jӱ�u?�rIe���^�6�k��o�9=��j�r�ķSK64ǉS�(P�cu�Q$Z�%ŽTmR鴢2f��K9��?�!��!A���|3Su�dō�w�7�~��oz+��~y�{H�t�<+��C�����-���q$k5�O������][ge���R�Bk|#����
�:IN�쭣��ma�{��!�~VN�Th�~%-0�ƹƴ^7/c��<o�`S+��L@��W�O�P����f1r@4jI��M��E�˸\���7F\��g�s�0%��!n�piK:!�@<�*W�:�2ڲV��Z�Dh�h�G��EhV�m险�?����%������7���CG�|
�j�A,�>���yp����S�p�����.���ڌ��Bi>��C,[����F\z�n$����
W�yD�bIhz�uӵ�ۼ��w{BA	��>׻��� s��5��c����O{��L��b�ڹ w�HRs뇹{�>��1�]'A̛��O��>��=2G]o��]naO��J�ٯ�[��&��pyd���) �.~���.����s��w�˺��e"u�7JRd���������t(;���%��zc��Vn�qd;���p}���$���#M���|)9D���|�u>ҋ���$�ն�)���<i�x�_��-/�R��Y������j�_��>�g�%�u츊a��V�uUg5�hSXDZ�"��̤�����xM@;®�d��\t=���VZ6���b��9��N��/��U/GІ���#W@~��U��z+�2Z���3c��w����`�X�@q?)Y�9%*{�hY��v��+q��>��o�3�ܢR����FW��b�!#�.���꥛�*�>G+�n�~���zf����S"�Ց��ZӛnMu�2�K{���d������0��eS�JOQ��U��e����JG�|B��d�����8�ki#�V��P��/�b�y'�HX
�vq�����������?4�W87�Aj{��'��d�w��ô�;!E'���i�)nЧ�x����m��I��%��s�NR�JV5��!�����ԙ�U3�ɹ[����[�XK��I�h}�@����%��}�6�sz�_�Lc����O;�-�(�.X;�8����9x�z9�ؚ,�2�ݿ�(��ޓ�B������4����P!oE�9�\ٰ��ii�d�������!x����Y�h5C	$b���Ч���8�&��b�p�4/�h/\҃VumNR��IU�K�\.m%�V�����1'��D��I#췜qW�ʵ�j5��/�w��'0k5��E��8zd�Oa��x� ۍg?�yI�"y�u�,���O~VV����`R�,��l��f�f�mo@���"�����l�p���_�|D�[R�4�ɨ��� |Ơ[% ��C�>GP�@=ݖ4�}�n�U_Hq���,��/�e.t�������:D�����d�$�Ąe�q�������[\����}�����k���2Jo�Df�J�ٯ���u\�=�<�����:��:n]�.88ː�8%��M�1�p��(��ϊ�Ua����=ü>����l�J4�i�7�&}�>h2}/����� ����fbd�e���ܡ��r�MHV�[>����[X'D��%��^�e���{��.U�>e��?Dy�p"�2
�B��� d�Fz,���.�TY�<ϸ;�DC���GW_J�čc�>H�Y$�$с�r
{���*P�QA�p���3���L���)����#���g�S,�y�4L�H��&7lO��HV�ũ*q����� �*&6"��$C_��R#�=nHY�}%����uB8�v� �@u������?�tB����ѺAs��f�+��^�HWj�3֏}�r�Q�E+�Dt�p8.s��q�@�c����8���x4�4qwZZ�K������)O�u~��)uL���F������� �]ze�K6���?����lw���e`�V����Њі��t�F�iq�"�_h+����:&��/��j�`ῐ����?I�P)�Պ0^�Rv�� n3X�r��o�ny�!&z��|����M�*�|��m��V�[�q#��|� 1��#���Xc���ms!��h�<>�* �:C^�)S����x7x����/t�KA!��	�(.6���i���ރF�9���ϳ�O���gL7��}�"u�'�[Ѝ�Lb�E�[�k64��?���O�j#����roX��$��o�M�㱯�w��r�H���T%p}bD�VO een������O/Y&�nr��?뎸�D��΅0�{�o�㰬_	U�Ǖ�p�ӄ�R����w�{A�ܶ��)E���jE��j�����x�ӒR�K��6��3p��*��̫�e:��\�[��3��T�bz����[�%����C|íO
�Qϐ�����b0����\2���(Y���<#>�V�8Y$��X��E����N�`�� fy�4u�x�<*��y� �!H�2�ϧ�'�W�����C�N]v)DԮg�ٙ�ѧrSN�QlfI\�"Hy�<�|��G�;����	����ra�-\�����J�S�Zw��;���-��m,xZt�`�3�ɴcJ��]��5lF=(������ʧT�R��������;�ex�
�"GO�Ai֬^�R����R���	�90�и����4���Ad#�P�Km�~ �JfXF��!)(<Uhg��P�L�ڍ�Q�kWŇ���[���N.�v3��\`.Ckn��R�������5C
>߹:0��wT����ϻ�0@�q5���~w���0O�d5��埅��ֺ%���9_���{@8g-O,1nS>sR�>��Ѕ�Ee �P���23}�:�|)��1�нO��h��Y�m}�I�l�`��
��E�Te��~�g�W����ꭣ���7P�iAT�Ni�����n$�A����CAJi�a�B������]��yך�X�����~�}�9�,_|�;vȔ]�ؽ��G�&�t�v��f�V���3^�����v,�r�xo=�-�i��һ��n?���B���B�H����@;�ү.�T�>�O��Ɇ�9�n�K�2f�$W+�*�>�	�fQ\=��R'�(�M�\I��η���v�h�<��Ag0+Zs֔hCXw�1b�?�@n�{�vv� <�y<i��ѺN�"+�!v��r�!���lk�p@��7�Q���E�k�=��ƿ��L@�H3ߌМO��FwH���^R��CN�#nn"�%wt�=����o@�-����}�k[�o5>�<���?|^^��H|��ap+�!K��2m҆�y�d�~M�Ē��+Ih�.d&��<��7���+�c�b���?G��]�
.���:��u�3�s�K3��q�dd$4]I���ϋo^=듹��}Hf�Y���?���H_ϗI"j�����`@Tc��񈅘3�M$�m�1��=���! �a@�u	f{��G�]�
R���}96���i���sQ B(���\�߈�LC��w0�7�u
 i�V��\�+�8mw:���揣�|�Ԟ��bXh!���k�=V�O�9���V��k�v�e����-�I���(Y��>6���,A���F^�����C��!���R�����'���'#�W�"+�ْ���b\�}$��d������VH���~S�b����iFş�4�h��Ӗd٣�69���.�gu��Z��D�ц��,�=�jrw��.��]cL��u4eY.�[�D4���K�+8`��wI����4ŉ�Y^�.�s���$
�K��o��}û�=?	a����50����"�
���$�!�����f��K�l�?�IВMm��F
��?���4�t��Z�-�d��.lP��{�ȖT4dg��{y�3������v�����o����R`�L&�˗R����/u$fj��-����Jɯ[�u�7�i� ����g��͡7Gh��.l��A�������߲�����Y#���S����(�����`d�-[�j�Nڑ�t'.��Vҹ������)qj�����pw1+�3���z�	΅��Byl��~���3\%qEw}��G���(���,Um-r>��BH��P&d�2����@�����8]��J����S���lw�/ڎ��H`�˳�^F���׆����������}�7j.�R�H���a����L	�vr�k��Jf��EJ�̱LŲMN�rjcz���)���. [��d���^R�K5�6ms��W�Mڴ����D��~�jmB7��(kBA��?�K`��a3�o� ��bC�L;���ܒ`�t��E����0�]D�n��}�{4� 7�#�a��ɩ%�T�!��!5�Pk�1"���)h����C�pZ^�Ʌ��p���d�OV'n��5ǋ�xOM^秵&��&���u�����X@�u�sg�>M�A`u������&�X]7�������I��r��U(�y����8-9�Qf�4<��-4�V�=��L)�%�]�xQw�H���i>�I��y�Ö%�$�W�u� ����`���
�����8y�{Q���҃U��<�̘;��sꁟG�tZѿ�����O��;6�0ި� !�;�wH�<�m4��.֬��nˣכ2~Jg`Y��@�ö
Kx���ϕ@�W:-�9U�{�1���_V�:��^КA?�j�=��$�/�1n��K��3oAZ*�QX�\�������/���J�����}��t
p*O�&�ҩ'���!0���H�ےc+8�NI�����;V�ms(F�S�r�R
h�m�zR�!H���~��ZJO���>�� �ݺ��Gǵ"��lgK�H~(������(���x�Gw��A����!�1J�sD��3j��IҬ߬�Q���U���r8O��z�^�{XR���Z���Zh��0��{�#�e����P�6o'	}�;�`/��j�yL�I	Y]�Ә�h0z�)�I�E�������x䤪�E�c�14!ݣ���n�p���(qU��9�56�t����"� A�w�������}iԢ-e�-���?2F����!^ǟ,�4U��j�l�M����^�S���V&:�V�D�����a����5H��~��v�H�LG,��>$?��,5e'�t2�N�/�m��@[����:��lk\lc�d�-��N�^����� [�<��Tv�w�g����Q��$�?�i��'J�0|����P&E������j.Y6��J�����^�J��Si�2���+� Ф�'��D|��ܹ��z���úN_ƛz���j�>A6x?��8��nxӺ���vH]� �Zv{����/�&�b���a���D-�3]#���xa��x(�3�X3`��Y����n(�$]8��;!Oֻk&G�)?yx�c=܎���?�C���wY������ag#�,��xz�M��&�QW?��%��6�J�]���w�\��(��`zu���{��y������Z�8�c����-R�Ӕ���ݔ��z����:�F�!g��!D`��&�!�(Ύ�F�#u|�; ��	�/VT	N�g��4&����Q��(ѕx�'2�3z�#ch�Q�䵼��J{
���w�mA Lg���I����J#��L�c�o���#�׾,k�Y�źq�{2�Ɂ�����z���>e��</ol�{� ��eq�t�|<��Un���T�Πz�*�ek�4��roa�mj9�\p�c]����2�W5Y�m���Dw�d���$|9g��]���/w��>�?�Ń�	]�V}�+�D���Ÿa���6���:�1Hl��'�h��@��3]c/eY�_���5��k���V$�(lA]��O/1-�����-�����b �<�����3��X5�:�:k�3ep�%5���}�ɿCn�S�;&9�ߡ��2�O��oi�6�����t����Gfp��.�[�gAa��s��������"o���_���F�<�>�gU�J�v"j����
,��d�*�R8=��k�6����g
N�^|���[�5&i�b=���z=���ƣ����X�$�	���_��Ҟ��I�~b�W�{p5�lK�ys"aruP�!?����l7&)6Ң����)"�=�7��47�~����\�����"��ގm����ZC7�ϖ�׿Nc�3�!7ߙ��e���9%U^_��ɊȄ�<ޔP�+�֟�o��S�g%I������3Z���GT(~�I}��?N�ؕ�R�?̚��栫ߨfwJ���Nt-����{�J{E1PCot&^���$��o�b1Y�n1������wx����==��X^��7O
«��9�b��6��V��}�n[z>Ps�`�Փ��l2P��J��
�J{n��@��q���ܛ�F��F�P��H���
~ .,�)�s���j1��n3�d�J1˖�*�匏m2�;b�f��V󟗺����h�������ˮ��
@�3���Y�dJ�$����t#DD��OmO�b��X�j��~�r.o#*�	giz7D\ra�������:�����������Z�F:U��ʊ���M�|�Ws���:�!w.g�Z�ۺ�
�1�)Sx���a��?h5F^ D���7�X]P��#)h������i�1^I0�$$4�dY��k�vp�>�Y�FLy��] j���W���>��=)y�q~GSL'�Gmqvt�st��"�C�����C���`	?�i6,�I��󛲪���A)C�I�>�
����eFW���i/̜=,�)�����fݬ��쾮�fP��F��b��#�^X��;=�M\������`2x�[�$���4�{#5A����������2�.I����2U=5�Ͽ����e�:� Q�ok'm=��n�_Z���pj�1 a�:U%}�Щ*�I��5�~UvD�5��|�'��G�
���OLrf���=�.����ZJP#X���b��Zyu ������{z��>	ʃ��ոG?L�G-Z�H)��i����AS�Ύ�d��C�G��dU�}�1B�|<��	N�+X#�&㉤��}K�� �\گ�_2��w��]~v��3��q��ӳ'k��yT�'[W[O�:r}7�� e�u�2y��/�.�l
@������.a}�]���Ao���n�4d�S;��*�4̝���>@pN���y`	���5r�O*����t�{y� hI��?i����$���D����n\`��=�2+��/g�^��n\aoi;~�_��Fd��^�	�G���ꄰ�p��Ə1ׁ����9r&��̺_1 Cﲢ��
&v�L(	@L.���%W�13���w>ZO���9��(DK���"7&�i@���ܿNys�fj�w ��(��g�rnd�R����8��:��������>�J ��Zh���h�Di��ӊ=T�7J�{��.�(jV�K$��!���`��������3"�.o�"~����ڤI���vlN���|�0Gz���R��:���w��00���@'�,���!g��ى�-�TI?�l�����s���O��0�:�F�����Ze���_+�q�K���WM,ڮ\�5�ׁ0:yå0���Vͳ�%��Gã��$qJ��x��]?��I� �^�_�+pt
!d�ͱH<����	�W{�3iRS�/uq���F��u���%��(SNJ
gB��-N���y+�}f}�zM�Pm�6S��n( �Ϣ���+�i*��g7�� U��d��(���/�=5� �WJ���kp5����K,I�+�׈s=?]�Ճ�z�q��qbF?���;��3)YpEk�p3B��ތMR{�:��d3�x�,?�����s�@���Z�aw�mwh=ȡ���!���V)���`Zntt-��Ώ5�fw>������o���4lm..6bBjQ��ܔa�9rt@�x�d��ۋ[wlOY3�l���5���7�
���h�Ǉ7�p�������r��?͹O]H8VO���vb����W-��L:�*�oT���0�,��W��ߘE,{5FF����<e#j���P��>�5.U-�������g����1���@�{ZMp���f\��d4٧���y>�J1/I_P�D�1z�����m�~j�H"N3�q�t>Q��ѕ��5b,Dkʄxy�ɓ���똌�#�ǡ���t��"�(�~տ:mxE�MH7��=����Qt��ѝ=͆2nD��QKɆ=�1�UKör�'��qJ���
8�Si����*t$o�s��:�~�֥N�S��4d�p�xD�A�|�}�W����W������':�E���FA	��o݅v����{~�K���z��#�(]�J��x�t��	e�P��~�B��BP��Y�9Hj7V��x6*g'���\����>�U�}��5����_���<v��סZs�ڂ�T)+L�AM�~PH��/�����u։�j��y�?��Pb�=0 �L ��G���k�������TsR�t�p��X0a'�}��4I��T�|ND<i�7��Fo��������|7�S�y��?)�$�mk��R�L��Z��)���z/S�o����8'X��G�6'�SQ2Ň�iy�ks�S��&���Ƌ�߈|�v�3��{p�x2�,Z�/s�8����b�Z�9!��\N��������:{�s���~��⹘6���2��&N�{T�Ē	��hV"�W�}���r�HV9Z�$�*��yֿ���� �Q�j��I{���z\��%H�Wx-�7�wLKV���4��8bQ�j�L�<J1rq�o��<�d�\_¥������i@�����#2���"��Jj���]a�%���ցB�Bȍ��K�E�%�/3�a��E���뎌�ж�ݻ/G�m.�yA����?� щFD%�]Z"�mda���P���"*$`<�� �;�9m|In;�1�{�5�&F�Ys�M[8��x¸���ސ�1��}z���s2ȶ)jcfQ:"�=�]~[��!��];���d������?��l��.�����*���H����a�����ݸ"����<�,��s��V�\���oO(�=¹��,)��J} q�2o�����>9�)�|BA^����cjW�xC(�æNAa_���md �_ZS�����|�j���d�|�(�=��6M��!_W�o��ۜ�a��@՞�׋�෠�bv�`�Q��_--#K���9\dt�j/U;j�Z3F���]�����o_E���A[�FQz=�&��[r.7�9�\kG
�A������:X�`��~����8�g� J qx���X�J�nb�_*0aU�m��3?_I����,s�I5ͼV�z;����^��3)�x��s�V��K� �Z��?I���.!b;���+�k�R"�w�jċ����	��I'L�)5ZT�0�F��=�Fy�����o'���������� �(SB���D�##�;T}��v~���P���̹��/�������U���&�J�^�ނ��?� �.q�Ʈ���>�)G[�ϻ����LGke���q����\�ӍSϔ#X�1�U�Xr�1�Fɱ�:`\nx_Va�b�̇��􊻲~��i�����!��(%>���o3#X��ʙ)���jז�����߄�[�wtg9U�}����.w'ؘ]����27w��(5�w�缀_7�U��O���h��a��m#���ϕ��̖qjG@��a�,����#���>���A�v�BO@L�dV�sl��º��q!��z�wI}����3l#$G,�8�{,�����o@8c3��A�?�����[�[�m�_n\�oJ�7�S�>��[�N=�!氏��iq��Z�%a�Vh�����&d�^�P�[��HF�%�f�cV��2��E�N���c��V6p/������l�a���[�/��a����������[	2�ka��k��f��;�j<s�E�}G�k�"sj�C��#��q�L7Ă���Ѱ���o��� ~QdC;L��w�f󏆍@ ���1r?r:AH�rCa�C;8�%�'�h�L�L����{*��o�@Dt�Ies���l�:�}�9�"�$h��t�NwRXZI���$�cv��ч����I�5͍��s9�B�~��m������O���I�Z&ݢ��v�U�Շm���[A	�0ha�8@���t��r�4�!6)g�L���bNyA�֝�/�s��^��ү|O�� ��L��*=�4t|��j* ���RxN*uŒ���}Q���봞*� ���v���mZ����v��ݦrM���U��f�1�����X'}��V��Eh��8Z��d��Q�Cf !���G�4��߷�`� ��R�{R=�FVv~7����|0Y��gEU���H$"ǡd�,��Cק(�74�b�듇+���>&7�IZ�MvZ��ڣ����������!�F�I'm�2Sﻡ��&�w�g�kL�I�����%X���װ �h~d�s�����H�מO�7*�a�?���YV�rw��8�����7i�s6�E �j��4���8fh)��Οz��׳s�p[����\�u�Pa;-���X	ZX�6	<�*C����H���U�	����-a+�A��H�@ta�E�n�ud ��z�=D]+�u���^<b�%��n�
\t�_ܛ�@�f����:���O�[9������-�m���su�B�TO .E:)�OIP+�G$S�����`/m-�I�r��'v͈��ڍ��� ��D]�Y�D� �Z�v��_P݀Y�cCr��g_�&�#L�8��'�>��A��oL?"gE�ť6q�N���9C����e�����ц?)���.���S�"��96f���;[vA�/�IF�����D8e-w��9���:����O~��ۋRL~g#��XO
0���i�y�RW��	�hV�ӭ
�:���{���}L����`��4�HI-ڭ�1[��օT�l�J�#�2�X�v�#��z���`B�6����D-���!Hi��ɧo�f1_r`�����U@j&M�YZ�nٳ
�'�3#
[���p��8E��bT�o��f��ƌJ����c}��O�Z�b�T��HK��E�8�N��ZA�&cu 2 ���FL6v)_GF$-�� ~D�8߿��~j���Ů>d�9����⮡8S<��3w�~=SK�	�.���Oe���X����oĽAb	H��x�J��;�N������)�ݢL��u�_d_�*x�(ĝ~�f���J�Ƚj^�N�,��Ci�o����S�#�f9UX�e<2�����`�طIe��.���x�x�<��L�iz��;�C7�g�ZN�Yo�0J�Ț�P���*Y���I�>:���ju���M����t�������|��)&�w:L1{.?����׃���J���S�_�j���il��c,�I)	��Ӝ@n'?Q�6��(�N�g��ACw�M�ly?�3wûQ�fT\�����h��T��O"y]�"��⫷�=�m�I��`�1e��m�oh�7�W��*�`���a�?��>��{Ya�6x�msSz̵V$�'�u?�;����w(�
(�hν�[s鶒D0pk>�2�j�[13�E�%1�qN�zU��Z5����U �)�Jg�K̳@�An��`�ޖ�:p~eX_Y�Q5��_�y���>kEn���&n!\�]��l���G�xU$��3*	����5��!��~U����q],B��n�釘�4�n����Jy�ދ�W��i�i�{%���J�[�,)0���Vꨇ��8�bi��8�JZj�O��&:��z��;��Y�)=΢�z8�\��f7��������\���'��I}�'�Ļ1����P`�7QL%v_�@{��{� -`N�G�0���}rϽ^4���q^9%M��]�q��ܓ�XHmPI����[�(�[�L�<���^�䮊ܓK�)�<�]-K]�߻Or%D1�')����:����;\�4���eS����`f/Zvx�B��N�����1!��B�5>���_�y��o~�\����^�.�SQ�JFT�M�#Cd�6����I�T���%N{S�A�4��C��rX+"@M���q�{'s�Dw_,n*`�?��-X���8�ͻ0�e��ۈ�ܖŉS��Kqq�8�j��l���
�à<�F�ԙ���pE�NP��I\�Waקt]��4��+��R��I4�勆.�����hN�8�~����Ĺ��I�4l���x���Z|��/��@#�W�q+�&U+t\�Y���� n�K5��jՐ�6gS��0�N�]"Џ�hգ��!vU;����i�*�0�9�c-�	��\�S�W��%�p�?�z,�8��Ҭ����W+���P<I��ȕ 4�,d�_�5 k��-Ε�i�@0��	"�OT�*[Si䜁G���j�	���%�AE-��Em���E��"O?hB��Q�.�虜v�` h�)~�ôፂ+�#
T�h�`eڭ��CV�h��C��,��,�����׬R���7d��%��?��q-�>�u����$��<)��G�;�8���H:�c/>,�+�減F�KUf�D�3�\q�_5�p,��/̕KL��zQ":�$�9�
ޖ��v��� ��tP��Pc���6	 ��>�k��C��2nj���N��T���B�=R,ع��r�*mRyk���q������¡�~�D�pt������c��f�k�Ϙr�/f�ݼ1qiH���6Y�sR��p�Y��R��i�k�[�֦��x)jS���"��A��DD�*�F(&ob\mW��ơ��e�3��"GkM�m�ŸMc���ڎA�Xn�˜�b�T����I��CF$$��9�q=O;�ݘ�I�4q�\����*�7v�Lb����)�N㵅$o ����� �NU�'��D���3Ȇf%
��Z4<��FȣL�n�R�J�mG��O�:��h]�5�y����ۦ�Ӡ�����^j?R9��ۍ@Gɦ�U[N@��Z��W��P\qY����O)~�FnJS��R��P��^�LƄBC�l��GSN��9b�(��=t��DJ$\7ǥ��y�����7���Uva0�vc��Ѻ�W�ō|���@2���Xe�h2�:ǄBbd��%ic�tZWZ��J
���ƛ�~mM)K^<��_N�jζ�_gn?y�,�$�.��dW/^�1�݉ީB��l�;���k�`٪
+���>9����O"�G�0&�5I���Gm�t4���l��"��v4��_����'T8���":�v�C��O�B�R���L6o�c��r�z�ދ��S,��'�}Wҏ'��Q�g��{I���b��t �k|�u�AS��|�_݆��_��6x�g���$����[_�kG[���i��Gw�1��\��J��K�<��*�S������R�N����z�Q��)LE���(T��~�$����G�
K�lN8����=_���|�"���ϬW���9E���2���|4Ԭ�9��ؙ~�OK�*K��F�B�D�("���T�iI#��?U�	�ԛ��w���̽]_��t`�x��^c`I�g��IK)E�L���
qA�)���]��\-�ϕ��g�Z։�\r�PM��Y7�Y�C,B���� 9	:�dϦ����9b��z��D��B2�_ўK�ܥ���D��	9�]��|h`/�}�{����T�={�9-<���%����X̽��1����|�ʅ���y޽ir�.� �цh�=�+�ɲ��^%@E���r���a�zs�wT�����͖f�;����}��c���XFt(F;p�$'`������Q���Nbt��#���Z��ױ�􎀝�\��Tk���}��'U�c	:G0W1��Z��W_ �QCU���S��E��o�#*Tæ��9�ϫv���R�ߛ�?�.����
Xǒ����-N�Q����P����\�	�r�`H�:T�v��R��'%F�iX��⽿����0}�ӗkH�#�$����4��?����͉�CF��;F];�~'��_�Zo)NG��i4]��]�ݿK��T����c� )E@��Dc�o��-�,ؕOIH" �~�;���� �7��v����h�{H?|�������6	�6�6cR$���*6D­H�ѐnŒnoBf+�2���'�&�s:Უ�%/v�}k��?�d�n�AD�O�n��̻	W:,���kY�>��k��Щʕ"�Nt�Mf���t�,�B�����0�_��k����%Xw=�o
��ί�:F�iHhTjIY�j�P�V��D�7�����}��i7��$	��A����Q}:�ɘ�Ǆ~)��dDkv�0a�?VĨ��"c
�;Q����֍��hːq��"q�:�f������m�]��(�븤�F���u��e|zx����Ӑ��;8��7�i~#Ɇ`��A��E���*Ro"���2]l�6�u��q��L�_`Σ��>��*n/,}���(Esp���w篾Ҧ�������)08�ײ������[o�b8�4^Z,�a��lP��	 ��\"�×�ĥM�hZm����,A۰mT�����4�`���E)�q�!Nr��F��0;�ٿ~}0p�8��?M�\\��X�DW��>����W�JN��*CQ��w���&k��u�`�B�L�{�����Z5���k��R��%�ũka�(�@p��A8^�%f���B�G�Q�����9��-i������>!7%j{AG�S1B�b���&��� ���|�<�]&+�7����}EF��GI�G�z�M�����V'dj�Xi�,�C�޵�˿��ތ�;߻��z	B9d:�Z!G�/��]-�\��&�xZ��F�a�H�_m2'81x��
���V�חJmp��5lI��T��\>�R}��9�c���YF���K%o��}��f)sR�u,ϒ�I9��O������ �2�8w�ܺ���~�v�`N�x�̩��^��Ǜ��|��7U��c{���O��4(-M����t����!�Q��,ȓlɞ6��qTe2Sbo65d��xC��Z�˱]K�+x��P�m�"�zF�����B+��[��k��
W�SBc��*�"�9M(M��X,#F�n *%5J� �Z :�}��7���B�UȲ�*X2%β]��b�� h���<����]3�@{˦��G��<U�&�h���p
�9c�{ڔ_����2�l6�%\EQ��3�D�J��G!����S��b��D�/ �7��3~���o��ܒ~��Ö�W�f���Ty�1� �0��B�9��R�ϔn� �sY�r�mB����gՐ ;�㍖�ΎJ����Ű���p��3��oķ��l��שk�m�J����Gof��y�l�a��מ��톖 Ŀ������g����ҷQ��&�����-�귋��+Q�gD@j`������M��<U���S+������Fj[{���G�5�o�%��ۿK�*C�$�)�Y��#V'F��A�Y ���F�%|����47)rq����j�E�\<�@V����Uh�ށ��V��Q��O��V�]��ɵ~��ܤ��3"t	��٠>׹.�qJL������|�}-����a^5��M꡵�����Ӣ��u���� /�t��'߆���Vd�zX�Aa���B����(v��=�tkuق���?�p�;���imWN�y�4(,\j�'���f�f����c�L�ɂ7�
^X�^�4�`�Avp��DF����헁���7�� ���1�>(\�ݹa�r=q���v ~3��w�&��R?K��8m\���V~c���z?��s��='
��M�_�6�;��R=��l���Oq�;�eͿߕҠ��	08��q	aR2��e�f���G�"Z�ӂ=���yfO�����%��)Ac������ʮ�������, ��9�r��I %ՠ&�O�3���Ј��'"�hco��i\�4��G�z�ZN�ݯ'(���;^�1|+�`���%����b!��Fj�SL�;���*����	�����7SNI�G�]�����bLm�IԖ<��S�S��J�ޑ����ם���mf�2�eCGA5}����g�Tk��ױ���ۻL(��*����[t[-좬�R3�:HCE8�[k��"T��2r��u{��ć��)��q�3���B]�s[����x��-���M�o�p�HH�n�o�s��ki]���՝:�x����U�谥z���%�K1o|�u}@��t��/��-�,5�A�Gѧۖ4�C����
tW�N��9�јA fo��C����:rqkNe�g���o^(1���D�cˤ�W�;�.gJ�"c�q�G�h(\n�B�Vo�.Jپ��G�]kCv�B�Ă�H�'!pGJ��d�����z\�QpK��JНᤙ��Jug�:������c�XI�UӰ	�[���e,0��!<45 �Nq���1����,����6� �"�J��V�IX��Q���)�G�ֶzz|��*:�� �aɀ�:���p/�'�I��j�$���t6U"����p"�G=cl3��܏�>\�!�n��w�o&=#ylG�n���Xw�%@(�PX�K�d_S��7ίv2ʿ���%�Hq� ���s�zɿ���9o��_�#%z\%I>W��ZF(����j�=m�K9+bM�F���,�}WhƎ(W��% x�Y��0�)���$�z����_�-��_������c�w��l-�Id���zp�n�'��k `��x�@�ߘ0��(B~i��(�j��WȔkN�4��"`ɢ!B� $i��Ì;@�����!\�|g���b��U��.O��u��+���N�Ԡ���|�u
�y���M4>M�ʆ�d�v�~�G���`h��H��p<�t?�	J�N,Bz=6��W��TqH�`~|��@�FWa�w�OS�D�	��4�4f0i�-+�f�\���RӲ])Q+�k�`�+	��>7��Z��X}�i1���˧�DbS�ʛ���_��W�(N�S�߱���%-�Q�d�ŪW�:�Zhg	������7֟��@�
�Yp~�DЕjP�׬XZ��>�z�f�zW��E`��Ί���y�����::t���p0Ư=DpH���%:��}�s���9Avh���L�a+��ٮ6n7WC� 3%��~E.�t2��\��2�� ׺G�ّA��4�����.�c�g������n!���]3N-�<W�~~&(����p��2(�0�գ~;خ5Y*�j7�ok0�6�����$�XJ� 2�y�Ibj�n�H�r�N	aO!���QV���=�Hr�t^�Qu�:�M���ӧ$�HZ��{N�]n�x	��"^xC�|��+��O�z]\}�	����?��OS`d�x:?�����d7Ͳ�,��]97E��n���C��C��:wcF9�u�hi��z؋*YK:hi1f%��ز�-��R��h*{iW"A{n��豚����xo���sRSק���5���rI��H�
�ƕ�[�zu]�W�c�\�J�/B��%�q��[�B�̗��z�X,,͛�*����ii�8����Ģ^��j�q��B.�`�1��!�۴%RT��Ê��2 ��~��KC�#��\��I<����Y���E?y��[	uX�T�.�?�3�Q����Ǆ����q9I%��5�f^�όS���M��DQ�]_T�iS��P�̷��j���WsM�5
��4�u��8󇘽�]����*iC�.��=��k.ب���Iy���:�ߠ��ݡQ�y���c���%
O5b�\�׀��/�jۍ�%�y�ߩ�a��i���S�]���Q�<@b�LC���x��I9��|�:�a~ʰ��;u�s����R`]^���PSJ�x@�������m��s�O$
+8��A��4�`��@���ʙ��ظK�s�5�Rn$�n����h~�kdУ����{��~�!3%�2!�o&��FV_ns Z������!���c����'M���� �Oh�~n,�a;_g�Z��r��Gp��oA��%#��� �~��Z����&K�;��֮쵑 S��]�y�uc��i�ӈ|�;m����j*T�z�U�2���<-H����im	1�:�g�"1Yr)Ӏ��1�-2�_)� �-E�U!O7zY.^w�/)K<����Y�]ٌ.M�F.� v��u�ѓ�[7�]�3��kɓ��u�+
c���/kq6��
����Z��;-%@�.��	Q�ֹ۠W_�!Zd�l?F;i�ƹy�U���Nb���2�_+7��}g�fp�����+p���){�f��:�Z���eX�]��|!7�(�����+�+lC�&5�y�Y0|G�X)v���v �]N��៱�(����~ƃ�Qf�A���2��)A��,��Ja��^��7i��	�)-�?9`v��'�7띾���RŊ���c�����Ԑ��}@������pj�����{x1�Y0�D1�y��):ç��d��q_Dfh�d+�^Yh�/g��A�u!2�r�M��y�V#���>�0��m����ѽ����-&�u���*��x��I�jB(Xܚ����n;dQp��sH�&����#(U��v\�4	���m���1~0��v��hw��XhN��ş��"/�_r��u/�Ē�3��b��EgM�a��dM�2,���i��X�G^B���ޝ0!Ԏ�Gz~�z�'�M�Q�D�}2�J�#FUf�80��?�xa$�~�~V).@ ��dJ����<ٶ�L�������h�{]������s��R7��쭃��pU>�ĭ�>b��1pT#^Z�EYZ9�O��y��>�{r��<s)A�q�%/M�X?B��!��3>�&�Ls���h�?�H�Cؽ���%��e_��-��!����A�7� 3�-�]Hoo���BkQ�1���S_=�(�5���g��K�2�K��ՂQ�x\��.f>��+m����wG,�/���Ŕ7_V��31�3�Ũ�*��W�5l�{�N����b����i���H%���j�e%>zز+|�f"��w��r)T��p��'2%h�74(f�_��n����J�ѕٞ<{��"��I�f���E.��fp���g������t�^J����6�a+{t|�8h_[��S.}�����7EKV�p��絯N!,Ӻ�wñ�ݕ�U�˪��3�����}��O�^��@�*L?�~�j7�����(�:���%�Y�L|vf�F.����Q�eƪ?�=+����TP�`S�\=�P���J|'��mN� ��[A.A�X�(����;��[<X������x�\���*Au��"� 4�~�16	yE�#'��:�7#�O�C��W?x����<+��f;�����S�jif�/�
��S�z	׸8ÿ�֏d�c"hɞ�ڢ��+
.��.~��NR7�z���Z�}8%bɸ����u�s��(��Ά����ej��t��/ ��ҫ��2^�(�b��^�q-�tc�P�!:O��r�@�zG��ؙ��3�~䃒zp��:&)@�[��:�LS����{����TȇEe,�Ą�w��)}������/��͟~���������}�:S��J}���$*��F�J��?d�T�]�-LKq���S�]
�P�ݡ8���-�Z�]����Z܃��~���ެ�E��9{�����<	���`� u]v5Jh���m���"Y�Y�ra��(:��d�$Ƚ	�5�7�D��M/6�x���2@���zcj���K����G)�/Ǎ�*y��#.rȲ~��S�;ώ�9��ʼ���K��@1.sD���3-(��o��`c�DА{�?d��ۯ��	"��6��-�"
;8��=Q}�^'$&�HV)���eF]d�>��������Zm�*��B��~��F�Y�9a{~��Z�������P y��8���(��MPg�D�NC>j�80�.�@cQ�^���'����4�Z,�
*�kѥ�օ���9>_�\������m*����j ��m�c��#Ǐ4w��?����N˴4q��o�\�E�Wll�jG?	7�w�"Y�w��Qَ�I�[�f\f�Ϟi�=��g�u㐈���{���f65�~�	;<�V���w��������d[&Z�ߐƔQU��4#�(-��C���4�$��j��B�Y�8���4�� s�����+o��~��W:?t�������i>�&�c�/����e?Wϴ��~=�ǝ��NbS�G����g,�~1�v���H�ڡ� �vMG`�[)����q�+��7�����Nk:��j0�5����e�G\��Z�h,ߒt��]�(F��"�y��q��V��L' �!��d�.�����3K��� 3� k�%ȣ����ꉛ<��Ȓ�⊝��>�IRO�r�<g#c�-?��P4���Y���M�9������]��l\�Ÿ,��V�x�zHL�E^�~+����B,b#䌃&�1��Y�b�E�w��y������rLxU�%k�O��*�뒄�'�MfJ��h��Or|����Y��m	^��Y����Lu8��)q3}\ߦ[V���Þ�<����a�W�5�f�sVZ�$��ݹ�CZ��w(���W1������x� ��7AT�rlT����0�q��D�P"|u�~
P�ʻ@�6�q��o��J�H��p���k�C�v���5 ���s⢤@��)\��u-���O��H�[��SϠ�Zr�!u���xH��AV	^G����!j�ԃ(!C��l����w���:��o�y s�u}���\Hһ� Qi����sѵ��y�3���)^�g�o�/�B��4�W]�����$@N[�DsW�"�
CZ��r� $)��L�<R܊���~fƴ��AK��������:��[�}��`~�4����/s��-�����40y���W������2|���Uꬌ�G�:H]$G9�Y	���W(6����59�������G����j r��a�9&�_��W�-p���-	 ���X��[����7�/QZ�����%}F�����UW���Ţ�@uڤ��v�I�^q����V-�Br����F^`l8?����(e^4��d꙼���[�h�ɡ\�����y��]"|W+����c]�8�O[J��K_�梿��߬�?�BS����mty�AR���!�d���p*���0��-I�o��uJ!�0g��n�?-
Oz 9V}zy�CD`'��ܹ�@D/�����&�u������Q�]
Z�8��#%���ܬC�VI
$n�`U�X6�M���Qx��R�ʗL�d�̻��+=�񰳤?5��K=%����IR�Q
� *W�U�>%Ѣ!��%w�)�-З2O����]00ϕ�����P8��F?�EDEX��\�>S�+���wq�^���{�pё���٠��'�S���IĞJ��ZȜ_ix������b`���Jv>:R����P�axUJ��Gc��H�4�hiE/W�������C�[�25=A9G�^BF��/~GC���c��l[����r�|`H|y�c��h���T�ʹK�:8cM�;���5)��q%�9���3b��y��y����O�2�<�6�������=�{i���f�Thm!�9ou#�Kv�E;XQ�K�aEw�nS�K��Bv7��[��6o��.{	]L���<�|Ѳ�[��)D����뷣�	��Mn���n%���*���~%gQ��},'rƶ4S.���Y�͞�[񳙗hHV+Dh�ЫΡ���x'��(��.�'��Or��a@�[�NRiI�aJ��tȂʓ����;A�<��^+�1��A�[� ���H��#D�|��%�/Cl���.�� 
�n�5���{+!�����&mA�~����
��M���a��A�o-<۹J-�
�YҖ�� ��zg%�TAp�����s'x�R<h�5l��N�3H�L���Td�R�4���˛�J��o���`��V�;E�;^�b�������ؑ���-�/"�ɱ<[��v����I�8� 1�[�&a���xS���M�ŉ��OG��TiE?!1���x���0���E�j���nR�RC35J��� �Ț�-d��;�>z���~S��c�}r�iu>a?����vo�&j��~��AÖ<W��s�_4�S��6�q���n�L��H�^V�jq�#?ycW���MƵ6T"�:,N<�^~]�e���z�J�����A[ ��لqozt�W{�_@\ ��i�^Юn��N���dwoA�����8K����&d5�Jz�oLk��F�HS�zr4����4�m��4)��Z�}r��'ѱ����_'T�^�YO�ep6��r��{��Q����|�H�NE�P��q,5]|�娂��I��8<��x�X��Q�%c=���� ���h�le=�n�S���iEp�y��p�?G�yZ���[63�vy��M;�`�z��V�d�S$Ym^�W�.����AZb�;�h�k��Ԡ��M��O���L�n	��#\ӭg�t��$�����97��Pxę"�o��v�+?� Ь*1���tYZ^���
�]�����;u�Ǯ��`aAЇ��kz��.�+2���ӄ��޻
�G�9͠��8���7��|�F���QO�0�t=��ס4��.���x����]W
�%1<��F���=��ϋ�y���5�7������+ZS=���h�X�F�<<�%��f���[w-������K�Q(���e�NK���h�u�O��G�Ztg�-R�,R�Ń���ɴ�ʜ��Jw���bsީ*цN0��/K�kN}�
��l>�Sgm�т.u�`��5�W�BM7���Փ�|n�,YZ�&��8:r�qpbIX��V��F���6��O�z;+}"��ž���	ͅ���LћV��@wu:�$�4���[��}�f�D�w��ꆖ���zF'v=7� ��e^��)A�uX�v]��Y9�ڼ�� -�t������sK竬m�aq5놪V� 6� �2b��RaI:��_o_�jW.��1�A���U�Q8�*�P��Gw���[�����w��<����)ƉWJ0k�ׯ���{IB�g� ��hgQDY�13�A����uʛ�X�e�O���W�����8�F��c(���h/g5��e����3e�H@�Tcҧ���ע�����`�JV"V��E���9���>X�Y�4S}�A�0�_h���1�)��t�[:�o�K�)�bp��&2�g|n\�VW��b���B'�KX[{�Y?t��`��zǵm���|<��Ӓ5�r/#��6Я�e�!xÕ���x�	cFef�?_�y�u��?��O�l�#�-e��� s�Џ�v��=ז�Q����T���]���H]�,�Ǯ~?���>d��
J��\�o~��hp'L
W�
��[ ��v�ť�"S��\ -�9��� �N�^ςRn��3Y��`�02�`ba���,�1��V�����к�7m%ɹ�Ի�w߱��xH�����S����"_!�)�z%�5�#���Y��l�=�3�nz�jL� D�}\X�ˌ{Y�D�+����h��8Fy��������'��լ�g4Xs�������c2�����b����z�V��@�T�?�LW�´���v/y<���G�y�=\����\�,VC���J*\���[r碫�O��"���^B��t��D"��9Ok���ɟ%V�{�*?|}�P��;���;v'���
��T��_p0GvI�z�8N]d4����뎶�J=��66j<���:.�]�]�5�8#F"M.>� *�,L�7�;FԸ��=�&$���&a�9:�;��h&��%]��B����$$����jv\��F�J'��"Ύ�����%��k�uo�)���c�g9��p׀�S�z8e�Q4l�z��>�|���pl���B�� g��i�K�Z�%�у���y�zj0����;��͇�F��u|� -�΢m�c�ݬc�Aү��5-!������Y��lӚ}��{�aE�BC��ۯ�`Z�g�ou�+�=g9v��<V�l�Eg\�ܟ������g�q��X%=P.���_����o�`�+��Ɩ�%�ሥ��F6������V[��l��nI.T��2R��U�^�eObZ���N�|�5��e���i�m��W�g�W0�*�¥x���֎o�����NY���ك/�`@>c�uc��-x|Z�F{TX��VeS�.p.���R��}0��H�L�	���n ǌ�x`�ap����%�=x]�ٕ L�x:}�+a��4m5ˢ�ÓV�=��P���
�bS�]
X�DnU�0���9�r�L����Fol<�d�[<J!��}�I��0�����g��i�{}����ϵ� �4s ��~#x�|B��v�}�����8��#�k��	�%�Fy�j�-R��T��&�KZ�t��0�����P"��kTi0ź�Ǉ8��R1�� @$�[�n8����_�C��A5g��9d�X�z�E�P�!!�{3&&p;G���.q��̑��,��q���r��R�8{b��!DȍH�i���n���#�D��L#������k)�ȵ�����#Yt�6߈�<tH4�K�ƥY��cv����vy27���\�B�&G�N$���i�/-���u��{��U�~]���U�YYl[�t��Z��|n��2u��n.�p=�6u�tR��b�ݐ��~9���B�XB���l˕
��c�4�8~;gT�S�ծ��V﷐����7�녵��F?�Bc�2=N�s��&kv6(�Nɴ���>q}����Jf�:~R�D��IX*�����/��j������f"�J8p2�\q�l��)��D��;HÌ��@��9�f�0�;`֨��o�ʁ�~"c]|��\[9��U�B��v�GǪw��?
���3�or�!L}��X"᷺�
��ȑ�ᑽ�x\��N.����fU�(;�u�M�5��ɱ"O� ��� �nHW�5d		�M�)ROC��H�k=�N]l� *���!�f�+��P>Z����RyGj۳ż��GL)'���=�{т?�ڜf�{霛y#۟�Ei�m�Y��-x���	��K���l���I;���F�;6�����������Sw[���E�X+��I_�{
״����e�:
_gAa�ʴ����^�ŅC
��;�7������� �?@�r!�]?}Ü���Z��{�sӖYJ$����R����l%���6�T�o��������#��n2���C��X�U���w�A�@�k`ےі�3�����8�:[�~��5#���j1�@�y2����f��<:���:!���K��=�L��t�$��_�;���S��\�w
��mh�h'���k@K�
y猲k{��-R�0�L#���
�RT��إ����Zx1���W���0�s��{��`h��G�V���� �����K#F����}�d"���Ƿ��+�#5�jp�FO��ij�D?#�I�TZjDmӏ雛љ7.OsR�2��36ZN;���������4|���Ѓ�T	e��`a�OX%�%{!��H���ݘ�VP 4�C4*b
pvv��!�6��HJ�k�ކ۷�a������.n��<�LMp b"���xI�4jn5|	g�)����W;û�� ��nf���Z�JZ=��� ��Ot��C	#�Y +� ˨:WA�\ �)1��ZЊL�;�[P��/"���,ū묽��Yo�F2�?��6���ـlސ��t��M�:�'���y�'Q����z�X�]׶���� ��*�����S�KN� 7�'u�{H�֪<��*sXf!mw�M��{�������[]o���ĩ�d�5o#�!��4W7,�s=~c����a��$�2[�]�~�Gn$Y�wi[o��T<�ʵ2'��h��ZW����\���.�XW��+RG�Sʾj��Y��'`����e
MS	���Q�'�i��S�Ê�X�L#�yg��(n,O�V��(X�X��F�M����JRd[�E�i�V�i<�>�8�Cz^g���ml��ث�jm�Omtp���
=�=��h��C�m�鐔�C?�]`�> $e� ��*��x��Ar�W�j*�."=�k��Gg�#U��
a��Rn������YH��M��2�m�|����E�Ғ�7�V�ңL�@�}���O� ��q+�ΣUݯ�L¦��{[�}��U�n���}�Z�s�l�t�x�yb"{.쬵�Sʋ�]��I���0
��#�����̡�q�<!F5��8����AH�֞�ۤ,ިiX��Qy�v�m6��̀:#�l��L����$��q�9��
�ء��EZQx�<c�L�g��=D����|�l�3�R��H&,�vP��U�#ױxU��݅�9�%� �f5P��p�B�\b�>�@�cɩ�X;<��w*b�����,��P�_�D�hU^4�I�y��F۱ǣ�='�%��Z�m��K������ÝЊ�C�ԟK�Y�<����艴 ��Ⱦs��D�W�d	�#����Ǿ
ܫ)Xs=�8����J��9*8��M�D��DB�*Q��f���?�˜A�eg~�4~�Rӯ� ��b��������]����o�g ���P����L�kX)�Bs��ҖM�@�o�=�h*�x��Bce�ύ�j�-ݿ���e��LU���ڢ;��������v@�cLܜ��v�S=�������f3����:m�{ߨ^ƣ�0\3�dZ��<\t�v���p/�"��P&ɘHH�s$Ij��5��9Ue(C��kM ��paVA�g�)�����w�و�+R>Mfl���NHO����v	I�n�J���+z9������~�����3�%��,�O֚��ñ���g��L�>��]5;�`җoJ����h��ҩ�Vk��D�L�P7�{ϋ�i�n���t�P��ί��?�+�������h߳'G�V)}���?���'-JW���yDR�7�ɦU��˰dbd�����#�8?�-�}.3�y3�m��d�s!�~�6!�{ϼ<*���H�r폆{���P�~��3����"����H��yՎ=}Լ� O���YB�����ϸ�&�g�(\�����6?O&�apMM�*|�1_.>(h4~��0@2r��l��h� ���ǹ��^M��`�a�ڜUv����{]H��(ה"�:w̲b��~�уmD��&�]�/���_�c��{?����:p�嫻`��~�t��SCv�"Ay��n�CA�q	c��K�ʍ�w�������B-�sI�qij��!�AZY��ݼj��܍<���XL�}4�i��G�\�F*ٚ�r��)�Еv�HW��t�(Yiw7�]����V�l^ʼ�kh����sN.
��d�u;��:����a�_M��mH���w��I)�����Yx�#��!��x!��������Oc֣{���E<��F/��^f��т��nU<iKyZF�w,�.ey_D��<�<u�0��o���b���s��Q�;���j^D�v��/�78)`�� ��h�ŏ�܍5��}4mq�TFg����1lfI52��]���J<�]O�h�X�B=�5ʪEx���<c��Y��;�6O&<����-��d��P���[c��:Yͽ�b$�z ��'�&��z�
q�����֭/	�78x�p��5*H8;4yX!���H�|X�}�cg��&g=
T7�1;�)>ݰT�\�I1��hZ Hh:ހ��a�m�l�8K#�p�x��:���C�Uy�J�� ��`���O�ΣfF�E7��NᛦW�
�~v7Q��G�LM��B��}{���U���2z�u� ?`��Og���gp��M��ώ��Eg*u0����a��(���\�u�	���	x#v�;g.:&�����a�03"���BX�����S$�F��k������-�cF�N�C��5Doy=?}������RRi��Y�Z�u� 	B��� םa@�Ml�n�LxJ�1m9�^TQp<ޢ+��jcm���`1A=��?�y�VQ��|�3��|^`��}�Td���:]&0���W�
�h C��ib�9F��X�7�¿�_(�F�=۰�[R��L;�ڼ�nC�wo�#��#��ݴ6��f���QN��M��zr��V�:��)��!�ÍD-������$�6�/�$�K<�l���:��[,���nz�~��i��Er�R�b�z��I�sFٮ�54��2���8�#�[��K	��M��%��=�b|�z�-�J�1Q��F��=U[v�8��9�zY�����t��V`/�^�W��7��ӏ&����k7i��>�T�?�I3k�^�p*���+(�$=g��9Y���c=��~�[z�U��x�d�I2��B�~��y��匓M�GFA`d.��t��:�
�s��k���v��gA�Iw��M����z��w�ܴ������'>W���5�kA�NĲ�{؈�v��c����]Gm�BE���.	�B��,Q}��ܽT>*r�BǨ!��7��u��{���'s�A<Gn�״�R��D���_L�G��y�;	eD��)��uB+1
����CcR����O�PK�7L�k��Db��� ���  H �	��ms�i+B�Sܺ�G4�Z��^Kh��D{����G�Ʋ�ݙ�ŭ3:���Y�'��Ì�`zA �>rsR,�[��������U�C�͡��i���M⟓�Ք4��X�f┻��?l�R`4�C�l12��"4�g�� �H�Yz|��k��zۮV���U�B�/�-��jPa�Ң��:�4�@��?�3C1�}�ԛlnT�L���$�|�c�ѱ��Ħ��(��
ۭVa�ed>K�O�}|���]N.n�π���^�u��m'_�@æv$�~6K�W�|؄�k���=zm�0��e�5�I)z��>]�B<u�5>g%��k.O׫��<��h\�Vn[$�\��ӣ3zO��O9�\H^n<0�����
Z�	Z�d�����o��-�py���7'q����'�O$K�RS�對�Z�0zP����Ąx͗�����5v����t���f}9F��p�t�
�)d�s���t��tqW:�g��pl����B����e|LMH��N9�1���Xd�B�l���x�Y��1G\�� �꿚��R��&���G\~}���P�\�3�@%���l�����p0�t���hZǗ�����G8b��C<�0>0�'�k��Y��'�CU�Qa��O>��|����o���M=l:^���g|M�!*��6�9��OI�%������
�?cqȐ(������o���d]o<�h��V���6=�X�1�>6^��&�{������i�*	��T�`]������������}̞���eR-�@�Y&C�{v�+�_�\#��P�Xji��m��W�V+s�6r^sW.:�kN�<��z6h�o��D�}�X�W�,�ƥfz�]�;�t)��rI�!��DI�}y�m���H(�W�{85���M�kw����=[�������w�t�dI�517��*T�!��&E��O
�Oi�d�d��������D1_ƙ���w�~"�@�y<_�w�	lw��C�yko��ޑ����o3��>��G�G=�Q�q������i�V-|�Y��Y�(ՠ�QE�8�L��f��j��zy�5������'|�)����Mv�~�C�x˒#6Z���A(�ۿ���nYs:Ʒ?�<��=�������?�::�@��Q����D�r(ֆ3b	�H�m����-i��yտ��z��ҳ�[C�f˚�3h�I� ���)��@b\P�1&�$�V��{�v���S��g/·���'��@�C/����������n&�Z�Ów.=��>g��@�R��E]��n�(#N�=' �𦇪-�3�U���ߗ��E��@w|���2���y
��|�qwF�hݨN�����OR۹L��o?J3�h���r����}�j�z��QW�}bF20������/��jI}m;�s ���z��8�����񷕞r�|�#3�0�X���@A��`I�kQL�-�����q��FPqZ~"JUGm��R���x��G��������T�=U��o�E�~�]{%�c0�C2K�7�C��=���;r����[��p��_Р�F�ƒ�o���6�-�N߼������N	�%����5���bBˤ-��.�m��_�RM��1����r[ۆ-���RJ�U�*f;�_,��7ͼr��� �i�nON��t;�Ϙ��f+��3���|�_�2����D��D��
K�� Ōg�Mѩ/�ZOs��|+����cy[H��|�����'+g�:{��!�{���w��̧�O�ZV�8%o�q�B8� �D?����l�(�K"œ���(d� �s��4zT��v�b��CPm��9.�:��ox0��u�F�+��/��׺�<�e��g�'��7�OE�	�u�>�.��\Ԝ�<[�c�ƺ�P���0N����7�2�e6{�m�����@�� ���2��t�+�\S6���E�����g�C�9�\���!ӭ��.R�Q�Ё�{�\��C���$��y��b$���>�y
C% �̩��8�g/{��+޽��m�a¯j��{�O����2D�21�p��|R�j�C������V�\
�ot�98��e �]�puC��#s�`���
*�l����r>D��͆ �f��P�\��&�k��&��]zb(�wzXp����Aْ�,���$#�*Z��B����7]t�Ǹj>Z��[�sJa���-��9Gp���uWC9�+��R¯^
5NJ@��7o�A	�n`�e����֣y�N�<��=�����菓�8#GB;��]k��G��̟�9���87R����'��Cn�����Yʀ@�X~.b����q_�}Jk���QKs!gG���2�b���D�����	���.�h�xo��s���]�u�@k�h��t�B��ѩP���WX;Q��Ȓ)I���9#yɴ�mka�us�d�ϧ���`�2-�K�'��N����T<ש����H��M�:�?&�z��|��ם�4�S��d~���d��L�I�]���V�U�9?�Cuk�Qk���b�c�%��o6W�J�o�3yC�^��Wn��^�̘�Cfq����5�}&ts�S�}��Q��9~�|��Єt�@G�ĥ��5O���,~	CUs1[9�������C�/��?���GݍV�������GK*`5]�#=_˺M���kY�\����tN���	�m
�\�x,V(����~�}#j�t�q�@C[nM"NoG���֔&q(�q�ܹ
����"�_����۸%��wfvT�[���űl�/.>���Y �u�m�����뇃�G���p7�Oe����AG�z�w�s�j�w�5?�y:� �;E]���Q����S������E�W������}]#G�ͦc%���rw�h�����a�3�S��E�[,%mݟ��,|�fE�k�h	۵;	�z���S/�W���1���s���Q)�|,5y� �E������я<[j�p˯��oOܶ���q���EDAX7N�ن�]�tuR�qi%\R8�np{W�b�Z�"�oYA�D��,J���+��;�)�F>+�&��_��s�H�w��.�N�A�}��mF���������[�UX��D���w\g�q����L���ܜ���d␳�Z��Ā	c�qϟ���o�U}������x9w���dl�h�U��z096����/+b��������4�~�)�T9:�eOSe�Pz��v:��m*@`�����(���� /*�7�I�[)��D��C"��l���j�^�����S뭐V��3���<X�xO�I�I ���k�E�֡S{���6��;�*8�?PG�>>-°��1O8�s�Ō�lG�w�XJ�.���$�I����m`US�E��M��i�@u�o]j̰>-�'����&mMu�?�VF*�գ���黺�o�s��Z����,G��2k��B�t�t����V���؝:y;���:�nd��P	%��Q������V��~;&� ���FI�����!�` �Be�[Ԕ�h�U��q��6PeF��!L���A��S7gf�H��x���?�j܈���]����_�/#wWz�t=�5]82��>n��?���L7L�ֱT�(O�]1�
/�ᦳ	��x��Y�!yV�Y/
p1�[fs����>}���s\���g���	���p/�_���*��F�AI��D��d5DְJR����:�8�Mw���/����*���e8��4��]:�1T�(�ʿ ��1�Qȡgp+F[�"��,��b� �+(�8����#ݶ�_-�e�'�j��qRE2|k��?��F���<*�j�M7�+�����z/�����NO=
1�?Y��qf�H�2��i�lRca?')�t76�\�ls���Oυ��Ѯ��4���͏)T�..z�H����W��".k����|�RSdr+ǘ���sQ�$G�B}Xtr8[#+���!Q1վc�bbk��ʫ���ӅsNg��������.�2���w�*�K�(�*�W���_��d�RF��by̵S���VX�Ge~�<|�]�xe��E2�C{�'s2�#��@���S���ja���ԑÉ��J;�?���w��g'χ�Y�ֲ���g�c�f�0Q�3�������E�V���
,q	�% ��H\;MK�:����N�|�n��D۱��;̡A[\pbU��c�]	��z����R���ޓײ�"&��K�=��g���I�4.F���$D'�</m8�k�t�i��9?��p���P6��6���%����D���f����z��֌�Q��]"Έ�ݵ/���&[���ߚF�nG5���sd�ь��z`���՜0m�E�֍?ht(Tj|�b�6�d�y������2���G݊����d��L2���?1:�#�S�k�df��m2ۛ,�#C��>�f���[i�fO�m���@�>����>���B�{�b����U}߅�E>@[.�B�Ib3��:q��'��a�fb~xjV�Z��\�T<�ΐ��a��Zl?�2O�����'�-��r��{2���>T��>|�?�¹�q6}���|. Q��P.Hn&��!�輵��f/ަ&�2P�����k��ri�ގW�D���0s+sbSr�ϔLG�O�J�8A�Q2K ~gɡr�Vۼ�	��t)�����A�j$~��#w E���{�aX;�QZ�Aڀj"��?I����Q
�Ԍ�^�hi�;��Q?M���ͪ�^iڎ�6꾝�ѤΪ4r���ic�HY�:����������x&��\�ˠ��{��z.'d��묛�f��lZ6rQ���^:�(0�O�H�	Ӻ񷽦A�$�Ug�	���KWm��`vx���z�	7x�N�}besƘ���:��M�2T�0����k�7SB���e��]$�ƶG�Ƞ2M�dR7p۟�	�G�u|TK��e�ں]�L�2�
HNSp�ۈ���+���]�U���4�tm\�DO�E�;{��@3�B<��U[7�G١�E��nTj�Tk:[g�v0Q10�jO��t΁ɼ�V82�V��O�9rk��5/PN�6�/y�N�'�*1՚�������r��Q��ɡ��e���|�֫`y���uʵ�@�T,���<�@Nt�9,��K�"{1Lrhv����h6K�.�0�Mrdq�)�p$�M2G���f�>e�Rk��/D6���Mʱ�ǟ��:�%���B���I�4�)��gQ�Ć�B'���ozKН?
P�(�_�6��Sg�L�g)=�e<�����9u�ΰSK������<������v�z2N��"�>�~���`+��5�7�ă��">J��a�#KȈ�SN�`�����1G�8���"�ƫ�Ġ�x��J���ѷ���D:�K�n7��T?먛͏r9_���b w�w5��Y��Z	�*�/�=�7._�F}��Q��]#��@��+B�d���T�������Q(�oC������K�/�柕n��Ҟ�׹����r�eS�?E�{��VH�JY�>�k��O��#��O!�ՙ�Q'���W�������tc	-�� }nz�2�9Z�����Y�Q�k��\��A���c�n8֡*������ק\��mv�r����R�X����y�_۶��Xt3��e�5i��>[B�8g���=��$���:&�s�y������>Rf�q>n׺���v4鹜�qry�=?w��n3����C���_A��?���? Q�ɪ�6a�;��j`�Ϲ���i���~3m�wb %��:�L�L���
�}��A��1�����K�C`9�O��o�@7�����=
o7��a� _P)��\���r xܿ Q"�$��>n��Sm�I��U_rf�8���{^�IJ�G繜��9�C�t-�$҅��b����W��A)5����(�!Q��?T�2��^<���#�D���=Sʻ9��m
U������K��f�S�dO̎^x>bKA&��X��O��b��`D�@G�M����{�FɌ�L? ���7,�a��6Cg�A���(Ec֍w',k�՟�,;��Wl����[tW+ �O���3љ�w���U��F���)]�]�8<��&��/���@e7�I�����Z�Zk{��v6�E���q��|�h�h����ģ��U2 �MI�:XE'�+����_�)
��aASi1�;�K+K�sy��g0�L��6ѫ�����3;h,�j>��D��<E�{�UD����q�4&�� ��l�}<���#�&q/��>ř���P
�ܩ�'Ğ�I�+6@�W[b|�FR������Z�>h��q�g�񼯇�ߝ�����b��Ɯ�^uݔ�/����g�Yb�%E^���:�R�-J��
X���Rn}��`���oC��9��ʧlE���d��K�O}��6Q�r\�9�7�+��P��포�B�ܯ���N�X��	����l�G���P(����l�J�����!�l9���H���*�\>{k�q��H��}AK��"��r+��?�Ky1������W���+XAbDc�f�#���/��J�[�bu��y�G1i�J)���
�yε7�wВL��2�����֤H���Z\Pbm�ë��-�5n��+��U)��-��6'�㐸T�Z�M�]Ƙ�_+��n|�a_��V%���6W�x!�n�*B��J��g,l��Ѡ)�k}�wCM�Cdq���Й�1�w�\|���$E��џ>9��/:8r#7P�ę�{v��f+'.���1H<��'���2g#֖�R���.��J�M�yf��>�DaASN�k�`80����L4����c���b��R�(-o�p_� ~ۙ�hL�+�g��S`������E߾�c���Im�vL(�`��{���81�N4��0"�lJp]�.!���l[��T:mE��M0`�5�\�&��mY�f��������ʡ�7�L�ۣH�:9#6��?�X"p����r������DG�cR��Vdis$��]�&*B��N�ɨ����h��K��ą�i��K��ˏ�5K��!d�e��;���=�p	Y׬UZ:�����Z �Ҧx�ꭅ8c��:#V� ��eA�y����W�k��A�;���F��'@ܦW�Jؗ�u��O&B�:��t00R?KA��6�j������!x�u���d�	�Έ�%c��d���Ʉa�~�4gjB>$J^+�x�'?H����%�C��A�ߕ��Lx���W=�_Ģ������!��\�G)"���s�T�s�����2,���PH�5$��)��4e�?����R�.W�q�j૗�~�]q�?�;B�|_��῜�}h���R�3b�̺A�|�e�+�4@�Z-��bD]b�I�������p��E�a�%�v���QM_�@�]�7���1�B����QN/�����D�.EZ��X�X^�!8\,x���|��S�<� h�G��Y+j�����|��������3�� �
�Ɗco�(f�����`K������"����l�M	�2���)��'�=�&��Jԓ#bC^*&oO �>�W��X��\��U�k?��Ά��Lř�������K]&�9R-С�&!��_���	��#�L��s��b�����lCM���%��Fd%�v,���nT+*��4{	���W#N0�>�'ę�PQzK��|gTS�ҿ�r<�*�(��4!��t� ]��@h���j����J(J=�H�R��{'t�#�����?�k�_�e��v���<�L��<��|M֡�XV�����<A��6��|�D�U���i��iH��[����-�3H����ne\��/E\�e$����?��_��}|U��v6l�VH`�5�ז1�Ӧ�ݒ�j��6�QB|�� � L.�,S#��Q�v`w!�ZI��5��U4=�&���c��J�~$k���Ti���@K���~��O�{e��sR�-��(���-�$Gzk������^�iO�;�)��DR\i]��`f���,EB��'��g�=�Uh�����V��SQ9����y�X��@,�iD: �$p�����*0E�����j�(��h0oq�2Ъ�9�����qcrw6��9�L7�&�9\���]�������(# 侽Z׫FI��9�����7?�z֏fx�֝ �0��y �����)v-np�?�yGJ�i̒�=���`���!1a7X�F�í��*���>v�'$Bs�� �����$F���-/z�THl+���ϭ�T�N�@��&�\b�-����_6G�D���=>���)�5u�_9�#>d���0A���(�/�^���j���y[�%pH��y�Y�GR� B�{�,?V��3�C��X׼�P�r c�q8ޝ������(kJ����i��VHI������hw�9�Mb�>��l�jN�Cg[�`���$��\�J�3[����D)�!�ͳ��u�����fq���1+q����8�EN$>��<�ڞ� �u��{L�_=�-G��G�F�J��iih ��7��w�
ĥ��6K���~��Y-���ě�3,1|�w��$��*qI��;�&[��j(��H�y�9S$i�S��� w7P�Ա2��&'�����}�ei�q���w�W��{Vlڃ��Hb�z��]<r�D��H����; z]�����v�>L�%:f�6�`�kޕd=1l3U�����F���9P��Ʌ��(>G�ˉ�_��+6�"*�d.S�{Z�c?��_!�,x�绶��=�hH�bJ�I��/b�����5brʯ_��R�_AN*��Ai9ֹ���x���V�ON�;������~
��l�_��=�{�׊�J/c̸�[���Q�@Y���v�(m�ܴ�RI&<|3u�2�;c?Ѝ�Ş<��~>lU����Á٣"^�Ie�9�
lC������P�#L���*�s���O�^�-}�D��H�D��S�fyhM��v#�͙��e[���h6�j�N@(�e?�?���3�;���wF1�40_\sV�joe���׉ ���}��9�{���Y�~��I^�2���/��|+�����j����ҙ��w^�1ryO���b�]Ӵb~{�|�yƺ��&�l͹����.�q����6�`<�A,����B7�$�4�1DV�H�S[�)��(}M����f_.sq���Щ�K�6���;*�]ju�'�������0&ѓ6�g��?��ҵ֍I��k���b���j��9H�0��?�}*
#�Easn&��E�'k�m��vJ�/��yu���R-L|��%JK��h�'�3L�j��:����'�P�ӧ)�p��i��ީ�%o}2�t�|>e���:h�8u�e�O��בݩ�W%~��_ݵ}gl�9�@���,V�wVP�ӌ��B���Qߟ�sA�	�3V
�}T؋L�}��H���V�5g��5i��Իb��\D�<!�ǌ�.����Q��n�k�>�_>�u+ɢ���&z�����׾4�Go�p�S��+`��j{v�FoEx�
J���a���1��ԊL���!hk���m��޼���g�e��Q����齻���%d��^�	zb��fb���_�G�s>p
�$����ck��ɬm��ú
WV��
�&G��"2O�T1~JOfW5M��ΊSc*@O��7����bؓl�12<Ŏ�0����!O%|�Q3���7ν]N~�4r�CԄ
�(���<�
��!ZI�7����E�s
�Д�ɮ/�5Cc����<DAN�:��U$���B^��	�����9ܚ�����[�1!]�A5˝�-�Ԫ���!���<)�j��2�K9�q][��ػ�+�K>s��ïK�C!G��.��db�@��#+A<֨�[������s8l�,7|��p�͛�:���񮢼��Rc;�Q g-VO���	g��ᚾl@�ȎSg�N���qP����`�-�U2(��Bxn���^�ZB���w=�I�t����8(��F�Galu�Y��\�҅ ��bP�E.��3���?.[Ⱦ��h�n��E(��6�{�U3��V���:F���U���L^���;�����>"�xD$�݈�Z�gD����n�l�p[:J����у�^���*E徕�//:s�;HK��&���ļ���yy������y�m�/��Χ�PC[Wb�猯u������H�#�g�T�y�E�Y�ce��<>W��:��5�Y�қ�"_	�����g����n����8�n�nK󕼛��*x��Ss۝ �~n!Bz�מ�6��-f[����[^�s�� eM��MǼ:��r=��@��F��s�~���j2廬�M�7��E�|&x]]'V^�����`v�>�B���I���V)�����2���I6f�l4=g��7*4a�� �>*~⺼�H�pIM6�-iFm3�����]0[��).pA�u_GAAM��P&©�T||�kH-4=�:NE��8�H
296����Z=~����^7-��u�~>����m�ys[�� ��|2���E��+O��kq㥵����b�N�V_�&�˷�r�˴S֬��ļ��ng�����WE=�\�rݼ���6�ƻX���=�|��#���K�Yd~S���{[fl��AȤi��;4��� ���Ҋ�.����Y��-�f!�e�z��������Dw��+�V�6!�>�|��xW�ڞ���B�aޜ�a=&fEҾ%�w��H�N\�
q)�s83��U���<ٵz&���:�*&C� ��I��T���wW��t8"$DY69|+M��w�辯���?7q���cZB� �ķ���F	���᧪������x�EQ]ѓMz��U)爛t�B�6N?A�ֽL�`C���w�_-��EP�3E��N�]M�H�q"D����HI{��3w�@m���jF�$�6�ZJ �B�yx��-�Vi]�O�<S�~�k��]�.�I�+���e�_v�����z��f�Q&��{(뉡p�+�s�X�����H��B����j�"5��|Zk��$�=����+=��?`4l�k��"����=3Qx4�ܘ;��Fn&]f�V���Q/D��z~գl�S]ct��ڠ~:�h�s�l�ב�Mzѵ��W<HSUiW���.��aH��O&�0U߸qRk�SM&�i-�yxńY6��˜O�5!�Y���<�(����E-��=�~��ˡ�j��a�5�����ƩU ����U�:C}vaf�Z����U�e����(�TWTjm�*���"
j]kڐ#B�Ć�V3k�^��U��wbv[�R���UҦ���b^!܄�xL)7=��<Q`!��9�9���g���&��ز���u����(l~�I��Oj:�*q�-C�x��[����d�ƅ/o�sh�
��m�C��^*���yB�b�ʑ��ؼ�`��B�\���?*��8�o�:�vU���gy�)����x"ڋ!Mc$���.��V����<�v2�mF	p�9�'�f����э,�vj
W�����5�6*�����ٻ^D�ϢۣD���&S�Pz�)vz�dy==�����2�a�5����M�:�������p���Xt6N�3G�0������c�>!�UI)z�X�~��YNs!���86�]����$UtK��3���*������6�\���+`�xU3�UQ��#=->FnU͒i�I��z�c&�҂�i=	�[�����i�ڿO�f]Ii=K1�[�D�A2b���S�]���"��
f��a�����Fs&��E�9�/�!��]&�����d�J�=����V�����>G������r1P�E�x�A��za�����(f���0*�F0^��c������l�sE�Rm�������Z�ΈL� 0�e���!�*�>�&�N�BG3#߉:���F�4�ÖP>a;�L~iɔ��u�lhk�UtWN]jdcFsT�̚e��`٧
�i��}�Hk'�'�v�)�0o��=���ꅽ� �; �5��9A%�-�3��C��!��OMY���)��՘�oÄ'M1d���j�>0�vǡ�FV����'JJ�7^�d�K��Y��Ĳ�d~Ď���t��w)����e{�l�=���w��,D�N]��V�A����Co&~2�����d�%��r%]�9�_A��RZd�yv�L�w�|Z�?��u��f�BP"(�Tm�6yS�s�,�t�!f�� �^���e.�5�ɰ�/B6MW�>#N�ڟϷ�Q��+�MNoǐ�<�p���;w)9�T��%�y�%�w�`j8c����Y�SȔI;�ku���ܪdh��'!�l�L{���F�:�<������4\��v��E,�;�݅�Cx�./�)��.�����iu�����i-6��j_�;n��g��_>re�oJX�K�27Z=�u����7m��ڊrǂ2[��:�p����id���@�D.)���o0��ZX��q� l�bTJxs5�FN�1D~;ʜ`��j_'!n��y����XH����2��qO�к;VD9��]{zr��z����T�:9����t��M�a�:����r&�I&����Q�����up�r�o̠;�x�茪r͢}���3t& �縶��Eܕ .RW�\j7#no�\a��v��E�v�yr,�˒.8��*_?ɬ��厏zsಭE�؛�ͳ���<\D�f"�<$~z��N���y��_��Ȅ��/'�
�X�ŝ��G���Ε�B7zu�����q���� ���AG=��`ŪƟN���Z}з&b�ѕ���[ZY�4� �i��Ui7��b��SB����\���O7��6�%JZܲ`�������ycD^X�90퓺%��3��@u{=4��*#3mְ>����Gh����)�Kq�f���ex��k@��r�5�2�~���"�eI���L�E	d�|#E�vee��&�����:aj�s��[q[����S^U���B�bEN�V4�v�a��\T]�3�L�߈/�jh4�H�Zv`�X�G����2�q�-��b���<����c�l��:.���L�h��N���K�x�!��2-�:P�)�$r�ʺ�)*q	�mu��XM@n0�2M��ݍK�)�\���f��y��{uP)�� +�{�d(�q�n�Y�BT�c�.�	��2<���lz�-P�}�Y�
,�P�p�j��q����	BH;�P�N_o+w��2��(�0`�d'�9�**���f�9�U�I0���@N9r��
�������7�l!6aT�9����Bp�ԟ�
@q�|�i�L�OL1Z����H��ۢ�r��3{���]��ʖƬ#��g&�DA�V+�"��{��1�	o�(_����T7����(��#���L�c����Π�O����:��hs�\+�jZS���u�����?9d/F��<�j��h���D��U�_kDܪ�v���L(E�o���5���֐�<����\�0��k_�ݔ~�o�df��|c*��&Ҵ/�t��'����+��9��:�'�eEy���.`���x;�F���0N�wI���1RW�c�W4,����	R����kgZ����D*ՙ��fɻ��c��GX:�^�͹���}BT:v���@Q��Z	��gdϣ�q�[�2����\��+�}���W�~�<j�*��N�$�@ԑo'y�!X�l�m��Ê�q�@2�5�"�����+\�E�9"�� _�#y�N�F&C��Gt}orѰ���D-�r���l��-���<����'=�P�eq���>�K\���(�S|A�7D����"$5h\�h�z>�N��?��S���ʂ��������^�$,K�Nȹ <��/Y�<˥�4r_tg��(&���I�0qd���"���i�
��g�{"�b�o���C.޷�~d��$��3����}`MG{ &�E�25����Ĉԭ��M l�����	Z�g��.ўrd�r�Ϩ�Ѻ�gg�ý#-�M����w<:�}��Q-�b\?���w�K���d��m�R��YJk(��e6��k����KxH܎^8{���3�[�i8��%×Ff꙲T"��x޺f��M���3@���$�����0h2]�G��+�#���a�v���I��Yқ���D�q��!S}'{x�ی��th�-*�ś�w����g��@�y��V��BL�e����.B ����V��"x��˜��] �+*'�a��M���*�����#���s�c�A���Ğ�~u���Y�ۼ�1��"��Q�ǂ*0�`�H6��%� ��𲎔�N�����?��ap���)��P�}��	����|-u�� ue�%��I1=j:8�~v���[�~d�T�*槣�c�EPO���X�L�n$�*4Z��o쳎o?
Q�T��|HA���ˍ�oϥ~�g�;��2q/�������\�_Ey�������P8�s�bɻ�ĝ�)�0&B(�E�z�ü+��-/?"#�E���[5a��%�}ZZ+ e"Doq�g���'Rm�U��*�����U�Gb$X	� �>�͔S;Y�`$��U祿��r <A�r2��u������#��̇9��W{���"�K`.Xfa[�U'ٜ��R��bh<��{���
R���*�* �L?>]��L:�Oy���Ot�^►1��b&(��*=G�6����2^~��s�VM������K�1�X�����|��0X��9�Ogz��@!ޜ�0IJ������M���u�}['h��ow&�_�hO�)��F�_�d��
r|k���O8ߪ����CF[�E�	�J���!��ʕ��Ǝ�/ɽ�������ukך�i���b,� ղ�pkB����?���x�tu�DЭW�PH��1'������S�R�$xxU(O|W�Ş��Db#i�����<���^,���Bo�"���HuA�2���#�i��F-YC�!���K}�.+A��P&¦�����)!'�ȡ>s�'9��ݥ�jNsO��QcC��5�eI�pO�◱�6���Q���`��	�rLaM���m�Ԁ��%��lw��Z��c)ϕ���y
L��h.7yz��Q*ɍ��S��Q��l�}�XIe��Y���ɩM ��i�e%�4�y�_���	r��LE��E��!j0���ɲ��)��S������`׆�Ǳ2ޥ������d�,��[��.�窘�J��7�߽���N#eRǢ��ɳ�8��>���	z�q0@}����j]��l�t>�)!_(VX	ݺv��V�4E[�N������3 �������$_�.��"j�����Jd6^��&�~�I���I8�H@$GT�&�bˆ�Id̲(6]����3m�[�,(,I4a������DT�k�?�\J���=��(�K%�:Y�H3�u2r}��h�׼
Q��u��m� �82"����%��L���%M�����Ċ8T��Ha}���[U�dX�>.�6+��'��tN�ʖO�ٰ�4��ƹ�NJsEa��/��~&��W�������L���zD�!�-i��1?�c7o�aR���:�SGg���pY��C+߰N��4���m����CZ'��N�I܏�_��4�i�C�"�a��Ä�$��Оqn���Yg�m��Z�̺�����'�{�V�+��f���{.M�7ʷ�G���135}^+��B�z��o��ڠ�Bo2g{�>jwb$��Q'�̐��p �7j��PX���[p��r�Aw�5e��M��W'���������b�1�n)^[F7��x ��:�����/iڰ������k�o����A-�\��Ǳ��؋�;�ͷ�pK��z/{wk�N!���V��Ҹ��u)i�x!m�������A_�F!s����?�?���_����G�/9S���ҭ'���8�������N���H1���?\��7�s?�$��_a�}T�����\b�l�255��7f��
`y^�N~��g#�m��r��|�;]mdĠ��myy�����NNN+�!��1��k+�h�����Pt��eT5���P�/���b���/��?�1m���������_�/���b���/���O���˿p��RCE[9�����PK   ﴵX��ڙQ� � /   images/a16cea49-f54a-4dcc-9abe-0eb2facfbaba.png  @߿�PNG

   IHDR  v  >   �U;d   gAMA  ���a   	pHYs  �  ��o�d  ��IDATx��y�d�Y'��{of����T�J�ֲdI��W�[�L�hc04��д��LL����41A�=14���3m7�m�i�^��&ٖ-KU*��z��%�{Μo;�ܛ7�����8Y�2�.�����W��_���y�Y0@o�?vP����;��9\�����Ϧ�S�[?gY�Wߥ�ӱ�u�7N�1Nn˿ۤo��)���������L^z=���څ��|���crۃ	;��A:�M�Z��`�߇�_�2���}t�3]�_�,K��&��v�P��=�.zy�<��s?n�S���;�|�L���s����yK��%�X�'?��]�2ޖ�����g.K���>;�W���>$X�>��hC>1	�Ն2���&o�������_�z���O~�B��Bwc6��`ۿo�����2��}��ڂ��MX�܄��i��n�5J�G��^'7P��1tY����\|�V����^�t@�x��8�_����4��ߜ�������؉p�m������W	�����ua���e2]��wqd<�z9�Gy5Ne�Wt�o��c������U�������h����p~K��O��N�=���2�����1��a� $k2�7��w�<�8~���k�^������ �H2ʽ�5��s��FW5:;&|~7�=n'\���1�7��q����M�<��%a�~�ݼy	�;n�}�Ji�����2�p�>��\u�pq' ^��φ��������=�B �C�wAK	n(],��'��$�w� E�����!1�y��A�|����]��g�{8	S|��UR@#h䉝K���1���,��3'�W-.R��	 ���6\�Z-���e���<�:�m<�#�����b��}z�7VW��z��]�ۛ���'��?"�<4�H�>�7N�G��+�Jt\�G�k�<���nX�]��N�E�~�q�+�N�7����c��OLM���4t:�𾽽���+��8��4�]<D�w%�����We�t�A�9?/T|�x�۹���"�h���2P������RG\���}Y�'�L��c7~���������,Wd���]</�OvEwj�Bv#���J��h)��ȸ����~�sq?����� �\X�n�4�4c>�y,����$��"�O���\�c����PO��.'3���8��}�B�u�`<�#�����2ۍ7EfW�NZ�բ��sD��(U�{@�5?��.p��	�TV^ƺȅ�&�>s����p��L���q��U	�7s\��S`��th�K��y�3��9s�}IW��y��3�pZ��뫰��L�v�A���� �Ĳj\2��s�[ݞ'ƞ �%��"�g~qe�1��8�y��=������c���L���b��i ��\��Bp��h����ѣǡ31<�^9�	�!�_f��b�3��ҲLWM���tEM7��+�$4?3	7f����U �}D��3Fqݹ���J�~�zt�:K�H��y���d��x;c0W�^��	�d�,��;A����Q?]*��zΘэ��	���!���bq"rEV�dʛ��d�׿j���:���'�L��w�T�L��I�� �r�	�d�s2)�~���a���Z�6�t�X��[�@�{`��Px.4xΝ���_i��6�CU@��"�FNd�T��l6�� �=Ǫ��u����#pS�|���W����c	$:�AO�@�B����%lu A39	Ґ�J��!��-�u{x'��T2OH{0�@��/��A��Fn<�^��9y�����D���i�͟�v6��A�_�o{�K@4��	;���X��:�0�u�1���J3�׀�\s�p��q8t�������c+�B�m}�����q�-��9Җ��� �'�{]��L���(����+\\@������{�Ҍ>�������}M���%��'������"�O�U���&�K�/f��N m��oF��4��rYG�q/a ��E��Vu>z�f�p/m4G��Yc�6,f���,��|d}��j�K���A���/��6�Z�۞So��s�v@�J�x�x� ���0]���U��8^N��Β��>��*��״�ӹ�����Pl�oG�uԅ#/mf����<��Չ��	����9-���u�A�T2�En�'� ��s`�7���s��ۆ6���rs�~��`HZ`����^V/�6�k�h�Dk@w�t�0�PՏ�a�_������a�!��'���>D�D����1��E)��Zb.u�ӳ�0w�(��Z�[?v�(Lxp�Y�}��;^�q�G9����l]ES]J��n3a�����\�G�5h�Y5j�x^�S�0=F@*IG��s�n̋��'"/]%5k��[�j��1\;LX�X�qnK
F��>��L�@U�:�q�F�N���{M6�g!��Ǡe :zn?`Tm:ŭL=^kA�A]�d�|k�����8Y�`z^�uRQJu��Z�k7Uʭ�#����Y����T�s�v!.�ܱ^� H�M�"�Ғ��yHV���pA�{����!�@�oŁ��dq�I�`���7�- �u@U₰�o(q��fX�$R��k���t΅���ј�c�R�R/Jt�
��d��� ��p�Q� ��)����B���3�����2����΋����;x�	�v���y1*Y�8Ҫ�q����$Y�~�2hr6h�V0nnoCO�~�;n0'���Q�d$ә*���hߡ��E���N������a�s�s0=3���������	��1`�Ze��/�9��"+�	�U[L)s�ٰ�M����eq��bd��Q�ɋ����1�>n�,�f4O��%>�)0�(��h,���9�r����~��M64(�3��4�ǆK�̍b����h�!4l�l`�͢���U�{(�Kv�5v.�.էVt���5"�'�l�U
�u\O=V���"�A�6xjïzs���-l�NY�"�依p�ȉɫ �s@�a<�#����x�Ւnݰ�L�~����AW��)�;܆E����ޙp���EB�vX�{�\��o¡���TՆ��\*��K?V�$�
�ح�R ��X(
ҹ#q�u1�f��	!�,s����`��M?��z]��󄶤��jQ��4�'�?y�%24d2C�"z��<:6���[	�5(Q�QwoX}��t�\Den]�+��)��My��"�Tg:s�09w����^8�����gH�*0?v��Jb�
��`n���ՁK��y����y�{�N���[����hN���τ�GO.5�k��^8�W�A1��j�`�
|�=��*�C70�;4~��(e�s�O7�V��G��1��H՘���0����>0bo3��]��:Z#L��0E�y.T�F��h��D�$W��H��.��d`��b%7+��: $}�ϑ|�ê �t�V��%���9tN!ۀ �p��#��&�$}/�����	d���&�c��~���c����<�qT�53e�06�m���)	�u�dXYP4_6[�
�@ΏǠ�`> �A��~����H��n��EϏ9z��7�2�9�ޑ;%oK�K&�ՠ�	��u"���fЅ���2��}���YG셁)h�d�7#�V� PG��z�t{���s��������=���ֿ;�Ǘ
 �&�B�����y��s�w��68v� �����ZY�cӶ�E����f	��]OX�	؟z�	����9�ǧw��<��W�����(E��8�����]��[�L�!k���R����Ll�� ���G���C.������Db@�O�d �@$G�B_����_�p%ş���X�%��q��
�>nS =��Β��<kT�Ī@r�s����=<����h�c���M������7]9H�֊��Dzzٞg�E�r�$�#���T�p�觖w1��&��Mԟ�U|e��R�O\��݌z��w;J8�F�/��\�p܀ג �`P��ĝ���?��D|���DBd	qXʲO Hn������-kEʤ�����f�7Xύ��!�8Y��Y6���MԒ��\+Q�/tuDp�OS�q�Q� ���c�<q�n�D���4��Ӟ(�p��;z��p\�6�$e<s�	�,�����Bws��Ut���33Ձ;�8	��}��~>�W����p��8r�(hh$��H�w���De�@��bF���Ū��U��?gBpZ�Vs���x�0&��-���i��
"�ezM�/Э0SJ�"CY��@�*���q�}�̲-�¼�	��|�g9��I�#�K�͆u�"ɡ���?�!F��r��g@4����]BM��	�L��O��͂��>���%F���ޒΖ��t,
⦥A����3���d���6|��b�Z���i"5נ�Q7�nlY� ѣZQ�da���G�K�1�s��!���b}��5����\�{ȩ3�3��FL�X�(��o���m��Q�g;Kx}uwT��8�q�$�9w���s����d"!� ^N|�i|J||���� ������I��G���\_h|E�?�R�ԩ��:��\��G��ЁIx�̳�[������:|�+�G��/�̤�����8y�Lt2x�/�nϏ�9 �.���'��_������ ����o:
�[�t�ܰ9����8��Y׼���-4J8X�_a��E�~)��$I�p b � G��?Q��5��c�L&@� a���v;���G�Wf�X�B�#��?!�C���U�(H}�!qC*���0ܺA|O������$ �Aʹ�u��]� �F��0��:8�`Bry� 8�*��C/�Q����C7x�0�P������3$k%��^���j8���k
�F7Nz���tѕ�y�٠�ZT�#Q��µ5�Բ~��f̝ ������K�$��:�c�ɺ#��� P.[gJA=39qu�r��1���g�����BA�.�釪�<
���2\����b�#�0r樚�"!3l�K`k#iq���ۓ���)���S'������uu.<�8Z����9l~�G� ��d
�hAw�'(,�@��Q��ԅ����$��{�?z�~�-��?�(���~��U��G^燮�α��*��|ܰn����ҡ�*�PDh�v{�$N��U�z�8���f�i�v�t a�$���Lpw����+�cn�����$�jbZS���n_TM2�J,��7j�x���;���(A�U��5Jr^ԷG=q�=k�0�ɰJ��h�l���C ��FTI�,���BO�r@j�B�}� �y������rԸ��H������{�t��l�C�.����w����q�3��V(�O}4vF��J�P���Bnx%�;:�� 9�Vz.]��P`�x�(ǆR�a�=J���@.�e6�%�_��_�&��A�0���A�XG� [5Tٸ�Hm@�H4��v!��h�Ew�1Tݠ�#E��{��Q���������>_x�iX^^�v�S��^�0�\��Þ��������g�@�:�]�c���!h�u�38XY�D��	0ч����=|š{���
���?�����v	�O��K�h|R.p���ҹ��ܸ�,��MJ�3�������7]	�2/�W&�\��p|�b�%�D��E7��.=�;�ΰ�α����5�f����i�����L_����wz�c)@��Q?F��'8�G�q����hկ~��8,�����6y�X�)ϋc�*��!nb�
��̈́c��R�q]P�,���%�
��rL�q��DDz��;� A�%�.�h��p~����:�Y�i��`&�@^t�x/��e=�~��<�r��q��N��E��s ��� 5�xNM�}RW;�ֲ�r `�����e����1�3�H��"UN��'7,9��R�s�~�)�����o����؅����a��#�g�ץ{ c�0� s3S��^��\��g�+��1���%�:w�s�]�X_��	߇~������u۞x�~L�yN~VW{�������g�#���_�%�ml�+^�?r��14OD��ʩ�c�����Tps1��]4f�)n8�yjU�����⺠����E��L�{ c;���°�~���~�<�
=��2>��������N�߸��aXVE�:��}X�T��i�ͤ*$\eI{[^F}�ʒ�2�&���'�xFJ��3I5���kj&P��N]��e�5w��4b� �zM}�wE+�gQ};�2�=Y�zq�)hD���'�oó�+j�-�8�:!GB��m쮦�ojѱ�^3�c��N@��N���>���d9�6���a��{�@��Vsy����5���Y��&HM(���m_ꑮ{mc�u��S�07Mv�˗΃뗰��'������lx�����<�z67=�o�p��a��;�k:��0u�'w�-�spm����{�������0�Z��O|�����ݯ��u�'���,+\uF�'H�ɑi𒮺Ե�>9���(pe2�{�y��Z�r9%�%���@d ؗ}���n�6JSQgdG}�Q�4���jr��d.X����|���} R�[���Y���m��n}Hc#h��)��T�B9��(�Д\ įY0���Q�X�fi&��f�τ��Hs�	�4�
�+�Mu���J����03"Sy%Dʘ���-S��zj��$�n����q��0_�x���	b�k��J�:Wm�Dz*�*ҷ��X,0�r��%��
��~�!Wri�!�@8(�/�Ҥ�$�����ܪX�}�A���	�~N�%V9�@E����,c.
��EU]������O}���a������w�^8���Whkm�9G��v;�Iҗ�/C֚�D��;��ma���]Z��ǎ���{����R��:�9�`jv�����ԭw�/��/���ۿ��p��3���x�*��Mo�C����m]�K�'��;eVT��g���_�E+X+�aX�a���E��j��%ۂvV)�H6q�Ym}֯Y�e������?�4kc�|��EJ�1q�Û����^2����F�_v�l2�*RhH�Hcj��ِ�a\*8� ơN8~`΃�EqyD/�7#���Bʙ���j�CN0�*7j�z�⦡=��h���:�''��eP�br`}�F�q_%N�"���?N�(�S��������ĎZ�d���a*\�[EUHQ��5�j��6�)G���J�x�磉F���57HA�	Pٔ[�ĵ��[дe�.&�
 R�R�#J,F\�E-CQ {ˠ������.å�eX�nA^�FP����3ς��`��F���6LOy.�S�s=w��^��V&���,:0=7��<L}),���˯������rv��}|�+_	����^� Go9[��מ�[����g��oۋ%G
vYU5��#_F�'Q��$ˡk@��}�k��� ����WK$��M�֥G75�O����C�U�7�<���AaT��Q��Ї�0�W��B��FF2��Sfi����GS%�.֤����*|h<�z�ڭ܃�lP�*�4ę��DuӼ�Ha���y�mE��h����F����VƆ>0$�#��g=����� �.(�HM��^��b�,C������D �:����	�s�t~�m��e`��ϭj��Nc*��K�.��������D��F��B��J�H9����1j��\W0�9����4���'�N���WV�����x�s뛖=gr	�6%�i}�xv<q���[� L�k?zn�����a��޻�=���"d�6e��>������>q�$���1H
%F�������������� ~os�_�_��=��KF�VKu��"��Y8V�����Oi����M	&�F�$�$f��R����cN3�_�:\��zn�@	FcIYG[�����11�ڻ00#e��`t�`O"vw�ԭF;U��YQ�d��,Ӌ�F�T
��Y	t�E�Q�Fr�K�]ǋ9�E����4%d�S��g'�Q�De�� �C������k��}��H�#�\�c��1�^�K��H���M@��N����4��#��@�Y��%΍Z��p��s�k',T�_?#w��(46E���,�<Q��'3���l�]������X��ȭR\$)�]���܆k��^�ˋ�aqy���������� l�9�l�^)��ma�>}�����ԩS���	W�= Ov�̜�2��XȜ��$��&��Ox�bbfg&ar�/��V��w��ݿ��hO��������ŋ��c�=�?��z/���,�Uj��vD*7�]s�ۧg z�E�qN���D���Nq+̷s��!N>����ē.�7��̝h*�fd��=����Q�����5`���y���5<�9=W��H5���i�k9��BE"�)h�C[��e���糮j�Kf��画W�����(BYQ�h�ig.^!7���A?����<��8lZ�YF9?۬�n��=�ϖ�sH��"Pd=� }��#�T	�� ��2R��Ʈ�������%�>�Q\�lL��<��9U��-S�?�%Lʅ��w�?&����L׳�g�YL�e}_<���������OHhW�7H�r��e�x�2�on��>r�9F㖬�G���$��T�������v��ep��;<8O�*���a�	0��握`8R���͟?��A�F������y����Sp��U�9��/�S_y{����wB�K	�+L��j��]pJ��t�f�5f�R*O���������d�E��m��s��HaKҤ2M62��F�u�#4��ø�:4�!����]���S�F���U`d��{��i���od��<��cJ�b¿(��ȯ�Z$".E����^�@�y����ߥ�sεu�KU:)�ɤu%�b��)E
e��gշ���	Υ/Y2��2�h����}F�ԍ�3���̃HFYh�s� ��\ҵ� N�h��C�����tӆ�,m�T*s�H�S ��]t��	��E��c��j�z8�9z�]���x99*YG.<VtSb�������3��ke��ȇmaY�)�E�y^6�6�̹��穼�vw��1oL1�!UF��}�r��.�� ��J+/���p���p��a8y�E����|8�紋N�w�A�E�T��c���Ql���4�̳D<rʱ��8q�0������}�Cp��5X�v>��O��~~���G�z�V��4	pP��?���h��cM�V�9��@��Di�K+�[]�:�=�[����%J�.H�U��D a}�>Ĕ����<7A�Z�����ou��p���F�ta�H���СA���k+�0F#ۆ�/�+5�ɍt��>h\�Q/�y�b9-�Z�S����%�q>7�ѩ2�a��f�!�J8�U�yRoOG�Af�5'`��.��J��ƣ��r5��$s��$bK�_֚d�3-�Q�w����6'��m��t�ȑ�[�-�w]phJ4 UDҨ���VhQ.&�@��C��53�e/��jTSU��z��R�d\Ce�_�H��T���o% �z�㜎f�c#�.���}r�)00��kd�T͆�����L�d���(̺�H�^��<w�=5���p��h?����׿���ȑC���������)8z�0��-J�;���!p�LNzN�#�f|�ؓǏQ4j��^W���u�(yYgb2{}�߃'>�8�^[�����~������������pK˯^Eq呂	�t����e�h�j뗓������n���X�o�zϮlw{�kD��9F&y�H��d���r�2Q�����e7������m1l��uiZ�'Z��Y�U"��2�~ݘ�0	�0�Tg�5f�)Õ�C<F���؃�X���beŖ�>��nnH��G�b�[� �w���.����&.�9�3C�1�����KP��ʦH��)e� �#'����	��t���I��9ux�>p�;�L�Y����ȥw��$��-�R�x��*L��1G�qQ`1<2�y��>%-H�} .�.���h?��{&��I��R�]�����h�Fc����Rw�U.�F^$��s�D����8[~#w���3gᅫ�ط<����J�L̼�{])yN�\V�XI����ȫ^��g~��/{.{�S0P�[�Nff�)��w�l��&�9z� ��NM�V}��BL�&��5N
q��wK���}azlw
~౷�����_9���֯/�����&,LM�> ��uȊ�Ȫ�
��2j,b�`�͕�:���c0�6��΄��$��F���'������W�6(J���Ċ=�����qU8k7�$VT���Qj�]dT��s h����LMO/҃&H��ZL��O����O!��	����W,�7H)��tf�~��Q�*�p�@�Rx��8����64q屷)7`$F�s=Ł� @��F�w��;�(��P���C9|���\ژF�p�\���fTW�`��d"AWD!tC�����e�W�
��m��}#�W1W�m�,��w$"�'�sM�j��*��g�T�c�K�i*�V��6mt���6�>�ߗ.r�6��Q6!�c�_r�ܳ
�P��4�l.Wե��%�ϡ\O����Ϟ���X�x� �z"ٳ}&�����h�)Y2�����(�c�u;vN��Ν=�9�6l���ϭ���PZ|���A*���գcH�⯅#�Z��"�����r��(e��zZ\
}X��S�)x�a��/�/���i^�|�I�������Sx�U����"��0-��PF�%c&�$�\�Y2vSu����&�8x{�奟l��`ie�?WN\=���7�)1���2@8YVo&eb*���r�?O4����H<����k�e]: ��^WG��}�c$<���C�I�+�[R��u���W<M£�Q�1� F�^�Y�Ć~&�ӝ**�, f��a�]@H�Q�PbS���\�FN�����w�J�L�8�P=�~���:���j.����K��������N׿{��F�7��6 ��<$�����8�S)�� /�j�{a��p��fċ.���h�U��*�ŸR'�7�8H4b����"���+�jIxS���4e��핣���Q�'��u��Q�=qֆ�Fq�r|E���e��XtW�h�Z�'�: hTE/#�����꾧�m�S������z+=z,p�G���9ρ�����;���0��0,f���u�A��e��Ih�X�z����}'���Y��?�SX�~8 ��_����I8|� LMN���"L�'gb�z^[!�����B���M�V
xb^%���N��c���uX[߄I���� V׷h<�8��-�+E�,�UBK`��ע!r�U%�q��*N5 �+�=0��.쏰`��0�:���R�Ԏ��Ya�g!%\1FmJE��X�Űj0�8:\hF��I QW�nu�]�_��Ǟ�{��Ֆ�N��_��'u*L�[	��]�Q��&@�xr����H��/�J��eا`�gy�tس<�Xl��k�E+b^�q
,��h�q�"r.>��U�6,��� G���Tb�A(�"g��L�auPy!k���U��G����t��D�W�~�?��Ś����pN�
}⫯+Rn=Y4�K<�N�Yz���O���]�s�.�E�~�s��`g�T��QT!	s��Ad��WP�,�==݆^vz�8����#�+�� :E*��i�3S��]�=��H�x,���AYR:��������좴���Heu�=w�k_�x�g�ܹ�<1�|���? �;o�c�ź�m��D���Dے����b]�,�|?�-Gj3+�wp�N�v��d���i{"6	s��O^*��U��}����?8�)q1s�2���eјiE����E}ص kP_	3'�fd+�i�W\\w45*�0^z?����2	��z*��L����V̴s�HE��r��Am@�d@R~��vr6
*�L&��ڣ}MC�U�;���*�-�h��Z�e��Y�����>g�i-�#u�#�?nR2�ċa�ֺ���f�2�)(�T��wBj��hs`E�Lbn�����X�9��g�����s�@�����`���K��,�F��߬��(O`X��*�*/&��A�Q&B���e/va��k�H]��A����I>�L0�kH�Fk]*ha��U�\z�>�MK�Ą]������	g.]��\�K�����ƕ���I���AA�.f��,Q'ނ�o�~�!�/���$UtZ����s��L�t�+lS�9p�/7:��lI~�Aϫb7r.��~�[9���h����z��g����х����������~��׾
���y���[�܅�~����6\�r���쑇T��K�WOFc�VA����FCo�kpu�l��4p����'$���T�K-̔����D+k���Ճm�� �4a>Q¥<�\��� ��|F�\��c{ʩ[�ۆ��MRu�>�s)�\Vd���3'��XT��&\?y�ey��S|(~b8:�@_�7�HG榨��r���j�ɱ� �YAn/���?�Lj��ئ�+ȥ�q~�>L8�9]:vڮ���O��VP�(�4σ��F�`�$����`���ɠ(R�);Y[�RR%�=LM!��;�:������h�҃Fϋ�/s�����L�(�����U%1�/z�ˆ�\|��9���B_y礠3s�������4�$!�P�Dv�Fdېʃ���5�	� T��D�:�Z.Q��IUFE�As�P���$�wyy�~�q8�}q}6�����܁�T-�2��ۆ	�G�����~��,'��ӝN�\8*X}���m��k�����h���e�	�l��V6:��M�|_Q���㜬�P"����%��l@�ۇ��Y���y�'Vp��st�c������p�Kn�'�|B�����Eydb�K�|?�a���>� 3^� q��5E�_C�ϥ���E��J)k��.����'ar��	�lx`�|u	����3�P�||���R�_U땶�V�M�Қ>mƩk���ձ��!�;)hdnʘ�$U�X����e>�z��`X�j;R}:(#��	�3L�&�b�'�H���\@�i��钿�=�Huv���n>v�;�O��`G���6��
����;N٫B�f�C$Ϣ>=F���A�*:�:�h
h���'}���Ņ�wT�<�������F�K��wD�*=9��w��JBV"م���/��n+@� l�^(�;怢{����%��X�	�@�=���3*`��@LTзC�K!�DWJJ˼�J,4K-��S���Qx�D��[�G��=����z�+���O�Z��y�B�y��Rܔ��WV�(��SG���;�e��^�Co{f�5)w?p�p�^VNeD����CM��gځ��j�X��;Fzb^��n�=h�nl�z�T�� �~��P��xy�;�z���� _��3Оh���ð��
��?oy�-T-*�A��*��g-Jf�z�����=�rm��m�S8�0O���O�>8yϑY2���i/�LNv`ʿ�<A����L�30xt�D)��`�[дdB$�ˉ����+ �HF�n�kdCB5e��I9m�԰Ġ�� ��r�i#Ul�U�2�,�+ȇ �<r����ͺ��.���-����y|nt�#*LTio��;(�� y�KR��3�e�OF=�e�=��CLl5��0��	� ���K���1Lˮ9�agV 9*�����ت��X��d����pR<Ը&)�S�S=�z�h�sl�Q�G� P�3��މO����j�2�����V�Or�}��X"�TrN	��Gą�g�0&R��3$��:�M���A bz����1�9���U��t��,åkW���)t[
 ���߯�yZ<�������>?����h�����&Lu�~!�B 1JPu�;ۗ�L�8E��Ab������I`>љ��/���?�y�걢ֱG%��=��S� �Y23P5���&��g����=�r8��9J%�@T�ן9�?xf�ft�ݲ�R�����)���%���'TXL�v}�7���*L{�6�A~G��)���S
�z����d� Lt��C g�l�<��Y���uz�2������:v�D����2I���ɸO�tͫ��\�ZL���i���oB<H�h#� }���\�%���G%Rץ���2Ekaf�D�B2�3����>Nど�^���	�P�zP�N�W�{?����҆�����$P�xP)�ax�5�4`���YP��˱��;M��Hז�%(J|�3W#�5\�3��z��P���"�mp��������܈rB�L����G���*5@L^��䑁�����'?�<ȌyN0!:�PmQ��I3��~Q��&�H��d�,�z��A�ݱ�{������u�z�<��r.\��+K������F���>�9�m&A5�b���#��-������/��7UV2ġ�$�z�V�"0�>82Ns�|# �j)�L���_��KK+��N\9��}�纬�
�#�MLNB� a�'��c���ã��{�_<�x��8�-��s/���:��/��&؍2�g�H��[N�$�|5??�,0nzuc��	�v�b�^8�3���������li��X�
ϛ���b��%Lpv��9Z h$�uSI�R��U\�����k5��\X[.�$�z���5Ի-� k�^Bbq��V*���r�z� �g�DT3ՀK�1��=�bڋ;$b6�<�4i@޸3{�Ek�X�+�u��9vl</��p.�J�j(��@�Fq��$��Vkv�֐'�ߥԟ�l��J��:��)�ш��b��(�!�	4L��Ј\���>�]��Y�x+�A=!���Oi�2��W�bj=G�K�Ω��cb�!�(O������b��n�j �F��\�c��`�$���E%�cH�x�W�������_���%X�`���$�*����!5�,�8�.nfx���������KZYZ���Iz�*��E��R�T?[ �5ˉ#/�6�@�����34^�`��Fo��s�`��R�\���EHU��s�U�R2�HY2�u&&�<�؂�n	|���VV�����p� LOw����O����I8t�P�^��89���N<���P�`��"?�w�a�ߥ ,�	��Xs&���� � M��D�,�`�$Z�����������,l�����9e��2��˔�Vj�Sǆ}����Z�F��>�����"�#��E'��j����fYX����0I��Tj�V��
/�+�7�l�T?�`�(Ǌns/�l�28�=2��pk쵑�����g	�bsEh�׳_��J�1��;��+�ӷd!�&���#wUr�ԙ�9y0P�	�Ɖ\z�$�N��2�l�N�	|������X&����{�K�I#����X��.��ڌ���R���Gn��6��2@�6h��B��*J+cb��,�PZl��Ξ9�����'�|._�Lj�~9�HR��ff;��ڀ�M_�E92�^�����������n��Q�~�s�tӘ�A���(J�E ���mR}������V�8�m>�*��E�����ƅ�C��0��/|����x.&#{��spם�ᮻN{ �� �B�auu�y�98u����f�E��@�Ti�M�"X�X��m���yH��AǃuI9����}��8�5�`����Q*�LN�$a���ጓ�a�m��Ā�=�0���5r����dUF�=��"C�B�(~4~��9�� GwC�Y�c[j8e ��H$��Vg���c�TV׽'ר�����7�lPU)d����V��t3���^8� ��������< @�ƽ�+5�O݂ոH����DC@�� V���Tbu�	�]\�r6x�B��"}U�N	�Q�!��!����#F�� r>:24&&ia�p%��L~D��&����wr�u)RA�WbAn���QZ���������(w/5X�S��XQ�<W����@?��Oõk�`�7D�XR8L��y���`����p��[����C>�O�
=��#pM?JQ�ny676Ʌ�b�3��՛�g6ıBq|'W>�k`&氟6*�3Q}�#h�n���YK�qET ��S���sssp���S��k���%O�7p���L/x�\��{��VA\��o ǎ�{M��9�<K����ϋ٤/^Y&�n���#����4������X�IKb@$P�� �dl���h&bN�-�D�x�������(��������(�7�ݡfL�T��=f���!�<5��-)M���`t�#�"W�	DP�豬JB�63�p����vkZ�F]]z�k1�j����ѧG�?]�_W�� ET�UZ_���$���V��t/E��tAeY�'0�΀m�9��h���ž����*	�j�g�	��CB���G�L��B>�$S6���L~.J>�N.^�mڐ[μ�=�!�8Ι�Y��a׃����s_�<|����/�9��-V��K��Q�Rb�<��p�O���k^�*���p��A��mV���ʥ��Bn��ewD`?k�k��j�A�/�����T��-�!C��J���R��
�0��l��y���0y�1�p���}������	���̙g����׎�l0O�3P/�\�6�Z��/�+�2P�����][�R	�R�E%���z�_7���.E�b�@Ls��g�-@���3ԇv��a�$�w�1&�	�Z2&|yƄ��s%*<,-��k!qހ �Y��S�x�j'\/J��ܭ�\wh%�q�`qdٻ�ZA>�I�z}��~2��X8��j�swkC��[/Խ�k�q
�艍�t����k*0��>����%-7$�aW2D)H3��K�2%U�FAS��2V}D�h5��h5K��p�~|X<��d�5\�7��rPY-!�s�z��A��U	��Z	U0���<w�姾����c����������Ȑ� �t���0�Yэ��x現~���|���A�tT�llW�!����L�.�p
8���h�gqEH:
mh(�)E_tLM�4�n19�^��h�jw&�nJ� 隍'���B�X*�ʵ+�է�����",zi����._�2��Awh։�Z��\���율�6F�t"����+dٞ�=��O0�;��0%@Ci
]D5���N�S� �����D������A�����q-
a)�*���A��N�� ���C�nT'����w�׍Te�5i�:(�:�i�B�f���oث˸�"�JEG�����;��]���;7�P)�  �o�
&����y�$u���z@�FT#����gHA�?ea���%��\3�����8���ɢ�M�S7�\P٨���:r���+FId
���qA��ߨ�l0`���(��*���Z�$�@%���*��IN$�iJh�����+�/�3��W�+k+��H�>E5`zj�8�Օl�Ly����c�=��zx������#�(�Y�c��\�*�9u��������}@ ��@�'nM�+.Q�T��,"A)sU�6��Vr�l���HHQ�H��璹�;<�~
�{�,u��k�+�� U%��݃7�%����6זؗ�.S@��C�s��h8�^��@r���6�f	���ا��`b�õ�L%þP�v`�sѷ�}��%��s.!�kPsݮ�l�f�bVuij�����^p<c�=�D$IcL� n��D	��I�'��3�*XLUCiJ��5�H�*���!��Y�7�>�U6�0�s'�I��z��NV|�M�v �d��ϻ�g��q i0ζ~�] 9*L ���꘤>1��#'y&����s��+Qr�B&���+v�ù�~�q�)}f�� ��*Y����_OLN���-8��3p�����O}
�=s��1�M�y� /�_��ޕ�2��N|�kN�#�?�#? w�:IQ���1`��܉ؑ�99�(ɦx���qd-�dX<�>�cw�+
�gԩ"�[���Gm��hk��=1���	�9����ᕯz|��M�?Pָp�0�M�"����ƊA��)Z �'Q�d�VT�*jU�"�A���R�s�䝇�{��w18*'�s4���\̷�!!Z�"�
��JI=@6��t���{D,���,���\�I�1H~�̝��0�qiL��c�.{���fc��ҏ2Q��� =M�
��
/e�J�b�]xV���iª�s}!�8 °(�[��wpWqW3����
��b5=�^���@�+"Zj\6��XX �}OOl�b12���"���w37�\y�*�=w'����� 	)����>|��O��������,�,���:ϫ��
��qq�~��x��z�������+_� L��d�J����V\K�G�$n�jx�3�p�"�M��D]|(w�$���q4�#u	��T����2Uq,_�W§?�	�p���xΞ}�<�u���ͮ�.R��%�h�-����S�����J_~FU�8�� հ����'���#I�}�%��G2[m/il��V��A���r
c�����k_�gp�yR7�����6��c#������n�i��J$���IJ �+��S����p?��+�fu����U�O�Q���I�5�Q��8��b2�\w����O>���E�k����,�\�n �,ј���G���p��w}Ϋ}�D�Qb2��x��O����60��Ƥc�-��9�'�6�x=���xD���<w��9{.\�H��س�HP�[; �� ����o����=��^F\i���� cKn.ޑz�B��A�G�����sp�Y�H�N������*���vk�W>�(��#VEe_��ĉ�p��q����?s�Y��W���~;���X����!Q�)�ۊ��%��ie&sP\S@Are��8����$Q���wϹT ��ފƁ˂��*ݱD��L�"Q���EuTiS�� �uUL�>�A�I�6.۰��0\Ǉ��.F^��V�~8����#����r�a��ω�\m�C@�pLz����ޛ���і[ӈ+�Õ��gU�S�Tۆ���&�Tfh,˷��	G;JM2nS�\���&Ѝ�����8��tB�1p��야�1�C�?�_���`{k��L��`
G;�W?~l��`s�'��zx��^/�.`A���#i�H�7ĉ��6r���/��κ]-�B�����*�d*;@�e��@=�b���u��06L|��Aҥs���/��s`�` ����-U���*d&��i����R�.�HH3��� ��O#Mu���Aw���2%y��������q⚾.�y�{%Zj��$��X���p�`nE*�J��~��'MVw����F`mTz�a�D����HAXջ�%T��շ>��,������A���Ӄ����.���q&z�7��-UwQ��h���ܑ�|�����AB��ԣ�j��F	77�̻�{PW����O|�����~���0D�K����0�6U �|q ���F�W��/��-G��͕52P�Ֆ-YO��r���}δ����҅b#���%(n��e���kC���Z�0;C�Ç��DA��Vu��6,/9����7���/}���r�\B�����[���Y7��gKY��͂{��x9AlxG�<���[Rߓ���9E6z봠��W�\�
' k|r�8�|%.�)7ߤ�ƵTT�L�x���PUU��K����Q<��ę!J�"��ǎV����
JI�����aAfYV[(�O�����I��s������X-��|����:*�WnC���wN�\�B�W������5��];q����7%đ3ۭe��(bG��inx2��2�(vc/���t�x����h�����[e �s��]r�Z{w�]������}�/����ޯ_���͂�1ֵ�Kc@6`�:�]22p��$q�.a��K��kUJ�z�i����-]�u w��;�_���{}rb�{�}03=_��e��_��~<.yp�Wz�;�
|�4�8v�*�5��5��:%�@��(���Q�.$mDI���H���ru�C�
�7!�Ӝ~-�n�}�W�R}t�� t>�<�.�&jjc��Ӝ7N�FtYFO�r]G�)�0�����DGTC:��-'��)w>Z���T�10�߭頍%�6� ��庚6J��� w�/�ݣ�=$ N
����뿛 ��N����S��3�o%����>ubE�B\ߋ�؋A
�'FN�?�s�_���z�T�o��\��b��֩�ԭ-�W�����7�?������"laؾ���&&�X�GE4Yz�P%(bL�pŁI�p������fq^A}����^�u=�.W��/-Ѹ�8q҃�,lmlQ�M������"Q��O��>r�D� ��J���TR{�OC��x<J����H��̤�G+F� �ս�:�
�ufV�O�+3�5jZ��<[�P��9:�|M�7K�@O�٩p�BP("�.���\�2�i�NS���x��u n3L��1���T�
+dnܳ+ǒ�����*A�i��M\D��]�F[�JPέX��XU���ʂ�� �w=����	|�C m�� �>��&��i�E4�12��y�z�-o�~�g~������&Z8@�f�s��b�*��1JTsǫ�F&���"W09�@��iϓ�6s�����E�[�Ww�q��U/�{�>��gI��mÿ/y�G���>�݊�p�{w�>�ʲ��'�	�]Ŋg&� ��r3\dr��C��lt��S������5&���:`'g�I-;�*��KyR?X��?m�hD�2m�����Ƙ0������-���-�~<6����t3�e���檇�ź�T�!�z�<sa�TTN����7��s����XwJ�Hcv-l)'�L�,x�WFz_����}���p�����j���J¨��O!�X���ێ����#�s����=w!J����� �w�U�ln��9�T.$�4}��R�0��43l��a�e&�^׫H�{�c1�tu�CIձ���R8u�)���?Ow���쇩�Z�;DY�)7�L%��ޚ	wS�|+��;}q��Z�|�rE&4^NMq_Y��#Uݰ�A�����Ǥ�"�}>Y��a�g�{͸ljG(fh���3)�W�`B �:T�$5���Yg�N��K�y;3��t�rFM�H-�C���պ��BB>LX��\?�����GHL���F�E��IuI��v�p�����E`�@*m�8Ǐ#�u�g�{�t��I��f��.�K)�0?�/^��,�_�O�/��V��W�c6�_:E�|�)��̓_�����@+>)ː�t��=��=���X�sx�1�A�����s��q��g>��۰��Ny�gf�v�L��O��d���,FP�>�W��1"�~�s?gTm�1������0�$��׾��I��t���"V��5*x����%�a4�pHb)���Q���	�>|��ᣖI�?fΆ��muV
�r&4uH�+x�35�&�Rh� �c�Y���������8*�q	@�=�$��6��Q���11��?���<��a}}���7ƛ�'i��Ht��mԧ���ɟ�׽�;��n_~�޹�UNEA�k��M�x��S �E�ĻZ5�I4�{[��:��}-i~�X޲d�wfv^������+Ma��[�$ߤ��Y�6�X*s�F�2&8rИ�1'~��Y���jQ�,8���<�hIV1�>_�������2�.M����Ğ�h��mi|Pzn�rɽ^Z[c�Gj���:g]�fI"z�4s�{i���3���G]�Ƥ����D6Z�]������{1T^/F۩r�X^�bLi�A�8q�$����k�o~�7��(�۝�/���<+����	��D�{�������>���;����X2��8�����Ni1'��6͔II�2�D~#Z4���*�#�_���U.�_�R���{��_�2���rh�~9�~i��l�Zک���*�P�gP�" �1cГ�s�3�D'Q���병5r��Ӎ����m)qҼMyV�h��Ju�#Iz,�D���(_�ܚ��{�M�Q^qu���7^g�y������sd�|�HhR%�@��������Ex���J�u�M)�3L���z@�r�����;����V8u�8�׵��c�Ke"G^�ʘ�2ru�Nr�.��Mv;��7�e���^�~�BHm\��㸘����l{s8?����~��-s����<+I�3U�i?�f]���Z�0�!�FB�(cb�'vͶH�a9��a�K�6�& �2a�>��~�춓d[��1?{9�1ۮ�Z�T�h�|'�ލ�X�Z�����ًDpF5^ "��q�9���iM}v#٩5,��w�m���.]��=�5���������(��+
��8`�
y��� ��_��ᱷ��2.]�
,�ק�RX�!�:��Z�'���Q��A�u^��4���XU��\��9Sz�
���l��R��y&&&�h�(����Կ��eHAZ�w���bgDz�5E���;�<�zGcoX��җ�|�%6LFR���п�����&�ԋ�*�}����3�t8��uwѣVι	 ��8���DǺ��E>M�4����(P�i��}�T�y����O_�KG.�� <��sp��U��ɖ��3熩\-��.�v���	��}���>}7љ�b)�f)3J؅N���c�.T�P���U�C���.��TH�(����L��[��A���-�Y5i���u8u��<y�=��ki�H��_»���S����#�\ZpF�o2�,��qN�t:�����㮃�����zD����h]����_�A����u��2�`����j�!OS����i�F�9k$1�J���9x�$�W�[;g�g�ݷ�����і�O�ީ���_� _�����\��t���x��I�Ƥ�p����w��;�叼�<�%8r��`۬7� ����>���Y�8r�Lj��+����Y仲�UX!�Y��w��V3鴣�c��r+EO�f�-s;�^���q[�J�"T֑Z����1
���[M�%�Ѭ|I��o���c�j�ߢi���%�l;=�������m�s7��9�����^u��y�E[W!".�������SC�:���}������S�-�K��f��KO�Ε�n����������uX8��W����W#i�g�E9��wIkAU�����J�>n{_x�R��s�-ְ���<��BT�ϷG}��}cc39z��]o�ԚW�{� �9'v+��0���G� %�y�r��Rw��Ù#�kfV�ǹh�fn4渮�֠nxQ�2�\�~�4���ܟ�ז��8�&w����>��2���s=lu ���â+�Nm#y�)Y1�tr�R|�������p����]:���0�t��e�|�����{౷�������D�m�8QO��Q�*K�׌�0��X#���)] p�B���9�-�B��\F��G�+WuT١�m �eny�Gn�s��&;��}�@��)W�F���_�*�K�ڪ�����#z�،��E��JN�ݴz���v��%%��ck�T1C�o�Y�Qa77�����B翕����5�hvr���:��u�k1��W���<x����������k�h�����3+�[?vl�\Y��-�w�����*x��avf6�5����Ř-L&À��Y��4�L>�d��eY���7o}�\�J��0s�W��}���O0P���~��F�3��n��ڻ^ZA����F0��� �>��]�[U0X��|���i�p꤆d*��ox7��PJr�׮�çؚu��P݌������UNn�u�nn�ս��Oћ���@���]�@.�X��
�ڞI��$~_�������f�~�_��[n�����&%���ڄ�n��C7��+  ���n0Gn�Г޻ t;<��	��
�7]�=_' �����=O�,�+��H��1��ի�@�<�z�j��ǩ��48(��Ӕ	�Y��F��ĥ���gt����W44����XEB!�Z	V��uE��"O�)lC�Tz�];;v�s��������@[�����\��X�Ν������ѥ��(��=`rcb1���w/��{���_���iXYZ���9�Q����.���Z��u�衍�)s�EP��xf���i�l���I�w�W�(���~���S�oN��R6L��:��P�p�}�R"���φ����E ��Vj=�N�&��o��I*���MO9��{�9���{�]����x��^1M~���*翈����*�o���/Go�t~�R.K��b1�w�������~}>���sgϒK#�u��A_],f\ ���l؏����/��{`i�*l�0mC�
A � ���˚PQc�"=�z�d^6��W�؍��Z����2$7�gd����'��'�PeD8�K�ߵ4^����������ufad@�}���k��X�%�Zϙ�]k��� 4���!ZKC267ΰ�7�E�_訛��r���b�����8����;��\�]&=7�\���I����%�4�Z�|!����l�zp��\��.:��¯��/Cwk.,0Lc�m��Y#���B�zN�)�KX&����mR����ч�G��Q9�j�������q�D�y͑S�"Ѩ�A�P�X_�g�ƅ�Nc�`�Wg��ya2J5P��U���쪴�g0�fǯ�h��y]�*Kv�s��9�T|	���^A����Yoٷi��i����^|�"w<v7����Ç��3����4>���0��1�(�"T�p�}_��u7=���wï��/C��Qu���)R��
������ �Y3Е�S���E���%86s
�/2����a.�oA���`�������0�<&b�s�@"�P����+��e�D�V�b���zw;�C+)�=2�`�Y���U:K$��Lr�C��>�'�����Y��P90{���9��]��-�S�ѭ��-R*�(t�4�'����E�6�����>�I��W�
��qX\Z�#��7��:�
��e���}�Q�g��'07;K4��)r]���YK�vz��Т�/�j�N�$+d�:��g	�C@YZ�}������2�?@n2��:rOMZ��k�k^J:FU�Ο?O�X��giޖ��@�Mjh�����΂[i��s���x-T�ٛ����;�}��E�T��!�rB]�����w�N��7�q��P�df83a*��Ȫ����-F�ւ�d�9B��ϝ{����#<��p��E:
9BtK�1�jDh_my�~u�����>�&���^X^Z���5d������u�W���}���Rv!K��� ���C\�b���y-}k�vn�ϣ���,F� ����,^[����_��W'�7�ƕ�)�Z�����ֹ��5vaT��z�E������\#_���K����ms+,:�;��7zf���m/���������67���$:?�e��+�����c�@�������������ǉCGjQ���@L��ɤJ������敷����O����Ǡ���3s�����5�&;����ys�l�"N��8ѱg¤d��i��r�ϘD�x�滭xe��5 ~��r�����8����H���ぃ�6��:׮��Q�^V�k��ܖ%'k�X{ˊ����5���f�i%�P�k+��S� ��"�/ct��X�:7os�X�P�N-u�����n�V�Nv���\������I8y�$�������Կ��G�~�� _A*ti�]� �9�_����{�G�.�s:��+G`�@�:��F��uJ�9׋K�q�^̢R�@��f�%�^̖��ϯ���
�Y����^�O��ә����D��� �E�+���H���n�0:Q����|�{p���K��q��K���R�\�f-�*���ν�x�c�����f��W��ժM�v�ƸڍnF�7ԩ#��1 �n����JL��/��P���ֿ�-��r��e�m��¼#�禈nl�C��3]���_�o~ �������p��GCiw�\X��3
>r����\;o�k��h>��9�Uje�-������f4%08��_�җ`��O��zn��o�Zզ�w5���Ggdº������.+j������x����ۋjf��^8Y�؜��+��ܛrê�a
��F�q�en��J�oG���N������,Y.kă��O>I\��?�1*�6==E��z�j.,��0�"5������.x��ԹەJ���Ӡi \�P�dެ�J�`�A�d�ge���nv�J3�3�E�T�ڬV��E�e�26�����s�yB|��s�]w�y�+搫�PՌFG)`�HF t"�9�<W{�r�� ���yQ]�of����{���\�K��2��)��| ;E�� �����>�M�=쯛x��o�1� e(ߦ'��K*@�.9����߆������?�
��
��eh��Y�^�may	����?{�,�u�	~�Y��y���6 � @�ЭHq��$R���"&b��ؿ���?V�i%5�J�V):Ђ@�a�0�@hﻟU����=��{3��ճ�\���W�����~��� �����`�����
\���t}T�f95Yn�����#�x��\~Վ�����ݶ��u���+þc�q�M��:Y�&S^.F���)&fg��|��GK�/�Nap�_@߱����ҀdC߹r�`��kYP��n#�[�{�9�i��95	�u[A�Rp�+��n��6��M�� ��E���Ys݇m�fh~Y^�{�����кݻ�ڍ� :C���n:pPnм�I��&ì��j��~��Vz\���q���{���e�M9&.W�������,-�+�7��7����@�1�6'ъ��s�3��Qq�K��"r=!c�Q�{��*�[�'8�Ҷ3����^�g�}�{��2[��t��%�8qBd�����:��X6d`i��ZL��|�z��MQj2�c��ʪXy4��L��v�|[|�W3��jU�ZK��+�I��b[D�1�xa��h�����n`u}��n�տ>3N�]q�y@O���Vm�d�eڱ�a�Q3��1{*;�X�s��'&'��sωD �3�b���H aV2^�-]J�5=��e|�ӏⓟxw�}7o��gNcӦ��uIM_^զ�j��qI<b0���VazpV���_�VP��ծ�\�֭��j�������Ç191��۶I�~&��s�kЅ_�>A/�M��W2�p�VK��(�=%��zIg���e7������w�P:|�|��_�ǺH�ܾ> �����뙅�dbD�W}���[R#2&��X��Tx�7+M鬎m���cŐ���S���ַ���u�Z����Ej	�R�.ҩf�+����?���W���M�h�e�8C,~LL&<.U�:U�ɱ�M�M�YB�N�n[�k[+����l~��Z�F�������֛����Y/�~���144$�s�)���
~q|�Y����R=�+4�������hG�emU�Vo#��^$a�ע�v��u�#�on�YS�/�Y���BY�mP��_�/5�xi_ۭsֻ�,i-ǻ�vx���:�GE �gr�/w~(�c����3�8y_1���������Xt��6����hm���@��c����&�n��_�|������3���N"ְ�j4	�YR�C�+���ф�E��nt^�y,��gGZ`:����}D��+ǩ6�k]�Z�Yj��.�y.W�/��0
��a�\����Z��3g�� ����w_�YQDPD�m��,|�I����r&	a$P7&s�n��dI.�D:�� Rv�$[�S�JZl%HVr�婶=�������bWע?��mS7;��Y�rv+���L��(LL\F~z^�)�#�Hg��8?7�X,�h�Щ�B�o��e�s�>����!^~�%L\���� J�r����I���]pnЮ������=���>r�}�A/P����z7��-W��4K�2��X��U~ux�fC:��D8����I�S�D����V0)!�+��c"�����nƶ�6k��&����'�mQM��`�1��\�*����ˇ��#������y����麵�J
��S�k�?����w:
��iy��j�	7�q�ڵ��Bʇ��*��o=��ǎ���3عk��ߏ͛���!V�p�dT�ZH�@�l�o|����~Wdʥ������(4*�z��%Xl�:��{w����O|�q"玪m�9 �@/� ��;�8Z�&ju����ˬ+���^�R]�R&�YI�z2��P�B'Z���.�Z���dݹ�Zy�f�^kcSL����_�~jkSL�:'3	����&�pblco�pr��p���R��־ڶ$A]t�v��y�Sa5m���3�"��Nm�b6��Bc�9���N�<����{z���+��"��{����~�a�>4}Ӊ'053���˿���}LML!ӛE�� �R��RY�Z�K�a�&���������?§���A�^K��W�'6���_��Ū�&�ȁ9�Y�ﶭ@ٷ�����v�iQ	T#�j���(a�R�s��RՌz�j�$$��`)�`6g���}.������.)�	Y��M�1��fҎ���_��d9�n����~7���z��d�+g�vl�!�p=ZW`�� ���+��7���{�uS�3�uC�$�0���19=EL�Ƒ������'���?�?��?��;�"���_���o��T*�\���qX���MU/bLM�Zt�������=����*>��GQ��n��x���D�K(�L`;oC��YK]�( ��>�z���h��VnA���훏�6��E^V?��˵��ű��Dm�k��[:��\��}'`��Bm���XWk���7��~��^r%��,�t��1G4�?r?��\���L\~�;�nX�w��f���5���k�	�ػ-u�w[�k�A�����IZ�����B�<wбX1+F&���VC�O�?yO>���`���DM�o�(vN�����h�{ʙ��5�w��d�z2	|����>��޶�4�6��y�8:��
�E]��MH��
k� �����3�4�u�ݚ��.+Y�t�Ί@�޴�jn���0G�x"�����ٳ�V*���1��{�~>���y{��W&'��1���l"">�����ڶ�b��������1���[�ײ����7��}e�X�V@n�>w�\gUD�&�������?�z�I�~s�o��ŹFl)!uK	���nL�,�����mY*s�qL����׾��[��w�DY�Xh���h2B=[�4F-["bS斈�Gx]�uٕ̽|� �&�y�~z'p�k�^~�6_����2˩H(QM����[�$Z?��9q�:GP�I
 q�m��/d��&nT�d���֡5aѧz%��d��2����s>hko"���� ���@���p��i����Y1o���2�ҙ^�.�lSzL%(q;Vj�733�q"�v,y~�0�tf
{�؁-G��;���'�tOb���Q�w4�0���W]�8�ݖRw����%��-�jMB�R��|P�Q;��������
�	X�l�YcB'���2ٹ��H�Yu��W�}s�u���l	�s*tD��Ô��|��ը>�+b�+��>i�;�u�W�1�(�����@F��:�j��܊�Z_7׬�쥋E�D`��,D�n��[��,aoł
1��,Me��
K�^ L���H�j���y���W���)�ܾ�7�b��>�������㮻����[�LgQ�_��S���;���a���:qy9Z-( w�k��|���	Ä�&6��kiQ(�:�Wf�h��uĄe��=z�[�#�#�-���|�a��dTRZ��Dݖ)�-����0U�\I^Sl]*&	@�j~�.a���&�0A�˗Wʬ�/��{�lP��C���y~�ܮW����_�M����;m��ء�|�(�ĉ��ٞ̂]O-wY�˳Zb�4ʀ��L@f-�8�С�qT+.N��(q퍺�Co�	�8*�r}}����P�5q��E���p#�c��g��f���M qXq:'=�$8��C$eP�fY��K�C�]��Iq�l���m$��b���KW��Yz,[oI���-[ę>;[�	-����mۯ�`�'�
�ÌҘ<c�h�@�u�u%�՜�WҼ2�q�M��!L�[}k[|��3�űЮM�|��1��yI߲y$V�ֱ����d�ks[Bž�K�U�H8�s2X�$dQ �� ���W�\���3�G��+�� 2�"�&01����ž~~��s��%l�k������%,s���8���h�8-��C�C�O�`tl�RͲ+q�M:o��%҇k͆�ڀ�+�$U:OUR�=0�,�Ͼ��8#mu��76�>������L��|D�Ǭ~l��A�T[	򗾓���a��q�6	^��d�v�wTOm-�[q��T[��F��ǈ��
��q�׮E����3C��E�l�Z�@�,,-TD�/-u�%�~b��<�D2Mɡ�H%{�s�e�h�:�_�c��h�b�j�ZVL�c��� ~�P�U�R�42���K�����q��K����<���8z���Y����H=��������^�ٻ/8�;v�$.Б���w�\�3�`���kt,�z�UYk��N@j�*���w�������3�\&�p\�E{(�>�U6O��<mfU�@O�S�"�#�:#?�U,5�W��$ �����V٦f��<%q4�5Q��vЎD���b�6��[t�zm��?w��tx X��Uk�ކ��D��ҥK"�
��������v�M�}Gl��t/��G1<��M�>uV���yE"`,�v�٥�4�R/�8�ɋ�/W+����If|�VپX.	�rh#~��[ʜb{*v9����V��b�A��Tp��A��ګ�����߇d<�1b��oۅ}{��Q�a� ��w�DJ&7�r�}kۢ�Q��53t���m��ϔ��x,�&r�o냙(�u���7q�W���������y�-S��,?�	7��-^�}S�Z�Z���.�0�P�ZMA/���]KO�aѠ��(���zS5a�v��B��>~�x+5�f�م#X���󘘘7�������XO���u��d2�1��'��0^<�2&'/�I�Jr�HS;N[��	�m��1*�-�z�&2����W�w��cŅ�1Gl����m=q-:W��2['�ظj���ΐ��:��-�bQ�s
P�.��H�|�&��)���W�J$12<L���D����d��ӍM>���ax?���1T��*������@�
�Y��R@�:�@'����6��8�.O\ƙ�gd·��> �*3�M(����u��L��#!�l�7W��aX����`�AD�e�]�e�
�b��jS����w:W��nug��j�н32�5�Su��&�X��1L��bs�})���z���$���æ��?���	�=�"~��O0=�'�OJ"�c�v���!�e9w(�F'�����"���3�r�}���|���g�w��{|�ߔxjs��Ch��8yU�IE��n�G�'�Yz�i��M,�Χi�Qn��]�Kv��"�^�����x��OaǶm�����W���勨�˰yU@�J��d�0�qg�yCo�4+?[l��a���!���+߿�P�7�����A����FC U�8*�Ǉ�q�B���J��'u���98�V ��I������?dفy�Z�%%�o`[Z+fٯ]9s�R�~��垄����E�m�VK^�y�,�c�K\)b�m��
�/���0a���b�Jyb�Y|���������k<��8��k8z�8�7O 1Ic*)�x�Ѿ���F�,�N��ڡ7��/`dd���/}�K�җ����9��7�.8-�x��s�)ĳ4�հe01�����H|�칍����r��w�38x������}�3裉�C @�o��#��tQ���D�c<��#�`)�B(�J�Q��sF/�漸��_��ٶ���Q:jrh/�͑�^�Sn�/��g\�q�o����ea�lΪ���$˸��ۏ�8"N�Ճ{���1��J�e���c�(��?�c#�V���Ⱦ��n`�� �1�(�bd����.��߄�ް+]!\�㺯 ,�O�q�tN?1tu�q(q�`o��ybf�V�1��נ�h�(2�U�c�U�?�h�il�я�^��{�Gؾ�N|��O�����v-<��3XX��;＆˗'16�A�7I�M@(s�k�Kő�s������?ǟ��?C�3�L,��y�=��C�Ҷm��``�"U�u�y4�BX;I���w�l-"�u�혣I䟾�=\����K/<�Z��4���4�YK"1~�ЛˊI�#mF�1::�x2���ؼy3vmߎ��ĉ���;�|��Ƥ	k�3�mp$R��i��+ӗ�÷V.Bj\eJBI#lQ����`kG�Z,��֋ŢT�z�g0;?���A\�x�?�n�}����G�OQ(Xy�v��y���=�)��-���[y�G�;4�-�F�ϭ�1Mָ������}k��ks�����-���q1М?����lkw0�`���ꯖ�M.����KjI�2YLN�?~�$���(�q<����2�D�x��?�k�@e�@��K"eh6�E�>�LoU�x�VSB�ԕ�A��}�:���N[��"�p�LTc*`l�N�C���NZ'AWV���S�/QmyHdr��9t^��Ҵ!�-VDN878D�ac� �:Sƙ��9�&�� F��\Ŧ0VKܴq�H��v�mȤ3��?M֤ҫW�3䨾I�dH��S��&��,sm�"�)p)g)�9u�@!�C�0��Wv�FM��*�
�[B�Q���Ӏ�jM.����՞�n��Ff�ݨf�����:��?�C��2-�َj��j�IJ���XSԚ�iK엶�NZ	$�v0�����o#��ţ�>�/����K_�]|�o�o��:��mW�=�	+��&��'�΢bB�u��*c拽�ρ?��(Bd	����2l-��/�(:�z��[�M���!�to�S�~4���Z>�dZ@�C-[�jV1)��q��RAd�k0���G�X���,��JH�lzZ�6.+�]�v�� ~�֭b����EP:��y�c����:�S��������Q����1����&]����7\j& s�m׺��ĳ���T77+���7��YF�b"�������x3�������*�sJI����Ù��$[��]���45�*��c&Y%f[�c'�#��y���ԏ�	/��<��!|�_�o~�k���~��_��%�t�	���z�)�'��q�%[M*�,Ó���d��uy^��>$+�.�� �+�*].�a�����݃z����\�#n�T0G��#W0O*
5	d+zBj�{��'!>SW9�O38�!�LI\8�8ۏM���Ǟ;�`��=���o�Xl�c����!��~7��� #�7�2�]�|IV�jg�Z�q�&��#9�66��=���mO D���g�r&��k�����6PG4>����4�}��-�-*���9�>�z��K/�CohhXۉ�z{�����j��ue���,DARk�F��@o���/̛ǲ��D�����Ϟǁ�-[�����n�[o�Nl�"��h6��]�lJ���f�^1�f"O$4S'?Iɶ� �6m����&�ʜH�a����n��d|y�_�4Q-W��f�|��D�(>~��[��@�J����K`�X5��m]���$۷T�,`#�L1gp��	<��_��kwuAf:����lظ�oߍ�6H�Yg�z�ú(Tyu�M>���j�	�Mw	P
���2�p������(VܔXz8r�Lƫ�}%�ȹ�}K�4d��a����m]m5L?j�ꦥ��;k�m�_�[�A�>m�C\���6ځ�1��Q��4���������/|�C�:O���"�Z�HRN*�T�F;Oe�~�K��<�U����KbT����R��1�̶ٲp�D	'����۰i�f$��	�Q.N�T8�
�-����J�XW'�H�@�̘[���2积���&u|������P0!slB����\��YG���\�8�]�P�b;+Y��5��p�]`�b�Fp7-�9i+Mq+ 4u��� �FE�Ă�KA�s���9;k�oێ��y�g�ΝR��'pG���8{��h�a@eg���XS�]ݾV��Ie�6r1	ee3��%�r���փ�H�Td�+�k��7�'�ڊ�z�f
[��Q,7�R\Y��g�B�\z� ��^�_��_�"��O}�Ӓ�π�۱�
𢡄/�C�:��-=*t�"c���ߖ2nH$��X�A�!S�I�N�}�fg6`td3��1:����l-е+�^V`d��+/Zʮni��Rta>P?9gmiia	K�M3x6����V���(9�bæ������U�&B�I���:bH]�L�,ok�O�-E��d6�q�}�.V��7�X��������Ӥ����|Ϝ=+��8�j���������޸q���ܖ��]�Bۺm^���1�Ӟ�s�f�<Yx�!����4�|o�1�hVh ��Y�y��H�e�6��v��iL�^]/8�h[-�.�R[���Zjl�پ�V�z�p[��5���iK��NG~2��Ecf�����i�<�g��%�����zO<� ����y��λ�-�g�>�#&v�𡀍ʵ���v|���u�QWU��`�����h���_S�VJ�q�8��'b��em	!�h(��kr�nK�ج#�r[��e����*��@3D@>4ۈ��~�j����)��%�ZZ�A��JI�VG�lOB+-��R��6$;�^�oq�چ��8�?K�wҲ":�Ɣ2v59����Dg�Uf$>�ɩ)q�3`9�M�6a|Æp�� f�Hy����L�N��(��M�����°f����r1��&A��h�w��m��	�o��i��a��Я�c�˵p9��˸9ڍ^]i�g��bi�i�	�
{r����@�}�m�������?Boo}�<���c߾���b�$�~e21!W�ݠ��m�0G�2�m�k�⨂���Lm���SE,qI��S�LP��c�K�H,��@OO���<7?�J�&�lW_bó�&�rj�G~j0gP���}]X�'S/��n�Z��V�,㩬)?"��c����u��8c	Ke�jۺ�
�^�w���UXm�H!mbቧ�3C��s��y<��r���ۋ�|�۴""F?8(`m�nL3L�$��`����fg�d��bUV|m5���f�4�mƝ�N�窏qo�fv.��m�J[�E�BΉ�.r�u����l�w��� ����F�c�!ڶWWpU,B�x�#6��~�;��?�^}�]��%�,�����S �Z�4xN�>M��EI�dB�`mR�#gR��4u �2��	�#W`*���W�Fl�:i��3咰7>�޾^T�U�=v��P��@�J��w�c��#�Ή?� �-��m�l�5�Yjٯm�t���,ʴ�`�a�V�n [V �r�BOƶc)�*˜_�]4� 7�m���pM��b{l�oʤ�&f�Gtm|��rI��?��3�9w�lMN�b=�l6��﹇�A��{������l��{�^��ٺm+�]8/�ɤ�˗.�$E�Z���ʄ��������T��#Bs�o9f�k�r��#&O��Bh�
�C�dJ��Ֆ���ۺ�JRޏ3�m~�y0��,d3�}z���O�o��u�p�"N��T���]w�:i{/.Bq��	LNN��O�����NШ.�Z��px%f���g?X!*�o�b�,��v*`#�ȦQ����R����b����Vm�`�*�e� �lf�%���D9\�UOKJN��5FL����!���u}1�('�>N$�L�������0�`�긟(騙�{�.+�-�9��|<��3�����lR9<��3�oܼ	9Z-�`�6�Y���v�@�|�$,�=sV� ;�p��3��ΰ��������݋�wbl|L�=]��\�m�������*���k�]�:�A]>���~3�u3vnK-���֮����X�S%����Y�k��?��?�q�����u���!F�(Z�1���Y��l�����11��ݳ�;��iAxV�l̤��%�b+?x�:�T�7=�̂SU�${�K�U0��;mހ`�idfC�,&�H�bPa�E��Gضkl͢W�+��/k�`�+ %���m߉�͗k�ތ��.-*�o�}D'V�LHQ�`��8c��FFdBਗ|a/_V�u�����=��ǎɝ�Z���j�?|�)Y	�������Q.�5�BpHH����S"�ā_�}���GŇ��G�`�$q�h%��\�@n��7������[�ȼ����#n���Vo�U��X�����Μ:����?�ɓ'11[BO�RE4\��A&�����2���9�����:���c�5��D� �8���6����"�����N�X<�G�x^���D���w|��SV{�6��߃���:y����b6R+qچ��6SA��u<��Y������Kǽ&:sLP����}}�lU�*J�Z�zЎb���i=w�f��]��l�����dRԏ���ER���㘙�ՙ�*Z+�H��طն/Q�R�a�xQ���3321��x��`ӆq��mt�t��Z�P�ӱ�:B��-��*޻�Z�6q�^��3!~����]����i�c	��8y��������#�Fc}-q��$R��[(c��Hr=O�	l< �9۔�)\?,��ÈM! ���k���D��'�,m�{��\���[�vZBO8�D�������z�ݛv�ʶ&��';8}a���[�s�b��=qY@_�]Ӥ\�4(�'q��)˰~%�f&�o��'�w��p"B�3SN�c�������yvډ+Q=l_j���Wf<�a��B�x�m�jR3簸2��C��c�z��d���/���S�#��s�ܹ/�FF�ټe����/�����M� ����H�Zm3=�F��M��~�]�����	G3�38������:^x�5�'-ԋe�%	�-�8qK�����}�a�歸p�<zh����"s��`g�.[�vO�b�a�
���y���K~f f����1�lD~����Rg��α�c|��F��ڑ�΁#bh�H@b�}��VǤ��J�Bzb�z�|�#%�|��mB�L�_�.��,T�CJ4"�ב&iL�7^Վ��f����ΊBa����d*J��{���`;ϵ�7=�S���'M�)�+yU+5�+��O~�W^:��_���ћˁ���UW�f�_{3��Zvb�ǲ�wڧ��W���xC�M�K�v�-��+�/]z���3�8z�	b߱8��4�>t�]b�OLa׮��2�s�S�pi{�	4�#K�U8�c�E�10Ř���Z+�CD�:rn�L�j�W���x@HL�1��1�&bV&AI+,m����6`�@Px��53�V�&�7l�l��Uٻd�}]�B�
'��Vfd������z�˙��M2�|�Xq��.���.�<��꫋��s�iE�ev(��E���w�cohX�4��̭h�rY���P��ѨU����bM��W������� �;��r�i��:��//���R�z\[��~�)���_E����
��J�����tU�.��]���l�����a�0���G�:�$-o[�
��9�$3����ƾA|��'1�٥��ݷ�NԈ�s�;���8yO=���P�su֛GB�|�8�pjl֦�:���b0�E3;�܊0ĕ�1��E�2�h�C�U$������H�Z�^����pD?`�*t�E����xJ�V4G��_eJ�Ǔ��
{�"L7�$�CS��Ơ5|L4��,��_@�۹f%FvN�a\��,���t�y5��(�2��M�Qg��ُ���f�v�\b�1���T2�2'1����?�{�o��<Z�G�n�;ܝ0�"�1�ٖ]]�԰�o4._q������A�"�Lajj/x�.��%j�RAo64ZH�<�t��`��voފ۶n#�˥�U����{�^8p ^|Q�!Kq
%���н.����:�G	.����PWw�X��#u0�`1����-����sXq�AUfq.k������!YV bbQSZ�!�F��j-9W�}�������� "[�����
}���a�fRXt��$iw��V�Q����ZFTk��������e�zJYY�%��>���'�kb�a��3x�h΢=~�^}�5����d͟�󖯥���=UXkn�v́�Ve�Ѷ�k���rL���\��%:q�8N�:�?���=��o���r��Q/�P+�!�3�^'��X�Z玝�(�t��djr�[~~������T�Ǚ2(`7Hi4^ �e���Dxh�/����_����]K��QT���BÄ��A��A]��6�p��f�-�m�$&1_X�~��|9���^��>:us_�>C�H�����k��e"�Vs��I�w��֋ (g��r}*��E�,�v�]CZUI�`��~&�;�V2�����'��8�J�ǹ��CO�����z��dt�nU�Z�o�˺q�ݮ�����0�q��ŋ�g�ŋ�zNb�����ʾ��w����9,��æ751��s��C�$��m@YJȩ$����ۦ�3Bf2*�l�ps��G�.r�:6d~��aϽJ-��P��:��{�X~�-U�/�����i���{l� Y�)%�&3d�&�
�Oe�����֦��:��ւ�i3����FW$˵��5�{t"�0OQa��C*j��E��:�t�������"._�p�r|�)�Y��A�L&T�\f�VL��DW	����۵ (׷����� ~���+m[��lo�����
�t
/��f��1�? ��J���`Bb�9���D����z�2�j��g��q��ILMN	�1z �0�L2fІI<L2��(���s����~S]Kt�׉��y��3��j��麯"��R��(7���LRA<��&�sѩ&�a���ֹ��Y�B�GM0�#$f�CV׳X�ކ����b@�|>� De.�H��t���䚭.L}�fj�b$��lW�����D������}�6���P�y�&��a=��N��5�խ����#+�@����oE�+߰׈E0���yzб�Y2�w���x������/|����B	�%�D��%�L���h���#g�rj���s� �7��M�t0�0K#2u���y+`�e��2[ȟ�އ>��|�N�^�c�M�v�q�*� �(�wIc�ʧ��~��լ]�G��,c�B�y��� �k�b�ϱ��s��C�E��Eh�6�w+���J�lf��Z�JtB��jO���ȵ�."tp#\Y9ф�.��}���w�����X��?��r�Ǐ��4�����捛�������A��h+� �`	��h7���Fظ�g��Rs�Q,���~�_=�,��&��[o�|_�UX�p��%�grHS�k"�^�)���� �lߎLo���;��.�6nt��*�b�4ՉB�V�H�Am�^
썍� �cGkS�K�k���w��6��F�_�R���Dh�-���*>I�LP_�jv�?�-~q[N�<
�V�����n_�ID����U6u��uhBa�s��E&���͛1=3��3�	>B���N�jEeA-"UcI�d6��=1'JZ��P9�}vfV
Ǵ�x���)���yodkK}���޻�����R�ލ[�ѰT��[�w���'�坸��g��;���$���o���*~�ӟJxX�G��ӗ'�sгi�s��K$02>�-;�#�JJ|�M�vNkz���6��:�K
aHX_?J�E�&�0�^�*K�F`��u����rm6Ո��*4�����Ab)-o�:��VIF* �ћ�E����XD�\FK��c�&gE�j��Q��WO���s������R]�_��e��Y���8mF'b�h�NzȭL+@���+B~�M��/��6�Bg���M����g�&~?�L��C%_|�eI�c�y�#֑Z���������z1o�b7a����=&�q	9�h[k��z/�f����}���]FƮ�K��a<��#طg~���azbR"O〤�pj��t�Y�1I,�EtÖͰ��WX��>?y��,Y��#�Uq�O��c�	@6b`<��(�  �*?���]b�]����9W��s�����c��h	[D_V���b�BX��%�'6�jz*J�S�S��؈�
���:O���m�S�v:I�I4ZqX���:�����Ȏ�K�.)��ց�6�?twG�ѹ�ڗu����^�D�B鿰<?�Ç���߁'����;XaZ�rh�y�z������������%��zM02��?p����q��i��?�S��?D�� ��:-G��*���#Ig��E��aq�������1T�&��2Ш��[o��7�yU���[��Q��X�ZR 4'���-]pY�%�R1���PgFߵ�ޅ@�%-
t�6h[�9˶F��#���!�ī1�l:��5�F���~��7���O�Y3�������K���E���?r�7K�^�uKls�{J@�uا�?�8��b��l���X������w��D�o7{�oL@x�$	=�`�5�q&3��j<IW�x�w��{�ņ��y�^;WJ�j[c������VK5��;'KY١)��@`����H<x�����<�..���<|�c����v���?%�2�F}�߶����t����c�N��%|��[��� "���1��_�Dn�*N\�Va�&zG1#G������Kp��*}���5>_ay&�D����)Ɠ�
���$���q��p�EJʸ�6-W�9>�#�2�*�pD"Fb�me�Q�(\c��o`���OSPc-�xm��Z8uڵ�;v:����t�*'&7X�kph���lE�UV��t��˾�2����``7�BL��b�2�MV��<�J�����L���x����/��zn06��Q}뢈j�f�Ɓg�zM,W��.�^nlΨ��P�8=���~㳟�_�:�R~�1?1��-󓓈	~z�"`߾�DU�!�)b�SS�� �f(��Hai�Z� ��#`�mܪ���g;:�ۤ�;z�j&{R�P�_d�
����W�����r>��WfZ��y�Ƴ�-E�>gF.�28$�d.���i�#��/VD,��}�LȐ�Bؽ�'�6]���k*s�Bxb��\�TE�p�)����o[�\m���n�sA����Q�`*E;��g�� �w�\��ɫ��W��Xh�A����M����sV���1ϫ%+�s}~���b8D��M���}� |�ay��SIĜ�n���	�z�M�^n�n�NΣ��爱�?}
���g�c��֗��������(�8:�v�8��|��C�6��e�� �G�:�la^"c�{�H��"�d�JR�����cۼ�@�P�$*��X�0.�ؤd^M4�oK|5�$����d�7Q����"�gs_k7a�ݚ����	LrD��f9�&*\�ma���*�.ד���8��M3�R���Sd��>>_�{^S��&�Onѵ6��I%u�TG&k^=ٞV���:*���M[G��q�א�DA=0%i�	��V6�T^��l�|^V<��s]����ͫ��C�����I,�ΨN}0�Y0�?R����W���"+J��W��C�~��	�w�]�'SJ.B�t~B�}{? �U���^�E٪ԕ;�;�VÃ�K�q��N��_�=���3��>��쉣 ��{���n�D~V_�L/��"~��_�v���a�ܹy�1EpY���y�
�|=�3�`*�z�˶����t��%����8*mߋ���2LV;2Ŕ���s��vKB0�I���MR�������{ħ�sIH���@��=��Y���c�j~3���<j�"}��0��`u�>�I���_��ۼ��t��(���^�:��EE��·�K��I'��f��PP֘��ұ,�����ფ�.m9@��πz�<T۵s'���T�'�w�y[���{{�y�f���̴�R�w߽�1�۟A��c�)�}a�e�q��C-���{���XHd���w69t��2�<rD�T\Ml�V��"�t�v:��J�J�	����c�f�Z�}?dh��:=����ݯ}�>����_����q��cx��������D�X�8�x�>T��7	 �n穋��;G�G�������g?�Y��42<�J��ݻ��#o����\�a��B����VKZюUp��+�25���W��a�J�O�ϲ�1���Qi�&a�C�,_9[���M���k{�^��1tp���+ч	���z=k��}֤߹^i���J�1�a�t�Xx�Z����!i�l��h�����H׉V�Y���$�uL ����VINCX�$��p�݈������\�gԪu����d�J$�#�g�:�aOP?���LTתg0�V��߇m۷�*�����_�KZ��I���ⷠgs��A���,Q��h��.h-ϛ�/o���'&F��oA ]��IƜh�"2&̕'�Z�J}�]����x���TF��|EXA�ڮ�[k�WۮW�Vg��򌽔�A���c�{�J[���j�_��Q$�D���_3b�Ȭ���jpU�"�R���6u�\O������ٳ�M�^.f��0Q�b����B����MD2�Ck(�<� ��g124$r����D/�4�Y%�o��Z]O�c����&��~� WL�"<Q8��JK���۾Y���C
�mQ�T��em��6t�6�1�3�$$�x��O<�(��$�{�S�L���{r}ط{��l��2�b���ݒl\UN.����#��o���e��SYZe�d��7Gz��&c(Ub�N�I�"%be�B��۵!�a������`Q߼f���(&f��h��i�������@�xV~��zD��W�v[h�q��[Bض>:2B�ϣN�0��;��A��^z�e�Kc�j0�QIp&
F��x�>"];W�\U����8��a<���2��tW��5`��un�&�u�r�v���S+9Q��:n�wkWr.&u�}n��ς�:�H�5D�m�\@�2��Ǳ����.<����a�R�S�C��@�XP�KO� ��A���;Lq��<-SӘ���I�}ڍ��7��sH1[*�1�:����b�h�.�A�J`G�7?;�J*��J@\����4�:�)ĉy�/�D���w��Y�Xt����p�G.��"gP�뷡�=�QlmCg ���n|/鼚�.�M�}����R���@�12�nߺc��8t�%�&Ш.�'�'�=��k_(J(]/1�;o߄�����>6�� �6��GW���+� e�u�ʮk5� t��I��%.@�[7��[��qF�����7��$��NlZa-כ���`�	<X�XfB��-f��6n�eM�#zp` �}��RH�m��¹Hz:��
IR����l�����@e�r�$�~�}�	���ϟV��t���k�xDsH'Y�X(���Ǯ�.�JH���o��������?%�G���k5�K���C�jW5*f5��T[jr�;�������;����o��/��z�@"�߇&kwp��C̰��=�܇O�sr��˗���,���e�9T�4��-��%�9f��+;��8eb`C�Y	�,�gd e��w4�2��i5P�'��B[Lh�48�1.:'qw��x�&�x
�� Ҵm��랻�<���2A�J�@��$O9�-�`e���v�>;|�������i�N"-�i5��fݧ'�x�<x^{��D]�L+����z%��f����ڊ�So�?�c(�`0c#��90�3�s��L�/�����Qr�K6�����4�G�	���J����3=��iB��C&���8!c7�E~;P��@�K���H�Y�o��3��R���������	%����;vc�ؘT?b�9������ٳb�B:��1u���{��? �$I/�
M�{���믿�s�/�*���S]k�[&qL@���T0�f�+��e"8���*��Z);;V��M��#�M+����;�w�l�[cg�*�F��L;�1�»xy��7�ʏ�F����cp��o�H@��8*ul۶��?��)6��-ci̗�8?_�D���䝣�?�t�@ߩ��-��Ո��N �l�Q'fˌ��8�?����~�औ&\���vy:��dO/���Ϻk�95зa��G�r	s�H�֥���du�q5�O����	9����>�PE�$"z.4�i�����ϣH��́W�I�y.M;��8u�-�<����M"M����"����{�#K��8:B�'vi�غi����#���Xm���ѹ�si`YB���`^Mg���!���5�K��s��*Qȸ����'�5]�ֺ�V��P�9��|Ա�t+������qt����XJ`a� �lZ���_<Ϋ��$(�q��b
c�];0C�͈��� ��2}ƓS�;d`��?���̩Sg�[�0ԍ)DDD]c�rU�C��.!�*�{M����Ç�;��6~�_�fZm�_�Z1נu��V7�����~�8q������Ҡ�F�'��	��s�w�V�ݻ�|	��A�΅IL�]���!�.�(��еؙ�)��z�#P���C�jUp�MhkZb��R9�P���p�e�hY��jvpX�ɬ�$u�b�q�Z�:���-n��NqAV$<Y�xFav^�B��i4JE4	P,�vt����\��K����Ƿ�(��v���N������ݯ���a��1O��$��i�B3ݓ��8v��!�o܆��݅��(���h�9�,ULѶt�t��0+��9�8��^Z���H%�`]�$��^�ސ�����_������Zb���)�@/�ظ��@���mJF��:~��ۺKl�!��'���-[$!�MK33E�>}JL)�0�y ����t� �y�G����cӦMj��c����I._X��o�m��k�+NL�]T\���r��|�k�	�ۑ#G���З�"����خy���f��o����NR�ze��P?����o���h��^$i�[i�$Z&G,��RvL�H`w���yb�S�3\&�R��X�BC}ܘ9_�xv���}�#���ۯ��co�!���t�挰#vr5���Q�J��фO�^���8�9M�A
�93F����A۠%x��,�9d�V� �c\ZB7i�^��v�G���_(���B�ѭW�Vo��q�7-4�����j%A�����u�o��ՕI#�!�����T���ۀZ��N�pz���o_@��kH�*ņ�����!7\�g��H����琬�%�f�m󸤴sa�Ι�3�ct�m�ሢ�n�d�����+�Yq��Taٯ��Jy��M��?,'�����`�Vz{{��r������������s�~�8}�p95A����LV��츰� 2��T�ɚ���d��O�=��15��8d�amS��-]4CA�$+�:�J�Cq���Q���+$v�҄�юm�n�_�`�ն+�%��&fG��m��QW�HJ`��!Ohsi��>�$�w����g�~8}(��T%���۱i�d��*�t�)b�ǧ�q��D��W�AS��>����I��	��m�g�O<����/bW��\|�b�~C%6����D�C����P�ruN\� mM���S<A�>�Q6[o+��UG�nE���A��x/MZ���z���x��>�ج�ha�Y'`���9�%.�AǮ�����25�"���C�̬!%��fásv�ݺq��	���x����9�S3p2è�x��M�=�H�j&�*���#v��tc�,�I�������\o?m���S��,ZUI�$���[oJ��'L��Ō��(-wq�Q��9&,*�8 A|�!OV��c����~&�)�d��/OL����O��M�p���uo�$M��78�N�lK����9��T&C�˼�8���/a���Z
r���Ae�ʶ��X�5A��G��F���E}�ϛW�{�����JBX��V������]�)�b�����ծ<l[��V��lܽ��hx=�q��t=q�"��s��2�C�4p�h��(��875��jY������r���sNv�L���#b�@}f�*�iq���������:&�I-�NK'��,���:���$��z�Ҵ��Y.u��I����l���_��L 1b�����c�&���Aɴ���9�����q��8��u�l��[)���A����m{��1*�MP>���=u��_\x咇��31����O$��ѽf�ڰ �6MZ��b:p��9Ic��r1��>��nC£]s"9�[6`br��519UC�&'�$\InR)�ܢ}�Ӛ���oK�A���՗��7BY��8O�D���ssy	st�0�,�Rs>Gsqx'O
�.�B_��0���_��Μ>�K�.��'���m��J���R��)C�O��\a����zG.��v�����ʹM�8��W�s�lܰ���nƫ�|�P���VC�-Xˀ������i�svj��V�%qb.�{U�Qb�C�͍��34�"�R��3�Ă.O�T��yB�RL������H���r�-�F�A쫄Ça��(汑����g��@+4��(�����]c�M"��-��|̢�݀#�)�7��$����"\�P%�^����-�6��6oކD*��oc����U�|�e���,�h�$3��i8�@�]S��SL.)ք�9��]�*1���,�'�Q(װc�C�K(�;eS��&��؁K��3<�+�y[4Y5+8tϽ�8.^,�|�Pf9����h"��h�">D�7�����H������C*a*=)��D	b�-G���f��-*Ƅ+Bo�R�фm�=,��)�e*��jS�T���� >O�&'t-�R�H@d����XꂳX4�r�^�;��	�r�Ǭ�����*���3�#�$$Z��Ͼ�z�D O|�R&:�������=vgΜ� ^5�m�cu(�Vp_��71K�ڭ���ux6���N�n�3��:1�*�n	$n۽o�s�[��%�~� w�Xƻ�.��>K�7O��+����* %l�����D����O Y��'?r/R�3Ξ:A�X��"�z�61��	�b��Ub�IT�b��9b���%O�
�1��'B�P��G��.�G�������F������هw�CӉ����
�	+ɨA�!���K�
�5xEB̍���:��B��z�Gbx3�ns%?K�D`Ԥ%;3�:���-�A�����j���s#	D��Z�2L�d6;YB9O��P�p6���i�=O�D�mݿ���ߴI7'^�YSz�&m�S�wΚU�a���	�P�ma�*OLb���pv�����e� �p\h�V�q���8K�jP��
Jֱ)�#l�lc�3O�M+0��D�3V9ҩF�0;��WX��F68:�;w�W&������^��K�����tRUUD�Qr%Zy�q�l޴Q��%�n�f��r{���Wj��Ր�]o�~N�n�f{����������2s��/�Rq�J�@ǳcHe{013��K�:w�>�07��&pi��f�l��Qp����|I���
(p&%K�8st0�"��%Z��8=���v!Ml�R���ɓX���ӓC��(�$6��ѓ��O��vN�$'�JW[��hB���>��G�ΟQ�Ύ^Z�M��t�u[rHo�,�1l�Ӎ�J:~ f�8/��6�җ�G�i��?���]�V 4-"�:3t����b��H���9ƚ�-Z�%�:��TR ���b�idF�$�բ��~�v��V�9�pzf��h����n�� �{���;]�Fia^����9���7�p�y���Nؔ�-��Uz�"�e��j����G�~��wS�m|�X��)�Q���&��2�plH��V�%��ǀ)#(��b+�%���z�ɂWc�\�a\���> �_��P�ņ��0N�IG�Q?�V�h6��4�4�2k�I�m4ŉz�=wKd��Fu��٬5B�j7_�Aj�u�+��*� @�Eg�Ц	�ԣ{^��%?���R�����'��(+�'&>40L�o���sؼg/rc���855'��+�2]wC�ǩs�jG��b�FDV���2YX�4F7�s,LJx���gp���#�)�j�|P���=99�?� �z��k.f*-L����F�T�[��Y�3�&�S�A4Wb��G��mx���A�b^�t�8Q4q9¢9��$��	/�i5m��P�a��(���IZ�Ч�Z5�Zbb�	_�-�*���b�E��3m+�w�&ѱ�ۑ�/gZ4s�qK�3lfr���4��5o�)�ap�WG_���搦kK�ҫ��G�����.q7%r�'���k�g�r)D_�hs��a�êu�<�X�H����=���A;��M��a-9<#y������^�Y���)p�K^��kuD`�6��8���y�?=��?������*��ma|x�vn=O�t��єL�_~C�C�{�F��E��{�ƾ�p��Y`=�n-�W`б���o۞/I9��I��V�E�P��-;pyr�<�M�>��
N�p._BŊ�fǉ��-W��A��tu$�4�q�}�ƒ(x���އ��%z/!��,p��%�v�XfO3��O�>��-�0<2��Y�g1�������HD�D����i:�Fq�=Y�q+2J��Y���g��>�AE�}Sl�D�hψGg"Fc����8o�m�CG��b9�T�BI����9х�f`�q��**ҢGʀ#|����m����{B҄�A2�g���@φm��T.p'�$M�=5��YX��Kǩ��f���(�bA�?�?��~8G�}5b��8�y��jWR�yڒIN.�(�+�n��� �x��1M*�U����f�E&	? ���<KX��Q���k��e�GQ}{W�i]���d[�����nt�}S����_�8�R��Ju
�dVX�+"m\*�����1�����xgN���3��o�>�_�����׽^vZ&6�d���Z��?��G��[\���y�d���m��˓��X�/N�<��?�-��64�^aܳB}�R��ۢh���aj��+���>�$m��,�}�~���8}��g1::�vhy��������h	d����AUuhB`&���� ��r��bI"Y���ąF���v�]�	F�\51M1���"TW5`�k$V�UϓK�X�^8��[bc�����JF���u:w�q�RI�8I��h�2�v�x����^d�����M�lM���i�B �~
�\{�¬�r���NO!?7/��b��z���w!�T���[�&$vh�~����J&ۧi׉�A�l%���=nJ��6mu�jr0բ������|	3b#���8y�N/�F�W��h�`��	���L.J��u�b-�%wMAqӗSI���e�o�E�=�z~2A㥌��id�,�L��5$���lN������D��m�ؕ�[��[�4ܕ���[z�p�i++����y$g��s�!�����Ŷ����er� 6{�m��6�:�� ʕ*��6�}� F�X�<ok��қY���ٜ[�#�\v�rlv"��:q�Rn�7 �I��q�&�/��(�[b�Odzp��&L�˸0W���<ʈK�����&_,G;�'�ۼ�yNH��p�	�Iр��F�o�Jl}@����PWh�d}��'k���F����`�4��s|9;��tn���8BR9�9�})�I;�_��#f.ȋ',v���Gl�ʧ!&Զ-�J�XU�CpOJ>���c�i��sP�����*o�����&���Y�9xz�����1|z�����d�r�>������#Cs&)�>c��lVD�KT�*�m�R=��-��Pz���J��&۱���Y��>S���>�Y/�UqtD镁����z"�l�{oF�Ҿ��<̷�Ak���.��b�����+MU�ʒ��._�$����@�p�N#�*��$c��t�{�o��[�9��C��{���v��>�O�Y���W"jY�z�r 'X�r�����b�4�����C��&\�����E������L�C,�ۣ��>�%fU�� � ���S��l�b�� �n݁���T��z��,zGQ&v��9L�83Il~�b�I:�&�Q.���#,�λě��W��`[�C��a3�;��;1��v,$h��|6������G���n����WK���,Ҧ/�M\������79����
�<K����q�tJjӲ�o�V,��<[;�%9˕����:��lQ�Lr�g�`|Q�dV��2��b��E
Y�3�w���^�i�`��$�!�3�d)>Y�mR\�������nۍ
oOKh�Z�� �f~C���lc�
�꒸�s�<q�۶�0�Y�����þ]�D�#}|C�¸�@��<�`��$P����--�k��J�U~���)��0�2H"�ѝ�I�A����%���148xq,���eN7mf�8�m��+�eM1���r��W�]�oE8�<��`{�_��%����%�\F�9�֓$K@��H�Ǚ�3��`��_z�5$����,���W��j�[��L(j"��|z��8,�d��\N���s�tmV�ɊZ�G>�(Ν?�B�L���{�m�b�TCbd͞^��,�D;&z4q�+���1�=�|���i`fjR2{i_)b�c㨦2�։QK��\	�#�V�SK?;����Nc�2zު� ��6nԈ�
��2�d�If�+R!�y��_*���A���	�Uk����[�)H�M~�\8���+���r1��Oc����Ȑ ���M2q7�uC����f	�*�.b���9۳Qg+3n�@�S�Ź�V��|ptL�w��
�@�]��%5M߫N\B�&�X��Ha�Z����vUA�����4�EH��<�ͭ����~�����'��HK�����(Y�~�Ẇ�+��e��뫕���@�y��V��LY��4}ΙϬ&����,g�v�K���:�z��0�6`Wi�ު3ע�My�V����������]���Ea4b���B[\�Bi�5Ɗl����7h�5ꪸwT#MZ&�>[(a��d
~*!�!���j{�H��^��%�UD�\l�P�ۉsi1f�q)��Ӭ�U��>\�����=,A۬apxPjY�,����c��xȻ�����!\�UE�u�i��<�H!Gt�����N�3��6}4�羇���C��'�Kp�Q�V%.݊��Li%���?w��$Yz]�����,﫺���L��`0 薤DrWڥB�E?*B��A��B������ƒ�C什����&��������2�j��c0��oP����g���s�=��>��L3����@g֤�@1C@�l�r/Ϳ�������6�j��3�H;[,��Eі��q��������A)�X`�Ϛ��8?��~y��W�c��=4�� �Zˤ�w�"ܧ������8�D�v�>��{���")�;�n*�(+�a)�,hhqT�	O�u���{��n���Y���K�LLȽ�,�=z�������/5G��0Q��� M�nh�q^=H�K�$����F�M��>�6��GXxU;ᘿk��0�u�f(�`s��T�u��p&�1Q��LL��p�O`���s��k��i�͚�����_�L'������8�����7��P7�,,߆��M��/ZCw��]yv�@?�1ykU����=�m1���-�(Ӝz��T�J
B�dRڱK��և"=2���^2�K#�C/���������1eM[�bZ���d�x#j�؝�A:+F�pA��[wWĐ!+�6&�����IT�:j"6��|������O⾼OS�.���$�&M��=$����{'�\"$���"�n��i�~��3��?���R3'3F@�n�߉�;��j��՟S�U���E4�~�\Qlͳ,�@s����d(æ�!l�D��5�JR����_��^�9�������(��\[ǻ7n��}��\A|����*�������"+�X���N&�(�3(dS���������-A��;r��fuE�9�T�37?���9�e#5AY��D{	�t��^�N��r^�Fb�Ym=?�#
�B�k:�ֱ�9'׳�q�R	�����Hп�J^��I�듗�7b�\"�Hd�6t5�s�A��:w�/�Iե��ȳ�>�:�rC?���>>eK?�#�26��yy�}��Y*�������U>Ǭ��v��ؿXT �(�@i�������L�*'OY�9Ǣ��)���h�0�m�%0�gkS���U��nl6%Do�5�6w�\F�b>�����M\9{A�enb.VyǤ�OZޚ��H�װ�V��C�h�]�
?���D��Q]K~�zNGj������#ݭC���ʵ���=q&QA�yL��U΀_�tQA�1'��(âAgA��C�M'��1�ֱ�*�|Iq,�F�?T��gc��_18���W�k����a��v����FEa;��Pe�d��=M��0E��V�S^kA�_K��`�	� �]W;\��G�~	�݇�̨5 Ͷ2����:}�D@��-$HT���F��`ji��H#�@�6qu���=�wgZI��׃�]l�`zn��y4���3�b+��i�NG�����]�N�rLA�ΐ���F}�5���5'�ώ��ˡ��~I1�r���He��+�V"��v=�U�훴�!��oXG���T�1��oѻys��}�z��wkk?�яt(���4~Ӈkk2��8+w�z�SZ�ֿz��7�qn�2��0����D�>�}-AXDe�&
c6�>⚫��!�n�Yװ"�El$N�Z�ET���6~�H8U�/2�h� �^ϴN�lO�t��bI
MM�j�%�vr4���L��l�fiO�mձ4+��9�)alzť%�q��";�߰�6"4F��zrޛ!��E{oS��!"͆�OG9)t�6���ۂ �#19Ǯ���F���8 ����!g���U�k��;���u�9)��M�jP�l*��}6��}��F�n, F[��pH��ϟƀ��S~���7��*Zotr�yp�g}� j�mBE�b���Q�ނ/H���"ε���Ɉ��^������&���;����t1�*L��5���u��g�,��|�T����GF"��8����	�!yV�6��
�P�HOML*׿|t�4���6̵9���W(�1���enEy���hhj�������5�~ȓ�0���I���<b��>��_ SO�ݹQM�9�<8����|D��A����*�&ρ����<����/��/�A����b�c���$W�:Q'h�݄ι�D�V�� �xRPr�9M�����d�dR��1��3�(��gH��LSTO�Nv�j����ȩ4��Qd��l���Ç�:w��I�RMu����@��w���#P�n苭���.2s�H����Lt8������}��=޼loPgV썜���k
f��%�Y�;\j��÷~����[>��s��\XDJ���+7��0�e��Bm�ǆՇ�`����uc������1vƉ'7���Ƈu��I��Utn�/�iLY<-�i��S1Fp�D�E����!UP���/a��b=��i8[�<�sD�N�bW����܇�De�|��V-�P^$��+��D6�����/<�?����8޿�'�zX�Z=��F�f]�$�.]Y���֮��^O>���e4��;���8J��D���o�����l�BQ�uw���-_�`gC����ݽ=�HDP9��4�9\m�cJ�r4���v<�z�t���Ƭ�%�+�4�C?��dsz�9$�F}��#����y��aę���9q,�=��D#��v:m�[��!%8j�-���X\\R��U(����e����mD�G��T�}(q���<�כ򺙂q�e��8�_&-c&�����[�@��L3Eٟe�/7�v�'��W*�T��L��e�aW�YIml+��jc�����O�k��>��)V�M��g
t,���qs�+b��e7K� H��}[��j���V�.�>�Fr�9���ݻs����:��:�ri�dU�F%����n�b�C�粹��@UII6�^��o--�A}"|�� �������¾e������X�)���aq7��Q�`�\��O?�ph�c�F������������h�_��D57��N���C��||g���X޷����s�����?�֎<���ų���l	�ψ�=}s��D$�E�L��蓢H�z��iYgq|x�.�7j;ZQw��|<�m�ŬP����m��8��"��wx����Z��ZE�A��%b��˧�p��K���!(�3�xJ���&E�h�ym�kk������ÿ#DY�V������")��C��	��j�%B��Iu�"�y�|n,��e��e$r����ĩ�b(��r2��1�p�S\ޟ|~�JS���G�DBGr~��up,ߝ;w���Q1���}7l}����;�s8����{��z���"}#�qE�4�\�v���+Y	#t�����|5il~u���j3�M��O��"��mD�?e�j�;j�C=�l:#N!�݃�޼���U���V�D��T��ەp]6�i��' !7�����Q�̅�r=I��=ٸ�v"�_������L��c)���-��<�)�N��L��w�:�"��`c�3�McQ�]��k�L�1̰�u��'3���м;�c��aR*�M�|�����1Do�a�FQ�R ��v�g�Ӣr�X�]{�z�w°��#�d*�ŧ���w_�N֮WLu�p�"�|�E�:Q']i֘i� 0�d ����W���<񄼮V����jQ�������(�Q�Y�XY�F����� �-t+S����(�;�H���EM��LOabb\��a�b"�^G����<��R�}��".�;��Z�-�=x�J�)΄���QE�N27�A<[T5PGzZ�h &M���ly1�k��ZS�YX@�ZS�M�^CC�{G�ʾ��۷����­|f^E>aRDL�ii�@� ;N9���B��{H>��#<��3���U>�K����\_u��7ⰱ�3��u�*�b�ЈG��Ͱ0�i1EA��k>��!zM$�q͍v{�ȣ����{�L#�ѧ;�g�|z^rC6PC67ez^��]7��-���n�_���L/�������ɣ
^T�BO~7F�(P�#����z��[�j�sf�k�0q4��y�����((=�� �����9:������8@��nh�\M���ק#�Ke�޾��g�r�)5 Z�R�w�p�5�Y��e�I���%��7z-ᡯ,x2��m���yȈ���CZ���涎n�Qlz�n_yб�5:1J~#AU�� g�n�Ēs��z�|:���fCх�X��A�����bT9k^{JsKZ�\�˱nr~q1Jc��wK(l"g�b����ZS�be���Horjc��ĕ����7���?`Cp�z�J��[�!/k�'~|r�>�4ff���NK}J0mA�ˋ"�����q��u�<x��lx�:ڎUP�VRY�
c�$r�����1xK���y=��8A��c�:�޶|&D2�C�"x�)g�.d�z;uXB��9�6�hc5qR��q �~�8��(uw�*eT�emh�V<ߟ)N��G�s�mg�A�#���ݶ�܆������;_�&�Y����������c5.,��_,�X�5)��b܍Ű���c��U��)�G]+�Y�J]��L�0=hg<�����=�-����8Z�(�-�!���#+)3>k���C�T:@�TLY9to�v���`Z9 ]O6��U9�k���(��o�����,z��-DF;RkQe���i�����޳�w��ɼq �˫��PPV[��dΤ'�1�	$�ͱ3�N�v)ZBħF
�������r�}S>�}뺊:Y�8�H����P��	G8�tV���8ؘՊyT�w<u�h�?����@���N?�4��h�R����b>�j2�j���zK�n��),����n�0���%��*b�V��� c��M\8sF�t� ����[ĥ����/Wiw�z7u�mo�W�t�lJ�󎬯۷n��g�#����A)��T$F:\�{�������7���o蟛�~�?x��CN��NB����	,�=�� � ������(�@ ��h
����eu����>�}4�''��<��e��=35�%��5(o���7^Gus���0#�="�n�3e|2�TdL�<h�e����ߪN<ׅ�{�sw�ӗ8��QN#>����[����bN�ݿh�7u��38+�rq�ЗA�!W=LÐ�5蝃�cQ��(=���FY)^�'!}D�yw��z��w5ޔVUeCg���# {��E&Sl2���E(��˂����[ﾧT�f/�ȟH��s��aleC�:�&@���'1��u�ɱt��쳔'�jq�W�9%A@^�&��$_� �FVu8`rа��аSpJ�UX�-�$bbd�x�(&���p�������鏁����(-,�������C��?>e�O�G��c�R<e�:',غ�J���+����VL_�^��O�0cA.��s���G���ol��w<[�]��V���/.�(�Tְt�h�xqMN��9�۪�.O()���T7f|3s�Xþ���[�����
�5�.>��D~�* 7F���@kY=�!痺݆��''�U�%�n5�Z����Ge1�x�����kJ��?�������f�׏
R��ըs����s�:��.]FT֟#��t�(�ժ֚�#в7�҉Zdoq��~zĲc�a��T��Lq�x����\�������~I]F�VȠa���P��#mֵ��F%���!c��^o_�m��1?�rF�ǿ��9�c��\�O������Yc��u5LWz��vJ�və
�~a���e)J��Z�E��1�g�q3@���Dr��2`N=�3.a,?��w?���˩�qtx�ܒ�,Θ$��Ȃ�f3Ұ(e)|ȍ�aO�O#.�X�|m���n�-��ނ�lJ�]� ���Qx�L1��R(ǻ��^if�&�������P1����[7o`���Ĩoɿ�5BPF��]��h��{�;�~ ��Y	Gצ��=�x"��قi��0⋆��-�G�Яp@�mO�9(/[l<��'?�1g�1��,�� #f���uЖyu�e\æ
�~�<&N#���~�#)�$�i4���S�>�q~�n	`�pg{K�����ӗ�p��Osu����˯�6|YS�jI�엟xBg��u@r�k��)���Z?����ʚ�gd��tb�DV�rR;�9�`������=wdy1�=�PA�r�;;ۨ�o�� ���F�����SH��!.QH�u׊
;�1��,�nόx��Y��O垍
�(�g�%������y���s�����-������ɘ�'�S��/Jj+�o�����u���5������x�Q�c�.���u����J>��-+YB����O"v�N��4<� �g��y�wqa���,

]E�Z]�w���	ə�g�x��wq��M/j���D!P�]�cTd+*�=?3��˯�U�J��T�Xx�,����H'u@�6�F4)�*h�Y���<�vj�g�ZaRS4�J(����K�1s=�j��^��8����I�r�m�x�.S��D�S�����*��s	,���L��i6�q��G;�QIm�h='�'��[�{�h-�͊�Mj~6P�?�Y@�"�l��.lM��O$�h1�v6����4Y.���X|���u�,m�.�d1��\&���Ө������7^��/����@pY�Y1�W��Ý�vk�qjT<�7�u�~땗��m��u�K{�x��İ�Q:8��|�ݶ�F���5.�>&���kY�-�40'��V7�Caz^:�YA�_~��9ʢY�V����ґ�R���G���͏���66���?�L]� �E�
u�a����}3���ܐ�ǟ��`B�{��+X�qo����-�N�8�wgS�������PL~M)�3�O��;��u �:2_��e�a�=a:Y�(�0_4���-7�,�NYלt6����1��M�{VǽV�	"0F9l�&:��P���u�y4z�w(�y�������)d$,�d��}�]t�K#��WM�+�4�l�R
�����䔄�;��"�d�gI�eå��y	C��B��\\RP|:SD��������ݰ�:1��4���VĮ�W�����a��!9?���y�Ř���y�GH�k�#����!�CE���ؖX�G �:�(��4v� �	����#����r[���ǁJ&�3)}&��Y,�1b�Euf,��,l�c��DN��q���h��]i�%�J"�iDs����E���aS>��n4m��4�x�q-���4�����Y��{ll�a㠇o�f������<�y�{�U�,*H��8}�"�]y��\]��ý#̟=%~��s����~	O�Ì ��ￃ���ё1�Lfp��E���ᪿ��[���G�#�=����a��#�[�ov �evO]���HID������	��@�f��u1�+o��~�m��Ĩw�y8YӴ����+O!�ыg�����<sׂ�`" !͒J���L*������4d!]�鏱AƘ�>�\�x���rݩp�(bg	��k+##���)C ��)�^�y��+ ���	5���M˫�âM����i͝Ǖ��(��5���p֨+�6n2 t�-��,~
��@S)^�Q�j?�B96�?�[�{xL�wL��n�Q"�f�~<�N��h!)��� �{W�]���P����������͚�zO��(٧D�\KzrN�n�Q��s���h��'[��X���T
�gΣ[9@�aUN2���b!���7��)+X�C�c�y�nD��l����!�0�"=�xs�*)#k-I���0�,��hvů��j$e��k�}�>�v:�����6�?���U�Ք{of����bYۃ��dh(Őm��Q�=�{��fE��D�4��:�I�qT�c�gHf��XF5�B"�O�<��8�<[G֡�>uM� A���D�-��XEs��U�z*��/����i�=��jmŉQ`t7w�pm{��IL�=���{S;Ogf�P�����5�����R�4R���⌼��VC騌��#T�M�=�NΠÔ�G#�Z�;���瑚�Aaa����Ѵ��)͈������W���w?�\�ҧ�)âa�R�{k�f����I)�n��6��cg'h���ӀF0��w�p�5��'��[��<������iY��DDk�c#�j#����z�����%k�F"�t�����#�Yy��t��A���~�}�1��o�C�KBPyR����(�xTՋ�C���z
z��^ϰ]��o�ӈi'!��c1st���j���H4���&�<�c:�&��G�k�j7���$!6�:{@�B㰄�����l�F�
Θ�A�(*�ޡ�t���i:=j�;BJI�bc��9�b��:�|u鹚�t����g��L��:t"��D��ȸ*��vd[�Y����i	�����'ˎ\q Y��QqL�m�d�����6���Q�TC�<j�b�Ɇ��A���s���aȸF�[�Olj��U��^�nII�X2��s��Z�Ͱ�7Nc�2,u@�"s3z.�� ��-Μ)�H<�s�bD�Kˁi�R�������4�Dbs���:X�9Dp�~�~�Y8��<4Ĩ��	x�r�GR�񹧞F#���:.L�ص�:�bouM����U���^{���ty������~6k9��|�Sn:5�F�NË�ɏ`��S��ݐ�S�5�c�H�@�HD�5$x�0t�S�%��x�p�#��G�(�H�o�i����9f�i`S�aq߉$eP�Z ��ۓ/� ��>���`:�!ת���zVi�T��鉹�LF#h�`8'5T�?Ӭ�>��c���a��Z�@��;�����2F��`�n4����~�-/��Κr������30�L��M!5�,#DT��'�cq���Ь7U����yG��9����Z:��J�4���PMk�g.l��@�������v��K
����PA���h��-�G�tM^\6�ԩ��[�|���k����m�(�S>��g�I��nL6��$�K�p�&��9�U>� ��＂|"���FX�,wV�A��eU�R1쮉>��M_�\'W��`�m�
E��a���j�CuƆ�*>��Ԗ�AԞ�Lo�:~8����F}x����3�X�N?أ ����C��b�����:�4���e&�h��i�VJ��D�,����d�)��ܕ��u�:��&j�,J�}�"��'(ȗi����D^a+�w������$
��G5ܸyC�-�)��߻w~���B�{�}4;=��6ju�&��<��X���[���Yu�^F@	#�XL����8l���i]IxL�U�&�EZ����N]��MK*ea��J��v!��n\��Z4*�&���y<?��3���	�Wnc�ʖ#c�
c�'�Nk�L�#F,�qS�a������Er��W�oFC��/
��|УR3�\1�����=�P�Ⱦ,gJ݆�x}��w�b6�n�>�jx��\��n�'n$T?4�F}���������W�U{:\���I��=�nB��S�2�t��Et@��t�'���d*�i ���( ���.4"�����b0�T������@�k;�(���$��))�t�F��x��R ���P��F�D�WE�|hL˽�$�xG�K��~A�I�.�_z���N�kJ��3�V�q������ƽ[7�w��`=3����l�H85��0ܪ��>��kc�37�f����X�1�7�jc����4P]�pC]3T8&��^�wb�,R��LJ/��r��i"�$�Fڔj�:T$*�[��D��c-bso;w����~��%A�9�*�pxTB<�����md�\
yA�r-�S�X\>��A	�lFSD�I#�K�DJ�q޷v*85�((u�j�t177�씩�Q�;p��.�����5|���abr?���pw�*��̝�Q��s*΋Q?��E8��8��a��f��Z���q�.��W�#�>4�LF�����a�W0{�<r�3�[�%;�Mf�@1��~:��f�`0��)%��gV��Ʒ������ ;����[]�QݼQ�,�1�NC_��A1-�B���yb����E���i����9��O�����덾(K����n�/���v��+��z6<P=bU"�v�衘�QCU�P�#L�!w:F�Q�����1%hʦZ�?�n	"g�D6�/p�J�j4+*�k��@�v��kx��w���d.ո�OC6|ywKX��T��l=Rm?�z�f�:�e�	?FU�(�1�'￰��0�,U�je�Kx���ri_�j��s{F�@���ԣbRzW%t��������Hh�S�ܐ�;-��ԩ3�F���2�!�44pm��#����i�<�������5�y4����D3o�J̆�O�ρ�%�3�M
(8��?�sT���VL^��sI��X��7<XEerN1�b��!n��.|�U$��#%k��C�.�u1������Eq�+�¢jcY�5g�禵~��h�)Ψ�ES.��B/��s� )�{k}��<��=���ٕ��|��S�F��5�����|wn��nJ<�"�̘�d�qj�O<	O~�1� �<�O�{�)�:t�zJ9�\~
N��}�L_>�L!�FΟ>��K����o�4s��]�5a[��,�.e=E]�,�N6�+��qG�������r��1=3�<fm#-Τ�{����:��	cg*A ���yCk�}�c�g��ǱT�W1�_!58�磏�=�bc#*Mj����
�fb��]�QE�L�u؀C6B�QO>�L�?<�������*&͑6��>�r����ۂ[Z�d.�V��-���1%�#pU�/��#�����[xO���֖5V6"g�WΡ�n�u���,PGPs��'��cн�f�M�;@�9)��7'�UtQ�
�l贠�H��~��T�ł�6#Hͧ|�̼��vD��#h�%ⲑ㚪a��N�H����٦�/�sn6��Fu�'�k:5���OQ����0�V~4Oh���O��Q)YF,���k��a�ٜ� ��J4h�3�4t('�0��Q���q�W�����n��#[���Ę>���V�J％m����2R��vGFwmM��f�u:-����
n��6{�h�l!!k��W�����_��zA3WeG���A)�H���΋��8>��X�G-��9�둬��J������<Y#*]�q����_��K�q�TWM�p�� ���� H�<u�,�rz1Fl��G㙌��}M��	�e*w���:KߗS�����)Y��x
)���An��k�*���|�22�y�O�(2}+0��"�Q%aJ�ӳ��	v��?�#:<N,ԋ��c����o��9s�T�tM��uI��Ȣ&Zdx�V��g�N�4<�hFj
��
�юv�����ݨ�vOѓ�7 @�.�,k���\ώ�s��]�Y��PuG��]?�êә��u��n+�RvF<��IQ�N�����Ĥl�"Zb���!yT'�{Z�36˖�3��遄��1k[WeQ�v��Pa���~:e�<1�'9e�}l�ƍpF���t�PGL�ڮ�P����k8���t0�i��l�׷�x@o<��;i��o�mH擛����d;�u�VJ٤`"�	����D\��	��Ip�X�d�_�yn	~p������5����)�m1-�����C��βo(EK]�v.S�b��l~��>�`�B���<�������// >?+(|B#cD�s�t�I��ˊ����pD�V�'h^�ع�g���qE��~�ӟ��?���.�%ʊG[�	@鰁-�EZ���o��K8`�C<a:jS�5�O�0g0�
���j**!F<!�$�hC���g�$�0�ͷ��"�l��I��3&VMXS^�y�F�����3�!�\��P�qG;eþ'�j�����ϛ{��È��aD��6�FMw�	I3-�76}F�_���2򃊴9>+��s��,&1�94�{��Q4�� ��r\��(���;��Q�N�S܊��������񵨕�$�H�4}�Б����9=dbԔ�"@����[7���l��0.�9g��x��Ulonf	;?�!�k�(?�(![� Qh�-d�&��t���}3s ic�Ԃ�O���W9@ZB�x��t�h�G��DXp�{���un�f��K�f0�IC{d:�T<gP������-N&j`4�Y7�	�~Q����vH�}�}
����p:>�w2P��.RO�>��N�N~���k�*�5j8�n8Y	f8�?�֍M0�+���K���������5��̉�������4Z���e= �����l$c��c�κk!wĨwo݆#+ ͊�B�c	���&.�O!�E˵zP����)��q~d�ʋ�LZ]I�b��iLOO��"�lp���_��s�Ω�o2ES���obd��. :2*^֨|���<�I��u�h&��Ei����%z�|�� �FMx���y�صm{p$a^�Dv�:Z�*�����z$'HD[�?���1*�8=��|f����y��f���;�}p��W�0�珍���-�i�&2�8�EVj�PC��w-�[�~lm~AC�?�xܻ~ʰ��1�?����OCO8�8���Q��m���n�D�V1GQ��Nx�0TC���"h,j���j,�QSy�_"�E������-��ئ~w��gE󲙚�	I������|�!( ��J�������G�U���7���>8���p�����H?,��TG=Jقf��U\95������,�����%d-��4��]qrl�f�{60CV1*�dI���ü�OUnK`� f�6l�j�rdr��'�Z6��T��}�	��6�rb5C�Ӕ�a�?;�O\+��bl�L��Q
Y

��#�L*�����ݜ0=���Qf�A<W�Ӂ<�f"�Ϗ�����(��a������O��3��  ��IDAT�<!�T�`|Sx� @�rc��U��#b s�*�Csn*�棴��=:{Y�ϜoR�uؽ�M�o^G��+����L�B}rѡ�L��:]:����ܼy����(LΠ�袛�b��9$%Z�0�f��P�����v�9�����T����u�=jc��5�?|�r��,*i��^y�
�_���jM���N,fXKjܣ����H4�v��r��=��5/~�;�%����r��&��p����aC�N�r�<�LO1b'��D�����un��A�Y���и�\�_�x�Ը]o�cj=�g�yz�F��A�2`Lg�cU���i��4zv3�nĖ���|�tqcq�S3�N�q-Jg���@�G7�#WH�D�O�M覦.��*rsӫo��(ڙ�_��zM�?����\�~��,�DR��uZ;{�|h˼�k#%��p�`�	ymLLF����۔���|_���z���F�� �݇�0Z�����5�����~�S�^{U�!��ќbKN�F��h�A�)Y�Ξ\������<������x:�����h;�N/P�OϦM��z��)3}vA�4�<�cYmK����_N8���O(��ӴX`��-�:�gب�ϡA��)>�S�y:@�@�ؘbcDxĢ+�	�'0�̳:�HQA#f�¹���:��[����:�x����s8�o�P�{(�<23��{w�{��#1�z�B�{�҈NLÏ��F�x�L
�[�޿W�{G�g|n�|�	j�
��Gjc2i�'�;�)e�fe��CE�drzE9gwl:0X��N��c���ıvd���)��Q�ϧq��_��7_G*�
�ސ��Q�0��S�1�)�H2�$�E8�$zq3(�f���r]���'?Ǟ8���F��C��F�A� A���'/ɚ�s��U�M�Q�){+��p쬩�XR��3ӣ)q4ܷLSU������-*Sz6E#�a��\K��d��F��ÿ�YĕG�����\��<�ᆥ�u�������C���Xa� x�$����WnӘu���$�d{q+��5�墆�,^��-�z:-�;an��\��x\�TRd��3̝�Ǔ1M�0�������ﭬ���E�:v �5lv�Jı�]����Fƈ/�dQ�����$q`��`7���X��ü/�����K��q�����\1������N��ƒ*�%�8�YEה:��f�"_;fBe�Έ�W�o�8�h#�¦��|69�ݞ�#���*r=M��@� Lqe���c_�ر�6诹~L#��l�&x�lڢ� e�F/�s�T(r�;c��$�]�X�<lX��0+��07�&�=S.���5��������T.���*{�*S0{���6���(3
tcj��,��=3ǔbr��:�ԓx��u�z�Q�pk	�Y1;��/���h�0Ah��>+�*���W_���j�Uܿ}W�L�?\g�z��W�:삒����f8�@��s����g<�6���T������>b�?7zjyo*����dݾ��U1�א�`b$���[�gR܎�����{�����-�#:RD�I���y}��d�w�a�� �R�z&=�� ��U��Nb��9��P�<qd>�潮^2���70hY�R\#HT��K�Na"���L/JZ+w~)#ˮۯj�w|���a?Y��赇��<N'�!���8�`�۴�oML`����щ"����ʂz�s��ʎ�)�WL�Y��3o�긚��_Ȳa
&f�#%{-#��׹܈��G\�`�7���B~�������ٜ��`���y�j؅ڨ6UH+�}�hS~��< �e�o�aeH�K�%��+n䇵e6��5�ߑ�h
��F�}�>>y�T��-�`�\�f��5MU���R9DSYAg��EU�J�p���w��5 �9�k���ꂨ�:d;&F��W�C?>V���^�A������4�\��'U�'��̶���"���u�-,#F�Y�XP����;��p	)�±�r)�@9Y�oP�1�Φf�|�0����i�M#&�v_"�� �ެ���8fi������Ie_8f&(���Fo��;]5y]N��ԓ��ӥ��D��2���c���H-/G-j�E� �"1՜ᘹ��O�塐K��'���{7���'��i��m�K�XՔe'j�&;)1��:���|F$}3}�}�a�ksׁB�m70��������obI��S�\@y#�<17��Q_׍r�cY�f,��emƏJzMQ��11�=9�Q�*�>����un~YO(��~ UTs�앎��1#�,%� �U,	�Q���ןA�����"x6�Ө�[�����q[|ոt��:����8$��NŜTT{Կ��9�}����� ԍ�n�� b���J���ĕ.�k�ŬҞ�ь��~�Aw�Ń��}�Ļ��y��t�Ha�5*��K�_���0r� ��	���+W*���O�h�x�T/�%���׷	����U�䍝��<H�?�tIA��^���ꀮa��Z�2�yA�77���5u�����>��]u8l����BW����"&g%�.F="���kb���@��ڝ5��܄������h�� #F>Z/�m��ￊ?yz��㵍��mx(�-)�k�c��ȼc9uS��?���X�|���4�>f�L�o�t�3�B�f����}Ȝ�Y��a�=|�3T��Cm�~~VG�UED�s ��������6�����������R�c
�w��aZ�.�������KO���ͭ��0��/ 91�#��f��5CR8��cz��]q0�����l��ciq��q�� ���UR����[ڌtpXAfl��8�LF���^Eh�t��:&:7�x�{���q�g�%�|�8�M���?�7\��k��Ûr��>��Iqx-699�s�a.��n�atN2�������I�}WR��v��rN�i��	�*N ?7/�s\�@��Uͤv�DvI}�!y2�w���l7�d�k#*g����B���I���"���a��q�����F��w���H���-;�+LCx�{���˕��cA��<82'e�Ҝ����:L���~P��&�h�k]MG���=y?���=A{%սNƣ�	�?��vG4;B;ʼ��(j>���۸���W��ȣ�"ϝ��� ����z�����QsS[�i &Y�������wK;-�v�5ߙ��sX��l ��!��%�B���@������� N�ԩ\~��ꝏQi�����9	ݣaK��|s�R[�z��G��=DZU8�R�$�^�S�y�����_�@F=��]ǤB�L��燍D'�7�sb��Ƶc�Ȉ�a'e�&Q)�}�<�>�w�6����lF�bږ�9��̱5�ôJ}J�i�bV��D�)�tLjȳi�p��Q���0�ɰ۴#�p�92?/ד��FL>����)��-S&�I��t�V��(P�E����(�B~�紻tkc�V���W%rH*��Z���?��������G"�������'�j��H�4�c���I��z1��&�l�{�}�h����񈇼��%���\ڥ]U�"�81m"y� ��D�k[���=,�Li�L9���s��y�w�U3_ ԃ�u�O�;<��W��t0N̍��o�:�X}�f:�v�O�Q��o��^��QyJ�O��Pq9�3��μ;S��;i�tʁ��=4�3��������N�|���v��8�[�?uv0�Rʹ�㘱v^_B��k؍���!-�3H�:�j��L.vst,2@����́�ofj5� �]>"�%.����s5Rf��g?�w���ŋ��)�������h�ƖZ�<7�����i�c�����g����I��j�9�Qfw��ldvA�k@�z}�(�SP���r���������d7����HE1�O�� Q�F���H�%��e�7�TwnK��E�ZA��!�(���/�ܨ/_�!r��)qb�H1�	L�Y<�E.{gf����}ՔQQ.Ǳ��Fp+j�f-�m��ܷ�����'È�ڨJsF�Ā�R1��<������@�:�9�Jb�����07?TS����=�xV,s�����Y���0;m��k�7�����h�c-F �3lu�!@@NwO���БȬ'�@��!Fg�A�L�������y
A��k7��ڨabrB��	Y�-9�1�.Hq�"����쉡���fS�����}KEU�M#��Yxn	P����"���IY+7��D��������N/��/�������ϩ�Q\9s��[\���V�����>n��DZ���c��t"��0vN�{�Yq��aN��aĈ��~�U|������u�pMQ��2���!�v��L׷���Y9k ���{ݬ���)����~^�B.�x��8^�:�7�?�c��ųP��{P�WN��~�!��C�٨A�D\6QA<p.cF��4�Qd�h�N�a� �������z 2�\ �ϰ�_XӠ�>\������x��g1;;N��	�gS���n\�n�����j���I{�êq��,6�����ݩ�/�ؖе���S.��͍"���!���n�����.&���x�,:��k����k�0��Kؒ���'W1=9�w�y��Z:����8\�F��R�tz�1�-�8`N�\�����0&�TeO�����9='������6g>7c�Q\ӯ��VX�/%D�ǋ�Å|C9��q��jwښG�B�M�/ck#�\:EwE��6�}˴9��^���Nh�ڪ�մ�T�j�
�1��xF|��EWΦeq��X�y�v�����ވDS�D�Y��Tĸ�i4��8��q��q�(a>�e1Ь�-߼�̈�My�\���4x��+*�FCtg�F� �ٛ��軈�\{/���x�Ś����9;P��qH���)\�*�|�S����#��{o##����vq��y��?�Suƫ�VUR�⌚����*H<&(�+'Z`wsT��%�jtb/��c��9�Jԑ�3$�8��:�I:?��@��as��e���6�
��e�xf��g�PyX�;�w�z뵺�c�~*� xv�Z}����:�(zrS_����:;P�n0s�̷�}�#�z�h��JS�
�8� ���r1�7s���b�sv�P���7�z	�F:�Daj��s��h�P��/�NS5���5[���۷q��U<��������j (���'Q�oY�I�0��E���]�� ��y0%���̦v�vw<�
�gCIb|��%Y@�9Ǔ�Q��_[���S��$]4��n�_���w�P�ӛ:���ߺ�R'P6���	�{jD�{!}�l1��Q��#��6ğ�������W���:vJr�b\�:�)��ϖ�8L��]�v39Ǟ|0��q�Ms���q���"o��P�'���~G��3	K#�����i�զ3h��YXbf���7���@����H�9$hP�:Awє�[|�.�,�@S���锩��3FW~���T�#�qg����(f����/h�\ŉ|�|f���ב��L�ﶎq�������P�����&��w~�)?�_�b���/�B��~�F�xL6��M:��kTA"g�
�/m� �����!j�N_�$`��X���aM��gT/��Xp@:�������������K�������w�V����Wq��i<!Q�Z��� �����i˵��zN�g�cV>���MMU�-3
f�/� ��⤷�= !?4�&e7�s��%J"��He��u2h|K���F��������2ǯ����>,R|��k�M�j���i�*eL�߱ΡF�`P0�E�d@�Щ���X0�mGы��n�C��щ���Iga>��'��gRֻ�`����>�������\�+
������4o006����5������j����^Uᰆ����eg瑗�$=;�����6�%��HV�1��R���ҍ��L��=�����C���[x��|���3Ͻ�F���I$䄨�����2�;��@z$% ����.
�x����-�w��CP\c��NB�cb���(��C�L^r �;���p���"k;���7���+`-���pjH��bP9� DP�9��I���,o��0��y:=��3K,$���p	��gĩ'���"�N�
�q�z�5k��sw%A��8#�m��
"/��r͹A�p�{
��UXLJDFm#�q�s�̰s�TJ�{�u�*��|��B��>�f���j���G��?'�v��!�"XG	����^#)Jc��|%QZS��_��,F�)��#d������R�����
��p4�s���U�n���W���W��������x(k�r��~�!R����>��Ʈ<�&f��.�Iԩ}��FGYO�D[�)��/u/Ѱ����U$��q����z8�0��;��A���#v��b�YQ���6���MD�dҨ��Z�K���c�\��R{nX+�?4��16#�p��Q�?�,T��\�SW�E��00�P�?Cc�d�Mqm�N�7��@s����uD��|��TpL�����	y9U�݊+B�t<�7�RⶐO��+j\~��ںM��4:[�ȃ��:_�9a�k~XC�Q#�F�^A�w�+�c�+�u{��q��j���D�������;���
n��N^8+�~�g.�`�H�Wx��JSb<؈�@�gg~x���l����ES�vC�\(#e��E�6�)�1�%F�/_���>�n���W�g
�1�B�<Nk�Y#�qџ�:����yc�EɎ�lR��X�W�Hx,�A�)�suC�G��wm�R:�Q���b��:u�=v��������>kI�|��7HdӒ/��V	�	A�3O^F"#�J���vp��DG��o ��hH�PH&�9S"���lU��k`�YFaq^����	ep�oν@�wFe����RI�@^-���Ks���� g}�䳖���
z=��4�e����R� �1���9/�������?��~�&p���+�ާ���>Z_����L�M�lP/)������>����4�X�^ĩ�ps����n˟�X@={A<�*vq�#x����"�񔬷�:���p2��Z���q����S8,ʱ��M�:���F=\W'�5Oش��⎱��aS��`8�ؾ�A�i�oLǰO�{�蝩B]��4�c��u���a��RA��ƽ_>1J���ï�Y'B��N��˄9Փ/��X��T���fv�4#����c`�k
G��1�Dy�b��]�O����m�����C�=�l�:z�67wu́lJV�`�����O�DQ����������9��/�|S�N��r�"O:��D��Yt�����Sk�hP�1&��?��ulO�:�\�#	�?���s�̦��98�6q��=LM�#/�grn�3��׬=p"=E�nܾ����X8u
��<b���@���TE�<��3�n�1z�I��(������]	_�iA���GP�_�ʦw=MǨD�c���[��p�g7�d���Z�7�s�A-��l[���U�jz. �D�j\�q��q�:1h��B��fޭ��i�H?j���t�5�5�|�r�r�,����[��U����X�j�yl��C,=�"��.	Z�c�]B��lz���f]<j	E	��I��	SS����8g�!������DBw���s/at�J�*�a���D,3'͵O�F�"F�����"e,�x�u��<��󚪣��1��#�	~�)��S�:I�s�w_ё��c��P��Z��]m��|ޔ��m�YB�XvjN"�|r�:Vo��x*�?�������/��o�Y��	���L΢#����5t�9��fqԖg�&k�Z8fx��,{ƩF�"��Ĥ���qOS�l"���^<��L)k�정a�ap�����y-l����!nv��Ұ�3h��*�}"�'��}���>�;���vҞ���?vh�Y���3�_�0��2$�j���:�A�7�9/'bub;6�X�� o�5�����9��j�k4U�Ұ�������{!o���&'F�a�h�qo�>��)I��x
�О�@����V�n�-�jx��.�o��џHҲ��VH�0UkQ�>���%���*a4���3K�v�Q��,!��v#�*�J�U�8�1Q�#W��FEot{��+����dsAR�"(�t�Gnj�����i��1�9m0i����B��:8���Ц,ESW_^XͲϒ��d����s�HY��=��j�$N���|�H;5q=��^q��HO7Tqx^�6+YQ��5�}�r�G[Pd{DPoF~v��=�]��2dq�E5��k�v��#��jxn|9��mA�G���$"Ҧ#yt�L�&0����ʚ�בs�x���HFQ���WP�AWe6���F)A�����5�$=P�9���>���A�^��f%Syqb��9�&r�~��W���1�ۅI7���w-���lv1)�׈3
���p3D��.����a��EA�q����Npz��
�|�E,Jw���c����S���8���)k���;�I1�́�U�Ώ�*E����40�,�)r�\v������$2��jT`�}:�+T@�[)��C�یc����ش�Aˁ�3�5�L'k:X+�׌�䙞	g����S��Op�䵕w�����~j��7s@���'i���A��%�Н��Cn+ԯ�+��%վQ�3/̷�I8�!7S,M�E�Z��2ggD�^A�z�2��cb(��Ȇ�LV	���Ę���I���6�z��:	�=�
5=`eJ�o�q-:�62G�;dsv:��1\ŧ�j�LpJ��(�R�b��C�8S�v�����Z@c{t"iG���rooo�^�a,?7�d0%f�B#"�'#��u�8��ƦT���!N�����@�N$��l�Nװc8�bi�)sLA+2���(0�Hz��A�</%;�6�(.%?K�1����[b��b���jm�t����!�6�N��)P�	�7%�?̈́	)����X�M�}PB��5H�	WL!�K�h��r�]���ܳ���l��i�}!��\n�\����&���]�j��TfS��xZ�C[�G�se_h���$:8�����!QS`�ưP*��;��ZO�0�ŏO��[���tYz�v�z~��U\�� ��q�[>g#�8JT��i2Gj�9��S´I��i$�������ڑ��-�
��ߑ�N�I��:���G�z��,���.J��Gq(�P��Z�鎏�-Ǝ�X��g�z��S	h�0^z��[�8_�ng��8�DGN�Sꤻ=_�%�9����2�"���_!-��ԇ����#
������?��m�y�k��e��h]e�#�c���I�y r�4�]�O�e9j�y�Z�=.S��r�qO�2�]#ȓC����Ǡ�Z�j��TX"5�8�FP�Y�¬1�f�]���8��L��Ք�Ӫ
��:=�F*���Z	���p��G,�ޮ�!Hq�R㾄N<	G6	�Ǻ�����XD'Ϙ��s8X:��#��s��I3�T���d��bǤ�"6�͟�[m��\y�K��-��c��G�����(n��I�1L�V�A�)�0�����xyi��
ȋ��\J��W��NPn�d6Ѥ�1�����~��.N��nM"���욬�fm�h�����dl�L٘*�^`�a�%g}-�g��S-!h�0UL���<��z�)�?��P-r���ӧ��ݨTja�#��)a�����-FE��o�	����fճk�(�d�� �J���ds���qh��>��.��+W.�������*���E�!E�J��ժUPGn*_�l�R 1���=.�k=�Or����N`T�0�)�$O�/
ӍONi=��;�j��Lȹ�X�u�^���)�|9c��/a��IP������姰���Igq����"��IeP;/L`qvͩ�ؽso�_�?ܸ�9y.���ۤ��[q.G��uu#Q���Qg��"�M�:U�^R��ۛX�~���H��x��g�t�2��-6��$����{N��\��s	�XB(��Q��4h}�޹��!ƽ`�3L˄�ő��E��:�|��H�:�{���;̭��\��P�����}��a�gDX"ͯ�U���[ۀuB�iZ2F˵��j�M��xȸ�l J��5�*p�&�ǜZ�D�o��Z�CrY,/N`v!�ŝ�_Oܴl�$���42�P?�~� ���r�F51�MvH�F%C�i�;2f�K$LZ;B)4��<�p�# y��F�����"C�_�ȶ���A�~�"ө�2�ݮrÉ`;�|�&�,5��ds�f�l���kC��W�������+}ytY���
�J�je���4J�*��\�-�-1=TQ�n��L�,L��c��d�rc'�Hx�<=��]��m?��3X�����Ook���}�b���=s����ﻻ�3بqP�DtXDwLw�.�B�C6�D	#_lכn��nx_�d1?��'�`��}`���&�h.��r��zM��#q�uE�l])�`qj���<*�k��Y^ƞ �{+w��5�� �� �b1� ��k�.�?��v��%l�v�r������x�n޸�?���Q��o����w���$�/G;�K��?uo�$Yv����7�5#"��ڗ����nt��`3)�h6F�D3=�E���@3Iz�f�D�C�� Ďnt���Z�r�"c��.��;�FF
��<L�egUefĽ�����矓4��@N_�R�u@;�ui�����nZ����ޠ��x�����+W%a7:=�����u@@H�$�ƺ�k��tM6W֥׬���2	�5]���|�jU�7��BO��n#��u3��&�P0ՇT�3W�~"���a���K�o|A޸�!�����%SY���"2�,���k����U�9�����/b)�A>�i��Ymh�
,����ə!���g�:Gt9���J��Mh�����@3���I�XŦP�ټSxF��b�Y͵�l�B��gǦ��D�jm��3q�=h��8�m�3R�{R҇5�P���{|M����P��\���C������qt3��%��$��AN����2�3l7$��l���0L�w����-������8��L�Ā��ڈ#�s��KfBW�MeYw`
�j���]t@�)4�8SE�Ȉ�S�(�ڢ'�B���Y��H����gYO卷�2�u����J�7bz��-J�� g�2={5���+�q(G�\�s]>�9�5�N�p�ʐ)5���	E��qK^xyMn_Er�����Mi8~�*�t n�%�+�W48IJͯ�FE�����C�=	S]�!r˾J�[��s�:��h�s뭷4zs��w�V����n��%��.K��r庴F0A(�߫���mr����
����˷_��'t/ݕ�"{��j�^y�%��K��l7���Si���\�X�Q��ӰPK��B�F҃(�o��0C%Kt?cH6[�j\���J�]�A���Ϣ�k�^Z�뛗�� ��OѴ���yl��%,$�(6-m�j�~�I(�)HV����K�at&L��5]��p���Yضc��m�.p�������ȇ~?�g��GG��ߗ���W���$}a�EZ�(=���S�8�YC~��|>�fE��t�k�� �d���bH��Lȡ/�{d	� 3~��Mk���a����N|CF ?�u��1��`��B�D_Q���)���*�?=�=:�F������P䑤R�YTv�o���'����4�@<������y��$E�/�e`�<�pG�moq
:�DF��t�����lɨ�Re�.�n[|���"e���@.7�Z���h�&^��9&Tt�j3��\���93)�<���Mg�0'O!m��q��k�Q�P
I�̡[���)C��H�'�R,�g�����F�u��N[���DK���riY_H�X��z�!�bIڒ4��3rk$/����t,=E^���V,���:')�K/G�Yݔ��EY[]�3BDttp(����~�rA.���L���%�Rc��Pc����H#����P�� Aτ>Z����F���l�[�����\�⛒\Z��:r��fKE)�,I�Ve�鐨\�Ԡ,�������z�A�}��"儤r)�Ө����կh4�g-����ۯ0}�w���l�J*����i�IS���=��,[3
������λl�Y_]�aGZ��׆	`7oܔ�����򣟼'�'���bhE�^�����}��4Zp�F�;m� �� R�>	M�+a#��|(DD>jr���`�t���g,�#X[ߐ�~��7���&B���14<��u��#r�g��d4�s��}����O~"C���^/����2Es�Yj�:�g	�����	<G.�:��"���NM��c��Qk�j�ho�kh2��5�g��RZ1��9RL��|��3뱟�O<��j�7�,���s��Pt��,�E(�K䕣 ���ӠHq��o(Hn�e�u�v(r�S=Z�5�'jt�� �減�K�C������'����]
L-
h�9��BVa���SI�B�s!+j�G
��ⷻ�9>�
��3E�f �gH��ϑM��l�iE�����yVv��"N2���W��?VG��/#)�rMq��)=lI�A�F;�D��4K�A�][��@�1��P�@?��uՁ%2��.�TT��ԥ�TZ:{u�(�"�1,*�K��hT����<�/m�SD�0�A��ѝ�.)b���y􎤷��:G����Iɻ�������'g���ǺZ���W�8�yR?����(Q����0��|m���UL�؉�l1����h�R�����_��K%�I��>5�|�/
 ���8�FkK�����p,O�Nd��Lѿ��k�շ�̱����Ljp7ը�|��F�%Y[^�iz '���H�'jԑ	���L]���Ϗ�ܯi�=��!�X���Y[�?�1��8=|�XV�$�߇�$��l�>'FGn���!��0*�*C�AB	f��@�����ڻ_��ߓa��Y��a��kwt_�EN���ٔkNXG�`�ls&��Q�9;����o4(���(E�H��eNA��6�/kJ��}���s<Q8�ԡ�R����Ҡv�7
�� �)3O����A|�gC���3P�W��逡m�1yu��d������dň�y�����+��Z��l6ekk�BN�j�遴"x����mJ d�1^[���=9==��Ϥf0V���-����ʿ|[�u��rL$j���=Ȟ�f5U�E!�q�F^@U�R�N�2����+b�!�yz"-}O(��.󫱬@"2�y�0搐��Ml�Vb���%��0#�,p1��R�l1S�Y_����\^�����3���\�\F[k�z�9��N��iT4Q4�$�h�U���8 CE�ӡ�>�F7d^��Y�zS�~SQZ�Ҭ���)'=a 4~�?����C=��4�k����l	���\\*2g�vZ��Q���IcЗ�D�@�@���ѣ�������k�22v4z+֤��)�rU�U��ej�`E�|�����qH�ph4��t���⩡��d��^o��jGrH��~J+����*iE��Nȑ�u67o\��}�7X��ַ�B��w��.���Ko�s��Φ����F��4f�
���CG���x��A4�L�#6%1*ӽ����{�TvϠ��$�!��h�ϝ�=n�='hP����U
@�k��J�LN��@I���Oe٘SR�u��g����Ǌ��b�I�y�o�����-�}�7YO��;p�Z��Ke�v��l�1����sr�F>m@����r�7�q�M(�JD��g�Q�����3����sISx㟳��|���5������5���Q~v��?�����mn2�L�� �1pԌ!8��f���9�#5 ��@����{xx����`$����E>0xю�f�\���#l�)l����D�F�)��dw��kE6E�v�Q��:>R���D�RZ7�g�P\��ʸ�^��S�Ї���*��+�UKW�d�\�ݏ~&���L�w�w�wMN3��q��S6�0g;m�z.�qQ��^Q�]��y���J(Y�(y�(^!��d�Rc3��MuL��I�4���y�(�}��D����9���F���#� 2)���N�\M�R@/9���4r��בɠ���?ƺ�s�dq0E� �A��T��I�p<�OI)oP�T����ə~=�J�*��S�)����p��$jD�EE��E��w0�M�	�N]̆�}����S1x�yL�Wd��{L��o��I�Z��z�1P��.؂:���U��o�����IG��rp����浛�a�h4��䓻w��l�u��*x����.�^�瞥�|�i� ��D��B����D�Š�k�H�D=5�i�y�?�3H�J�2�J���5�:41��9}s4N�0��Ք���]����vx���������8A�t�*�C��I퀤 ���5���˒�=��"=��ۨdK����W�&+�N}JD;�e{є3X]�<[@��f?��yvd��O�q��B������M�Xp�8�<05l�{�%�9<��b��tި��$��Z�52��R&�����X���(<�
c� =�k4MW)�!�Ҏe���J�ӓ�r��+<���c9ST2a�U^._���h+
:��ȉ�e��S��.4S5�Fa���a����@��׾"ח��h�IZê����=C��_����?�D����E�RV�P�.I��G�xE��[��i�ǡX�-��zi���+�U#H�x�Č�9�&v�/�٩J�u���r��#�bd�Mo6�U�c�Q��U�v|3cV����|��r���wG�}�\_i��,�ٞШ��-�-5�cE��I$��"7�Sd�
��h�H�FjLR���ײ^sO&]0
�F��U#��;'�G�� ���~�.\4QeKj��z9S���ҝh�k�M��;r}5+�?�AJn��)�T����3�z�j@E�x�n���vd��`4���0�.�~V$[,)`(H1[����
��K�Tg�TLB�+ԗ��.ˢF����������%0��L^�|�K��yIꊤO80����Tj�`3jJ�!��c�^Ǒ���LC:S'_��<���
��ľ|u�m���e6 5�r��^Yih����i�1���O�v��3ކ����8=0�>;DF���=��~Fy�A������h ��ddT0��q���b����ݼ&o��+�n���R�@7/_���:s�P5�"&F�uu���aH��&��8s��X���>WA=�\s���}�#H'lN�V�R�������"a���s�>s�񟑙��v19�g�D�3ұ��f�T��c�a7q������X� �ı
\2�DǘC�=�؅�\�Y*�Kf�gKuH���р&ƚ�Ц�4�ҘJ������To��l��A��Wt��B��)�Yj��~��;�����lR�V��y�'�W��7_�V�T�?[����=tjX�p<���zx��醆z"r��m�o���^.V%Bl颤��]y�i�q����șh�nF�5-yH�EP�����ϱ�%Fs,�F���mc�S����#}S��zE~��ߔj�ca��I4jWfQL)�2�F���$2d1��ݙ2e�1ErjDkf����1}���XI�V%�FyI��У��ϣg��􀌆�\It!2)��Y�H�y"��P�>�S�?R��rX(LS�i��Ft/s�RxqnT����[u7���j����G�yZ�z1�NE#��Ʀxˋ$)u� ��T �V���K/R�mmm]�v������_{]�V�8�������6�[X����������-�$���I���֖������"<�Hrd�9='c�����\x�5y0E�k�������lL�R�n��k"g�rt�+9_��X��YhQe4��u
ԏ�B�Q%���� oV���qX҆�a�L�K˒+���t�$;q�T��?��N4BB���Iv�F	���> �J;�U�R�0���8�x��s������2Y�Ⱦ�����$�,�sl3��2�њ��lւ���sNW��|!5nb�����E��'C��<�A��9>�����<���F�lb=ϳ�Y��(��J��5�p�1 @����V��t��r}���ב4�=�m+Ɯq�<U����

1j�?�{_74�G������n�+�<�zLd���X,C�~j��|��/0�'�bc]��R���YQ��>��/�tC�������&RI)����L�̃Na�8bNW86� �p�l�yr��y��f���Š��QRUc_�rCmGw����ɡ���� �d�y�ι0.>P��,'8i�Y��I���\��"�K��c ����ܸ~I#�����z�|�@�EsF+@%�<�D�K�����H��Kk�ȷc����S]�\�gH�#r��,ԉ�t��nr���i��FL�C�
Bm�/�p `t��- E71������3�۲�|$��ذ1n�������X�$[CI�A�$�_�§�o�v$����*�(ҟz�=��]0XU&��`�Q*��2���YZPJ��w�G���|�7�ֵ����6yY�ܣ���G�}.������a��Pc�f���3�o��;?�����%�HKܵQ?-É�]_�O��,K�ZPd��� �su�/.�W�Y��!߾�/Iu���4�]�w
�z!�^kB$n�"�cik���� ��F)��E�\���/8!I��=��n\���_�֏(r	�����ݼ%7����~DVҬ��e������ټz+��0Mb4��C(<��A����rd#SHT�g]愡��Y��}��g?b��g�+#�I�-�fB>Y'y��8o���s���9���Ϋg=U\����e͇
f�d��#E2����>�c�@	$5ϲ]`����n�)�޳��&�(x��N���|I0ô������K�KA������W�Q�x|\�A9�7���H_#G���񨏡��$�+#�$-E��Q�粬\��mP�j{wW���+��:��H�嬬/Wd�|��4�% }���t�H6i�(L�4�e�5j�i�&��ٟ>s�):�X!�q��$��+�SQD���yQ���yOw$k��n&
�"
�1pX��MÉ��b�s�{1�!C5�`,-��c��%������˗7��g{RU�&�N��k��k�1�C}����Eq�t3z��(z���ZD�3F��+'�Ǌ&�H3ox�0�@�N�\���:�2c�ƂF5�BE��dy����/�V �L��_1����p�-i�e&Q�5N�`
��1�!��t`9��ar�x�f�q���u yǬ\F�wy���W��R�&C���o�d]6j M7,峭�|�[#�Ov����*}��KD��Ϲ*n�,M��1�#���Hu촚r��%G�{FC����G�	G�8E/��W.���*{2"�@����ǲ��s�u�$5�ZR��J����A�ד$V빘VK������K���/IC��OЬ��)�1DE�mD�z!k���]�.-0�V���*��_��kWd��e��1����d��E�>��{wNO�\�6t<2���;���<r��p��g�6o����3��;B�e�HD��IҤ��xbPLɏ(5C��K��֜_P�b6bgn�+<��"�<�KV hhǄ�Pv:�����m�_G\��<@�.p�'��0�7�ߐ_x�T�V�Ŝf��,�F�ߧA؂��������a�XN��G�Y�Pe<>>f"���Ʉ,��F7'�Ժ44F>��VQKxt>p*�VW�}��:ؗeEPUݘų���W��벤��o��O��~*5�G����уVпy���#KFy���-�M����K��)�Lٺn�ƨ��+
2P��5Y{����7����7e�HWa�l��E�	����c=�985Ǳ5���P^����=ut��~gYn�~�C��N���g��<�|��)�l�NIN����03���!�9��2DaR����BA�l���;n"'��w����h)�;Bq-2�aL2�>Z�Q�p�I�dZ��]�i4�֟�-{��{�����q�Md�E
���W�r��M9Ik�Tg��S��"v-�	S�I�z�4* ]oAr�fGV�e�hx����L݂D('$���u}����l��P0�R�|�^PU��O��Ҋl�Yy��Ϥ�����X�DE6k˒�jt��˞F��z�-0`�� Y@Q�Ƴz�����p�a I�q�H���u0��5�Ԗ�V[��>&�ƚe3x^��nˊl��OP���տ�g�W�>m�I��R���]�kU��g�W�|S�)a��
�S�<6��X j3
���z�8�����wK�ƺ�N'�Y�iE�xN�Ì���i�p��z�;6�����s��x8y8#�3h�~�>�|j���η��*�������^l�M�9nP�q��;�6���ݘ0��#`��g`̐O����I�ן�@W����S���@�����ɉ����t�i.
��ppA<?'d���9Eɛ�9�t����P�j�R*�$RCѩ(te0V���#ǟVc\(Ԉ��z0�#���ý��D�n�[#N��l�Z]`�G����\_Г��\\X(KW���\:bs�g~ {;rqc���#EjP�@5�e4|NP�B�wQ>U�'��i�L5���/�!
S�Ė�-�.��'�)Q�画�Mp��N�U$�/V$�Ϡ�җ��N��PN���0���k�B�`�#?;��M.L�r�=�K&ry%'����t��z������O8M
Y����_���X�,�ժ��ҟ���@�?8��6؎#��H��?�ԓ��D�6Ӝ����<�w���OE��`vq�:l/��<�dH�x5kXn��9����b��!��j���T���9��X^3S���  �Tģ�jLR9��C�F� )�)�=��f@:��)��h�n�1@;\_;v��ϤՐ.��2Jr���tVPL]\��jq?�����ȓ՛/�f�4藮Ի}�i�0�����q�8�Id��Ŕ'�:$/�s�}�s:����jD��~aS�UF����S�]F�Q����@�O����_)d��[h�� ��>h4d��#�j�1-I��x2��_�)GG'lm��ݻzN��>B��)���P;����+D�%��}Dh����C�%�,nf������ġ����%F����&}ƢidkM�3��kg����pf_c�`�<����0�L�+<�Y�Y��f.r�db���]��'�ϙ㗑���@�kS�9��i����e������6�����d?��L+�P/TC��L����<;�5L۰�ō���@h��h�@Za8Sp��E�����ӟ�p�N���0a<�5�+=X�wD������[O�EH{wo�N���^C�\Q�4e��ݒ+j���i��(f"����������m��׿����M/ת�4�,����9<�Ija�[�#��KOG,��0���Zw2f�=��/��F<�=ٸz]�CP'���qީ�LN���"��,ݸ%i}�C5���?�4֑-�p(	)&�<�x&%E�Ig(�2��HV�\�dt�FbȚ���vК�@��/�Rv�FC�����+�t�'?�H�;��X&"�j�_(�L�,�nH��W��t�H�6;�R��!u^�y%M�<�]�6fM1	c��i���iÇ� )bit�}L�N�X*I����ښ$2u��t���S�Ok�t��� �	�'
�j�r�CF��3s�!;�g��<��p��G�LS;�1�3D](�I�m7��^N�:=A5Q_w���vY�v�JĹ�I}K
^��yo=#�� �%!"�%�k���wd��d��)X;%�6φ2�6��SE��[�eu��`Iσ�G�]h�1�>�i>C�GЕ]��>��#�j�����J�ZC��[��(����y`) dÓc�3�VDf��q/���sA��OǍv��gPmh�W��@T-�D1}�qd�y�G���9�m�D��TM�Z�≺(��tU�G��\�j����y�i�y ���@���pb��ڰ$Ή��B}k��.�5�:����I @��a����C' �/FD�]��	8�(��B��8�1/�U�ykh(�3�bT�3�,�;�鱦M=0�-j�VW)��V���G��!(�`�'V���--�4��&j̻�M)bi��nw4��98%�?
�H��r�uY^ߔ��'�\y厴�l�F����I5���ڊ:�#EB#y�o� �H��O>QTX��k���VÕ��z_?�f�	�G'֏zӞ�ƫ�ٿ���Gz�{�Ka����Z���c�&I��%ΐG�,D�2������Ɣ!�m7[�/����m����D��'ͺ���@��t#�X^���}9m��J6�h'�u���� �SS��w\����t��,V+~xp,��ݒ����P�����3�$��[�n�G����Aڤ��s9�Wi�0}��Oq��Y�1K�q�#�~�F��~�^<a]�h,�zC��*L�@R����Rg�KFiK���N2 �
���!g�����~�9@��L�H�mb%�a��Z�
F`؁�=���.s߾�=k���)��IjD�QD�(_�G�S�ᐃ1lC����k��;?R'y��Ҷ>���f)�Ƙ�����iSF��$�ي"G؅kV(x#����7�a���:�f�BxV�J�C6˽C�2i�Q��O��1��5�y�ͱ�(#�7����XӗA�M����<�¡n�=^@����4����q��s�ET8�#�)
�a\W�L/���-U�t�9����������(.��kaQ-`�6�����c`;�gY��=g} ������ؖ'�sL1z�<8t?~,~�!/F�6L����W��;	 /��9O�.��~�b=�Ü�y�>39+:xw�#ηHC������@q\\)���7�rb���g��j\�?�8=��![ˁ����ġQ ��A��Lvބ�s�Mȡ���4$wd��kk�Pn}��d���r��=�bf�"�7oȴ{�;��FG����o}����?��Tj�d)`�PĒ²4��.�wO���ըSk%b��q��ݦ�S��=3��F�����j��x� /�x]�.�84�ɘ��z�P@�(�I���*).�ו���~Eэ/G[��8���9�=L�b�������k���'�!��q�	�?�������{�����铣��l�6���t�亡��?M�b�(��60�i l���t��Ht�b��T�6sh�;V�3��[�e���K�R�P�+�� �E�(�g�&CJݢO������p�+�>�~�y�5P;�YτcG3
�;/�>�iI����g�=���P�s�*�8֗�9f~f	~����5y��e���;�9Ly93�40�p�a�+B��<�`��	3��\u]3D�H#^y�MYH��W�����/��ɤ�$���ًA� �W��˖T$_'Uüc��vD�SW#�Kа����Lh���
{ޜ�5�c���J��1���V��Ic�B��N��b��F�90+�5��@פy���k�e1p�����Gl��3�;�IZ�l$�E�a���v.�l��e6���׉�:FOy^t0��$�ƌ�
�-@���;jط����,S4ӧh�&chGO'�#[`�l�co���4q1�Hӆ�����&�H�xP@�Dޡ�jȡ*B�7��y��#J���h�6԰S���vS�\LV�1/�恈L�4@4PZs�!sK������_�o�ɟ�Wɍۯ����},����rE�dVJKk2l�0�Od��Ƚ���?yW�ԇ�k�%�֟����[�d��|��2�����C�3��pf�hoo�ŬsBO��PCa�a�K����ɑ��0��QH���;� �Ѩ"���
��fK�p��eɕ˒U*'��zmu�zQ�@���2�(���G����8,6�	�٢�xt�s:�ѧGԮ'6�,����C�߁Y�l�T Z�ӮN"Dd�VL����/����+���:�)Kq?1�o>�;^�7�����R�:�Gۓ�F�(�����ۄ]���a�D��%y��ڳ���ݟ����Vwҫ]��-�ڳHϪ��D3�S�`N��k���zC��� ��JG�z��Ri>���y�����b��:}����E�=8M:���^n�|����kG�=�W����=��ꮸ~�)��R���i}-W��nRf u��:>ZoƓ�61�q�Gv�%��h2��r��"�K4��!�p̴r�e�����k�����0���6��P:�/��u	R��4��(�J ��f�7/�aJ-1?��J��[T穯���Kh�{�M��:���A���
�������~�?@L	b��-��O�[�O���a�,�"?��d{w{F�������!q���������|�Լw5^��QO���5#<��\2 ��J��D��+�1�����MYa��[j�vICD���7�A�����l�(K�6|���y$x<w6�i�\eAߧ%?��;���>��������ȉJ�<�U��M] �@�D�'50�u�4�5R�2�����ѬzoE<���5 ����1mF�à(A�E� �X��tH�x�؀~���/[�Hw"9P�ɡ��ou8�Dfhς*��
�1�P|��5췤�/ȁ������"^�,���^� Wei�����H::"�N���K��1k����R#'eaH4�h�~��9+�+	�@h@o#]L����>���~o�� �Q$��M�FǘaѯtA�S��(F�<��!1S��a!lơQ�C�ﵼ�*���9b��75�(!�p�bCۀl͵���*�a��NH�=��(T�F�Q �'k7(���j�1�����o���#;�����XQv�A����i��6RW+�Oǲ��*��4F=�� ���]h|�˟S��#�FS�k���&9Q*P�ޖ��1�s0oY���HwVW׈��뎖}�_atQ����Xh�^R�E[��X@��J�Oٓ8j1��t��{> #��ɔs�"qW��+"���a�hD�LC�5���ՁQqL�Ǌ��A0ף�c�>���|�Zxخy<g86��zݖ:�>3�QB��\*�h3�a�Ct��\G'�|8��.�yj��h�nܠ��E���w�}W�wF��?�&�U^����T������<�:d��������:O����|��!����h����&�����H#�n_Y6K�x>�|{M��;�u�YZS��Q>�Z40�	�M1
,����=tӠ3��߸L	V�b�|�M��	�:<�M�b���q]�t_�嬬-�%�a�����}J��(�^ZZ��Ҋ"�)זeK�|m��r� Ø����)��R��儐tʶu��iõ��c�0R�i��X��9n��"ͅŒ�1��ɍѝ�FcMY���{�W���P�^���8M$���$t��K�8�W'9���9�Bœ��T�Fw��p�x�)��p�Հ�q�m��C�y��}�[�|~�._D�Ccؓk��D_�(>��?��t�Y�)'.�!����k��5����4�D��L.\�����Ѹ�����E��OS��/A,�`�q0��@�,��(���UV�~	|3� z�Wٟ ����f���=#���Y?bA�({"�?�hL��wn+<����tFl��I��r:��!�-�9���'��+0�:�U�����
P{H7tC"��k�v���QX[A���*g�P��eƠ�\�Φr�)똨<�]���#�����S�l00d��R��a���q_N۳H;6����;���\ǝI��>��f�m�Wpyg�S�W�GUW�˃(���HeX���w�u�v)5�J&?�c�c����>����=��1���$�ʬH3`f�]�Y�Ed��0~�ufl�X&S�浈��ug��y�=w�M���5��PQc��T,�/����_��//���ꍆLԘ#�*2�U/�i�4&��(Q8�`ǆ)/�������%����ooL�����B�ñ\�zMںIڃ�]��G�����t�iY���x�hW��@0sh��5�u�E��`<�����V��A��)4��B]�w��aH�����O���٬���"d�*�W�+
(+��H�R"�E蠫qը��X��̧nf�š"�KhF��F%�T�Pt�\��z�� ��LG�58n@m���%9Z�B�T3�B��dkD���x!��&d	<7 '9�����v�Q���*{���)� /ܵT���j�2.��ϔ:}�Q~&2H�E8�Ã)f�~�o�����m��-���NA_�p��d�Id�;q�'b-E|H>�f���:K��Xa.и�g5A=�˱C�#�[��P�Ǫ�[fV`�@Q����kA=g����r	̝&xI�Ŝ|���d'e�	�_f~�|FhbK��1���_��D��us3�N��ƃ.��?��ӝ�ϲ�,B`��!��hťa��p�M�&���5��YDg��M�qz#����9�πmfWܧ��k�G���Uߵ��c�gD�2JG1;af��&�Z�9oN����9b��M4b^F��f��fHK��Ȗ����Jy
�_ �N�ثЂ��bw}4�ͧ�i�Q������ɶ����l Bq�Ln�zAk3�;c�������qO��(Pqq(��� �����*��c�(+�F_�4IT�]#�:՛D����|��:��@�Щ֪ԺF���HZГ񀒮���'6j�o�9��!a��Y
sP;%4G�]����W��+�ɏ>�TV769$�2K�C�:�H�S�ۃ �1r�5��d�����˅�Oe����j���uy�'�2�Ɔ�(9^� �^
�ᅪ:����K�@�Z�+&у4'�^~M���x���,]����{
�znids��6Z��Θ#E3RJ�u�?j�.  Lk����`�h_>���#����av�9m2�-3�x�R��R��z�0O�{2���[�eq`,e]vI�L�tҗӓ=YY*J���+R�Y�]t�F(t����������~	-=/�e4�%M��k,��=/�����T1��\�)�mSOh:+$cE��p;d����H��F:9�d`�&]m�`<�7;	c�<�#�9��ǧ[>��c��p�:�&4����������K g�oee���O�~m3I�r�ɍ�j�$����
�x�j���mt!'�&�褛6�Ⱥw�O��k�+Y��N��=���8<�<�Qg
µ��Ȏ�#*>��qw{,�G�3�`���H��Te�(��̗��>/6���3�)[m�Ⱦ}`SH�3R[R^(�V����Ԧ@��qڦ~B���GQ��s�e���|��n�z����]Y]e&YhN[,p�e�Y�8�X7K��ӷJ��E��h�Ϡ��� �������q���d���ɔ~�awϧh��	��c=�`X�\�IggM6)9���p�]��x�E�c�`����XߔK��P/��p$'�L�P)��>(�A6�У\ޓ��f������E��.a!�1qH��v�R���7�yE���>�����{�%YY$�-��r� z�r�FWN	-�N_�z��\,/����ퟜI[mW�T��@��X��È0Cbǡ';CS��*k/��&'���`O����+r��;����9�{�����	�������~翑cE���4āD�y��N���"�Ȥy���Rc9�h�1�Ȣ}�  '��s�Q5��Ɖd��w�������P�����>�%������Y��+W֥TLJ�l[
E ���Aɖ���5X[���//�z��'W/�I1���y�{ah	Ij�)��8�
��
,�A��ʡZb�X��\� ����`>��ѩ:��8��Q��|6!��>��%5C�8�33xM��(�8�'�LX���M��F�{0c?��RaUL{;r�{�j}{���G���Qpz�}��?��H ./�ͯ��8���k������:�?��*bl��7��[�Ӵߑi�-��4l G�)	���B*�D.��MYQ9wfl�d�L$�ق�;gf}��DFqM".�:��,r��!-���0�㘨��b1�*欢�2��\kRr�/��/Iw~�7ޖ/~�-������wfFaK�&MDH�&Y[�F�T�V8\�İW�<f��m�ܤVa���q�[gi���q�=Ra����^?���sAq%y�il8�F���1J�y�.9/�ς�wtX��P;�Բ������q��:<�װ\��R4��T
;x���)��3����n�B[4�Ƕ,	N�fz�#g���ЙiF�ҿ���ś��Z�.[�?"J?Q'��Wn�x�LQ�r��X����$�1�9L�j}c]
z����~R�Ԡw�k�Ir��H�:�|H�F�m���pH��r�`���`�_L�I�b���i()�WmM���0�������~�w��ŋ�}���9���š�<EN!`^�xܛ��7u�A�hH*�����gr]���:�bٌ� ��6�h/_Ȓ����x�2T�sЕX�/����/�.\\V�}Y�J$��P�\�ʫ����](f�E9>�K��S]3t�����׿���U��-R�:�y��	�����3E�7D�sDȞFX�"��0�в�R�}21é��K��S(�j�&���<�.擵 1;,0�8�d0g��&�1�� z�D�RD�!q.�5��L�5�K���lŞ�j�B��I�V�R����?�C2}���5]�Da$aztuB�w45��=z��>8��Ƥ��O�����,���̚�����=g.�n׮���2jXAb�v}�Z�<Wh�<�/m�atC��/ۗvc�)�g�F02���T"CȈ��1�#4e���r]���m�}�M�3l�����6y��=���	�r��~��I󦺨a��)t�9 4g�Y��aO1����ڏ�Rs(Ғ��ћ&���zG$ʵwi" g�%�O�.�_[[U�Ґ�7o���f�}���w�����;�b"��*s;�;sщ��V���������)@��)|u�&��\�^8�8�<��F�j��Lr��5��1[�����yp4�<1�����LW��3\sM�j\�E1&pCnr���)B3��T��4��9( %�q�|)�W�}�XX�xI��]9����.�ν�ci���"`'�с�P�,�:(LaR��_��XCZ?�aG���̲��3,w�T��)7X�id�kѐ����Fxu�!���J����T�9y��ۤ0���ߗ�G��Xg5ܞR����X��%�h4��3����%Nd!P��Sg��tȏ�0�Y$5��,��rM#��m���p�Zm��i�s'��y����r��'*�n޼,�/�,W:����;���~]vv��6SY(�1�׃�ሴ��+���
��LI!:�d�����((�9�� ${	I�������F��NG��J��P�r�4�!��z��mj)�F���p��Y��kã:�>����۠D#�XV��
�{Q"F�Q���5X]SC��Dv�m��a~��_�9�i
�f� �����>E�0��?4�e��I�Dv���描�⫑dS�d]��o���#���KSw��[e�-�Ec+��V?�����A�y7F�3�B<K�����s�"f&�3�\5�؞өm:~MF}d��~�!{-R��Aށ�>k����#
NL�{y|���֨�\&�������}9E0hlD}p�r�� ��Y(
MC'��H������(����@s���!�n�|�e{�^T�T[\d���Ɯ�|�чD�H�a#�f����+�]��g,�F���{��M�`��h��H�T�6d�ْSE�(�u���.�YVl���)kH��}&e*�8���Zݦ0��AhN�T!��}J�y^�'p/pd�,p�Y}(	4Z UCݏ��\��.9�>y��,��3w:��:x��s��Sttӛ�2m�Ix��!U���=N�o��/]ɊW�Lo$�l���*��C���i���#3��C�����P�'9n���YFj��d��W��/.�x >�{W|��,)�j�)��Gm=��d����wސ�#y�(�tR��#Y�)z.��҅�����c�f�3�A*�����,�)*�J��Sc�$�F�H0�0Q"Q��;=+q��h��"8�ґ@VG���
*Rzh�?9d��yS����=ښ�D�^�Bs"�+1�0��������*�H�\������y��C��LsC��>�L��u���0t)�h��a&cF98t@�~�un&P<�|������-ǮS���@��sY{H9��&��ir�%�6��tPf�XFI#aL�h:�����h��Pi8|S?ѵu��3���퓁�產eS6���k�'�>ْ�FVE56݁F<e�+�F!�k�ܨ��3�?r^p��g4Ǌ��uNlԭ��c󄖮I7�����|dr�LiL3	�k[ztr�5�s��r��\ҽӈ�R�HS�p�!ۍ�Gv ���: +(��Lhf����ّ��F��d�8[����0����x�)����f7��hl��3�t�Q��9���8�y��00�[l
M�٨	��cm��(�˗��+S�bN;�������o��ÇJ*�B�Î\��:�~������a���Y\0!<�0l��*�E!��YMt�r���%؜�R���hUvx�F�L�Ǌ3vT1�_�q���W�%#E5#R�"���8T��T�`[(dg  �f�6�zR[ݔ���H����p��ץ�냶o�u����)ml�o��;ޓ��?���=�_��Dz�@��_����h�1?���o�ya>cW�[z�,�0�C�t���ku���K�ߦi._�"Yux��~(U}ֿ�[��9��[j?C�u�d�%��_�uK~�7�����Ǉ $J�QTZ�wM�Ȥ30wriu]ш/�D�vdii�`r<��-�9�($�2>0ZML������� �~�j��}3��x�Ո�H&��5��(�V�U>�Z�����������{���!��N2����^[�U����XX\���F�O�Ͷ�{�/�{g2肖� O�I�S�8�s�O6vq �o��a���)ua ���������J{
F`\�#���#C�՟��\{9�>9��8�#��&"���R��ȹ��zY;�o��p�ǳ@��<��6D��4ǲW�����O��p�N\��U�@,�i�tB��ɬ��t�ٽhcwm�G��2�lc�k�~���S21�����v2�B�(�b��A�y@�p���z]Ac������~O�������t�	��	�{�hG���ի���&�h{%�5�C�,D�L�@֛�ώ���q�f���>�~!�>�+��$��K�c�
�	oBԞ���i t������_�2^�tI͆<�z¯�PH�?x��:*�lQd��;rxx̋�&6R#�B�B�b1p/��;�u{���b�ǋ�޹\�R��A�V��rmQ�\��C�On��q^�eȿ�⿤��lJu^������w@�ԟ�i!D"�,5���G�]�~]��%4����}5�@�ȁ�Qe��Qd�~^�pA����tCC�*���z]h4�
 ۦ���ԩ�Gr���&|.sl�������iL�#����-asU���(ltܡq/J�T[�{FA�G�*�ZE~������}KV�ܾ-��v�=�4Vt;��]6���}]��n����a���,��T\�a&�w���x�$���� �Zt�6[]�������'�e�X,q������̰Wh�/W���FiŪ���Y��@���{��&O����p2����"9m����*��?�Pg�Y�+OvOe��LZ�g�R��F�P,Jvmn�\�~b[될�e��+��7�6rޞ�e70��1����)�y�*���z9�P��#�W�$� �P���hj4V|HFD���ʐ0k!J5�"�6D��,�5���QG�5:��kDz^�tH���)�u3&�N��R�1�Mֈg����li��;��3m霧`�2~ԝ3{ԇq⒩�HƳ\Ix!� ݚp���0.EM86�:P ƹ�
.Ĳ$e�=�V�W��y?�9���F��e�Ԟq�O.K��.��P��~������s���ӽ��q�$i����/�,��`�1pm��3)���X㟈��|�Nz>��Z���P�j�F.�r�򳳆h`򇱬$Fy!�zOd�q���)��Y]Y�q�a��
��Z[_碡"�>��D����:mζD�L�i����<�fĮY��K��"4�"n(םqbgST�Y���xh��u,�.�����/ŕU9l��v����J(���#�����Z��W7��r܂0JJr�U�9bӉg熺}ء�&-yc�tc��G����	��AYCH�L3m� �]1p�E^ǆv	�>�%I@՞4�]}f��^�Ǉ{���_jE��׾&k+���'���i���O>�\�6������Q[[�����d_V*Y:GH2$6��YY�^G@�h��������[����K��Y��`�ɶߢ����UT�P]���8Y|�,��Ӯ|��#��t�M��L��9�#D����N���A�.���T�*Tr�(c]rg�������)���7��P�aV�����~\@5,a���.�}6���4��N��܉jBF�0yF�Q����H�5d��h�F�tIF�6SHN"%��ѡ�$���Ĉ��9���g�)#��@�����Z�&�s6�4A��\0�S�%����Cf .(~�^\ 7F���LG��;�^䞏|�<ɌZ*6UaSA��cg���L�s�O�0pt�f����uS]��P�*�N��%�856'":��Xc���Lvwv� ���/���F$-C��'vf�#6Գ���J�>62�ρ��9�	DJ�B2-��_��@�щ��8_4$ug�"��<p|,"�1�|��4�-&P,����X1-���͉߇�g����XS��<<��ٯq��^�>ѯ0��J����9�'�4.!5�<x���F���lod;h]�M↉�@a��L1�����r��4�F��d�=2�'�=L�b�D_����~(����~b*c}�u���&^�0(���e�,�p胺raI~�7M��Wߒ���wd�y��d�$���k�c=��m9[�5"���CCrA_k�Z�����[R^Ө��i��Dݣ�]�|K�'w?�d�"�o�HƵ�7x�*j(�!��F�)�����,�$5,��s�ЙP�LV�GLn7���J���{E�>}����ʩaB2�%����{�|�{	��t얪�Ʉ���:�wdw�����aA��o�`����$u���=Vg�0�bn��(�^�͂b�(T�|���L���R˜��"��@���p蓘��5C[\���ˈ�B����1�����M�8fP
v5jW0z�i�b��|�Q����v��}3K9�����(4��k�<#m F�5�VMC�c4�������${r"믾!E=W�Q�{�5(t�!z#��h����#��A���T��7h�D4��P��d�A�UAY�y����̆r��P�4�9���уC_�V;���M�bҥ�����'��'�0ԑ���3�2k��]y��H���/3�2/j�{�s>P��Y��'��<e�#k�c���4$�#9�"�zjW�)���7]��O�k���9������*,�*��	(n|������Ȝ:����.15(36�VV�Mx�zq��ً<������Q�����h��#���������f���j�@=-�U$�'�Cm a��T;��P���y��Б
�!
A7����]}���\{Q��u���C#
�LڕjyA��Xv��SO�$	u�����:�tu�34�h��Ŋ��{V����D>U��?���Kqؖ�����)j��Eq�U9V��v�U��&�Y`��y�OL(E��'�X��]5��/UR^\'���?�YY��5��ե�t�t,Ǉ����<��{���P��F�@v�ȕM��T�����6�,���P��E�bFnܬ0������*�%���ԭN�D^���|aM�WE�ח���t:q�@7�[���o�<b�y 	@��������\�rY�1��(��B��$� �&:��t�+�_�7��e������r��#�S>[��D��$����d�р�q:����{;��Rc�<v�	c#J
�9��^+S�r}�pAǩ>����p���)�aߗ4��;��h����C��!�zO�"k�#���E����������D��� ��|A#�UYP	m�luQF�C�LJ���o�탘: � z�� ��C����YN_2�*5�,L"�I��D��8��������o���^�8��R> �6j���h*���a���sb)��&<�	��Gݓ���~_�oU�����_�Ap��u�׎��	ʋ�҄��R��h��@�g� �3(�m6�GC�&�=xZ#Tq_U�Ey�$��3����>�{�:��a����Şh������DVM�ABG/��\�"��*�dP�O#O�ǆ�l69���bc!����3ӽ�Չ�"�޳.��qA/N"#�������ht�wrJ-j��1 ���}��ݸ(IR3^CW΂�t�D�йB���εZ�*�5b���ɖ�����T�a,Dcɸ��\��o�&[�	%Н
=��q��pD�r���j� �4p��������撼��D���;?�j%W[7���5����������Ka��z�lU�+�G�l]�*b���o�{��Һ�3k���n,��u��y��̉�^�6JY`X�F�m�ĎN[T~L���^�v饠��KR?��+�п7[ +�}&��e���E<�E_� G��Gʰ�}�����ץ��$��*����23�U�%��	eA��@sH�vz�VϜ+"O4� m2H4=g`a,���Y��]��B������3t�3��6���#6���L�&�".tj�籮1q!>��G��v���hN���
�����:Y�Dd���!(��"�8���eg\��6l�AM4,����z7m��Qt���D6�53<�M�;T��l����u�3m��.{Pfr��u��R�3N|��<�w���{�b���S��CƤ+����?��]�|��}}uM*e�q���L���;�}�3O��y{?�y���@��]e/��b�ǹ=�JĖ��~�B���ߝ3����c�\ޒ�ZnC�T�c��8�:����qr�Y��+5ӽCS���UCu||���i��-%-�ȉe��4>PG;itZPX��%�Ԙ��%̖����*q�T})�-�-h���6����
)������M���Ht���\3òqڐ?�����_�k.Hs�U=��\u�����Oz�t03_�_��"B��V
���j�3r�ʎ������ZE~��o��ʦ��@:�6�`� &P������!$��ЫE���e�
H�!��~O���R�K!G�Hr պ�\�^�a����JFE*���r�g�g2V����~��^9��:�#��h�V-Ky��YEn)�v�!�(j/a\�>�����a
�{C�	X
��3GMo�nрc�-Y ���d3�My��O��,'�Mv�A�h��4�~:�"�zfhK2��r�i�7�)0	פO��#�Z��i�tNm�>p杺�(����5�^�ǞIit� ���C+1<���St�ꛔ5BbD#_K�7H<�xbSLs&�&����e�H<$�� E�`$~WѮ~�'�,�Wd��<u�PBD��#�@@뾞C��&��BF�ǿC��v�o5�B�9>��rbz��i�c0�t�{!�l�5�f�ӧjw*++r��,(P*+P��gwr�l�>��B�` ��+t\p��1�!�Ծ%k|����d[_�i��zn�HQ��X����X{=&)�铙��%�Vs&�8?�զ�M�5� %�Y���u������}.�+q�̇1������!�GѬ���
�1�vl��ܠMZ����W����<���6��4)���9���㎃AL�H?����y����3��IZoJE_o(��]��瘔M���5X{v�1��v�u��*��Z,$�Y��kh�������eY#'���H�_=IKا�q��wyn�L;�u�������}dS������@z�z��e��}�����YG����B��gG*D���P�F�5d�MK>)r�ɤ������Rt�\��.;Q�I�;Ҩ��b������"��^�Y�NĎ�B�b���|v�ҢT*��\˒p��a򹘿�&=N�ۢM!$�h;�A��x�Z,#(p�Q��=~�%{��v������*4:�)�(r�v�Zvy�&�����4�!YK���AĖ�������%ˮ�vD\o�����2��|�"�ݤ�&���@_ �� @h��h���� �3Q�7���=�l��??��ES�U=���{��q��s��WU�O*��e��k"N����{���X��p)|��{s�Q�����9c�=q2w�#�si��%�QS��>��4��h8Y "�W�/,�U4bD[&pc�3��q�R���$%�Uo\Z�iB3v��8B��y�4.\���K@�Q���zNQ3��<�(�<�����!���3DN_�B��,4#9b��Ы��$(Y�`\�����J��///���2{"�*z1U������p|����ٓ-D�kP�M��bH��[��&K��F���c浳���6�}��ϯ��Շ���|�%�Jo�W��D�s|J�D�Yk���� ���c� B�� 3kQm&�/�����9B��������pg
�i�M�{$t)�

%�M#�Q�'L�Z^^�Do�	�"s"V�n��Ċ ʛ,T5��R,��݄��o,��,C��v�����LI�,-.��M�j�<����D��#k/��g�{�q���"��pn����V�`i~����$ں�ң1�ݸ	�/]�N���i���~�cN�>n��������Aep�	���3X�[@#߀���BǪ���)�.T�ܸ�0lC�k�����|�>���!"��}��!VS��*U\L++�o3��>�i#���=���3|�!#�$n
Μ�߯�X6�6�������x��5Ō��EX]^���SDa1� ��9V��:��B�.s}�k����)}�-P����B!=2�\l�'��I��Y��#."�y�2ǩc�@!�B6��X4?:l��C�J����wd�����l�X��h4X�mLDҵ)	J�yM9+���G�z��c4�̎Iu#�͆�h���"Q�6�dХ�C#����OZ0���#ES����@����{���L�S�s80B��r��F��4@�㶯���ky�&�\`��u7��l�[4����M��I���Ӛ���Q������EHj�W��D�:���7�$�5�o���:3�.o\�ãCsڨ�>݄?� �67=�����,���{���7_�o}�8Y"��Y��)�|n��_�-�νn�޻�Z����{�
�j;�%�܅�H�y�~[f{���>f�s����"(~M��ta˫+���Xd,(CO�LrY�x�Wp����
M .$�3����S��ه�e4|T�ԦJF����X�9��8�4Q���WpA�"��̈d:���&�_�څ����Ξ<�4��
G�P@~���"j�`IW�0���#��8?�����K1�� >��u;�k��^�/�|�3�p�ctB���%�X_�
���#6\%D���Ub�0?K�
m>�Ý�p����]V]�WKp��GbT��]v�Π�s�r��&I*"�'�8$�ed�c-C��\bQ7������C�db�X����P�k��/�1a����xOZ����?�q�'��%�鈹�=��XI�$�MnлD�3b~����X�	��T�9��k3vnc�	j/h!R�({��-��O*9@�E���<��C�
�h�?���I���SQ 	M1s�1%����TvZ��h�)l0,����J�i�͠�p�<#b޷p����p}�F}��4�p�>��}*II�i �ey)�Q��σ~$�A�����K�G�C0q����(�fgau}�=:B��ژi�=�uN�ɍ*
�$�����3��o+jm�W7`��!��>��%��F�H ky�A(�-���NƞP�~�G����S�hJ^��V��\��Ype�9r�����0a=�8;�־|�$M��9O���g|�aqqk��&v��7�Icm2��#<�H��6�.��I2�St�I��v��X��Q'#W��Rݥ"���X�i�Ttu�}|����"bOI�'�"2Y��T�\/�1�;ȄZϹ��#�̡�Q�qp���5b��_Q�
��`����:)��^k��S���,�U�,��8�ϭ�&�h���H��"0^'M���n�)^����h\�ʅ2}���"����]H��C$Nr��i� K�R������E���6�0�.������ݟ@�}Ɖ�ǫ�������6"�wH�fb��"�e��\�Pʦ�4E�	�n�w>�w�8�5J/fB�\uI���Tzt����T�*^�~G39H̪ި1�J[�0��da&�1��ΑZ6���"�(��Fd�I8����X���~C.l�|M=;O�H��Ucj?���n�Wj�1m����^�D���9�����D�Ї:�C���llx�3�]`ܝ詗T*����O��谾�h������#V�	��Ý�x���"'ށ�����Dg�S4�	���n"e,,-1�az1U���p��݉�v<��vڢ�<R�,����a�~Ϸ4SA� Ta@����[ �*%�l��8	��E����p��J���t>�}���#<�_��o��_���@7�c���Q��[�?��MӶ�v�/�ӧ��R7Pw��[�tV��\nQ��mi��ъ%���2�WCA;p�'�cR�|=%�c�j��ł�]E#@\y�[S�l]����W�r�}�F�jAO�~�i���A���-Y4�Ø����ؘ_�z��|_.H�6ZG6�Rs&��KL�C�Bm�=X�W!..B�s�-�Q��<�����F}��˜,&o�L��8��93�.����z�F)k�4f���U�^��"��S\�M������a�볆�7f��0u,�4�jč7y�(cf���B~==����It��S<�5�' ���Rh�S��gO��(-�1��9�cM���_T��l���� ����DǸ��=�4��/*��X��I�z�Q�+�e�)��:���7�@_\�JIQb��0��Lrl�ao�V��z����J�&Ml�P��P{��y��c`03�@bm0��^���,�A��F�̗ekk91���D��^�xraC��!/Hx%"1�%��"C.�Sk�(%Y6�!2O���y�L���T�@�%S�j(.�w��(�ū/£�87F�f���g�����UX][���@�U�b�jTSx�կ�������t.FK�Z
5|��!�O*�������t��#4ڟ�����}-<�f;�羘�kfr��4й� ,�t��=k����3]l��<֍�9/@np��#��..�eB��$Z\ݣ�4u���%���#v[+UҀKa��%XD���kId(�Y�ʟ[�ٞ��ie�����,�'%[�4? ���lb\ ���̣=s͍��>89�~
Y;U��'r�ګܣ������p��bny���ˈH�89Wpa�ll�T#����.�b540�T]�{�>��l>~'�.\�������q��X����s�V:2���q��I���L��6�(�B�@{���l��n_���Q��O�3KPG�D
{$-<���=��5�e~�B!����NxC 5N."���R$�՗bV&���L*:��|c���&��`r���<~�ľ�h�<V�<�b���p<2��z/C�u���O��Iڐ����梨,(��Jc2��2����x 3�4��q�=c#�pn!����7��|Mt�9�%ߩ�v=�zJ��p���;*bgГ�^T�
�X(��z:̮���T&D±���v�h8�Sb� 88>9����d��ȫ�os��� :��$�š㕯��|���?�C���8�S1�L ��H����[^
�y�V���S�����3���������ʤ������UWV���Xc��=lQd��بƢ��.��	��"i�7و�TʉaQ*7n6�pR�k���+��Z������ⓉB@�P��f>K*ۂG,Rk�Ly�$}��[�x*��4������� B����Op��VV����Cܤp�7���G��Z��k03��r�B��F�C�pR�sG�(�'�M��$S�
W:g-��ڬɱqqn�t���ܺ�	�yeDF�I�l����7�1�'L}X�^�L>�h�r���V{�F���$1]���Κj��V-�Ѡ/A�1��\���TFc~~6�U^։"`�뤈��6�:)�E��+��?��w�tq#ui��qci�����͖��6bi�V�3�O!�H=�X���G�&Qq2���}8eo��U����������uE �c� ��ZYs����D^�D��$�7�nL2�ȅX�zQ"9���N�KMyv�cC���P�BC�J��&,d3Һv��(GR5�t��.P��	� h�@��} ��@�\�8�i	ўQ���,h:�0���cn�'��h�'�)�݌s/^����߁���{���蓹X?��n�ON������[o��kׅ�����"��{B�Rk}�C��ժ묘�}З�ۗ9���R�HqO*a�;\�-�P#�.7b��X^#��
5��1�0�M���9D!1,�Vq�����|���>,D(cNP���I(�\A�N��9�1w�!"�Q���Ȍ�\S|���E�ƙ�%f�"��t�	H�g�t���������A?���%lu�:\~�m��%qq%���Jy�m���"��I�α�}�NB��p�^5��{��:�������qc� �+{z��>7����b0�6ܙ�k�L�������H�4�/3�ʡ�/�T��D���#{��-&���H�Q�h��E�O�du�$�r2�l�$>kq"�jU*�&tz� έ��b̪���|��f�0��� ��/V�Dĳ!�4%��Á�^bu�gAV�=��0�y�ҩ��|={�F<��kƥܨ�ZN�ˍ�}f�pϏr�l��qsmR5&%���w����8�$� )n����!k��^U���p���ճך�T���.)�W1`�2�4X'3������*�>���z�Iʒ�̚��H"3j��v�����m~�����{�zp�IH��-�4����?uZ��*ܹK�Ŕ��1��-��4��C6�͗�3�>}LT��?﹡L��t}�0��Ӱ��U�S��'ᤈ$�h����"�|�Xp�����*h HnuK�=��Y��nUDrg�iG�ѥ�w�]PC�����ܒmV+`�n~�Ɖ��%�R�⋵�Z�����;uy���7St�g�.�߆GTE�;��<P37n��/0�$tZ��R��^���&�"&�2�$�N���7
�S��>���mB�V���̯\�*"9��]ٸ��֣� �8.b���C��+l����*gm��s F���Ǒ�+b����\�ڜQ|�X�dWc�g%ObבD1�dg��(4R�Uh�k��r�)�Mxr��&�X�����~��ME������zJaA�`7�/���f���P

��-��v�^m�2 QR�/��uA~'�����e�m�����hǬ���m�g���2X�t*��d�f��J5h�E~�(ǴFI!Ѫ�#Xc	ő��s���i�J7k�n�B�%���؃!��T��d���85�"��N�<!��u8�(���mxqc	�_��!�?�El�%��i�#���P��_�u���1�XQ�=↴ڐO�ޜ�?�Ꮨ��˿��|�&�n~�lH�/�夐̞�B;���t�v���A���"E�&�x=Z�+CNw�L4ų��p�:�c|MJ���V��l�А�s�eQģ��76��R��^k ]*^$h�h�+8����=�,FQEf���Ĺ���qA6b�ȫ����6��q�.��Y@0��iOG�h���,�&T[�W*u)���o�nR��l�b����C(�#x������=8;��k���Dh��^�uhVL���F}��L-4��f�	t��u`��vqӨ�$u�J)�U�A6L���Й!EA���ʱA~�H���h�@g�h؋c	h��-8>�ay)!UeV�h���r�TJ ��)2�",��K��w�uS����m��Rej+�@��QX���3K��7趩��I9�H%�X�',��A�U
"�ڣ
`j��|�X�L	��<}/�D�����E�oBK�ӈA�:�í�pq�
\]Y�6n�~��(���%QFUF'�f$��T��f�m[j��\o��ĩފy8��#�E&!�x�k!֢@��\�7ځ��S`u�X���o�.�����w簋�,Y:����w�w�wyN���@*NO[�я~W�^��+�u:R��<�*e�AAAջ7�g9�	��7VC}��&�s��#'�/|�y��������u�6>(�R�"�U24��k�8�H["��$���XQ���I�J.#�X�x�|eyf��Z����� v�Y}��w���u�����0Dn+AZ�p� �f�,�ȏQH���Ԅ�k%�������1λ�X�l0n�eD�!>1Q
IK�� �ژ�7��Xi�Q���c��Ғ�`q���=4|]��J�)b|i�P8�$��@q�C�(<8b�@�р�8�{Op����tk�	�
��A�\�B��h��j��&=8��m36o*���Q����i�+G�4V\yH�6f�;���a'o�X䙑�٠{��1���n������� ��sk}ǎw�M3tΑa㍂6.�w�YLpO>�9�ʨ�V87AmI+��UP�n�e��O1br�q��#�؉���ʏN
� |H����/z1@$�i'��7EzN=���}X�ϸ~�
��.��>tF�t�#@з�� �\��:5�.�5W��kF�i�Mǝ�C��Y��*3����f%���3^��jI<�tP���gI�ϓ��P�|��2����q��=�
_I}c��%Y� �?�||�0��4������g$%f7�Yu6�"����bM�t"ŀAA�b�̪T0�K*D$�w)=��h{�[�w�J5��e�2i�)�G�ɠ	��sh渳���>3���ϱ���^ �P+&PF�����\�����`}��ܼo��B\����	���pL��Ɉ�b;<ß�����@���
7��GR|Cv���(�K���J��4,OZA�.�rc�m�
�\w�"�C�t���L��
X��/�aԃ*��Q� 'vQ��Y��*�*L�:8n1C���^-s�Aif1�"����?8���c��d�*jM�$|]sn�]�R�|Q�f��L+�tZ��!�CcCe�1H�Jzb�c���<�fό��O�%#��Q���gZH�~�PG0�_�����=�����^� Ҳ|�^���H{�:��9�[@.2rB�n�[$��} �)QU�1ڈ>R�Qt�y�В7%ZS��0�x�OBF&�A�7�4��p��L��!���X������*�]��\}O�I3�����7�����5�i�~�vǣ<�př��L�f�ބ�1k��ZR�eDz��\�	5�1�P�2P����.T�^���K�Y��d�������D�WJ�)v���}=~�	�8ί/�Ϧ�1�@>���\�v���JO�)�B���&N���N=9��cϓ�Ц��]�/w|���0�X�5��{�=T�8��H�b�%$�R��δ�%CtN�А'D�b���I8�J�#b>�xB���>3�(�R������`%�\i#:x��;h�6�۰s���	��r:YN�z���'�R�'1Q�_�F#�j'��k��  �;�f�m�]$�Bv���3��$Da�;���{ոׁ�����SH���d���s�,s@��;ã�-x��!TJFp$�D��dԥ���Z)R�%�����1z#���H 7Gj�G�VJ�o�2�DB�1�1q��pA3d/�y��#kh�G~��B��9	8INŦO4U,£����#s&3��02ßo�� �v2��� ����X�����̯Q�D��bj�jG5�.��yTE���X�Q�$6�7�q^���0�*։��Fun:�߇���EQ5�X��d	
S��J0�t_��i���I�4�k�Ӌ&���N��b&^B�*O)vt��)���@ca��Wa����{�����o�����U,	o�ƀqj���R�[
f�b�$ ���5��c��ϧYᝡ���M���#ц���U�_2I���?���=V/��?Oվl�ւ�]g��ʴ��f�}�x�1�L͟���գ�� �����i�qXCMR9hz��CRmԲ�ig�]h��?�qP��B!����x<bEƴfr"��љ���n*Mɠ:	����{���#�<h��i���)uQ�v`�}ƅ$��S�HD)�I@&�(��Z$�Kʑ���O�E�Q
�xx1L�%F�R#c�(�d�3��g��LL}����:z���x�9�.i��7G��Q',����#�����=Dj�֦*SJ��1x%�Xh��<��)��x�4�BZ�Œx*I��'���Y�yY���h�e�e���ϑ�H�!N��������R�E*:-Z��V�ya��#�k��ԯ�`���Y��5����5�z3�5�`C���m�j��2�E놸�{�ϟT�3Dl#��-E�R�m��n���w�œ�=p�P�)�4-o�YO�� 3OD��Ďtj|���޿<�:B�t�8��}��Np<$���S��֕_�E���M�/����,6a��%h4KTچ��x���</��0'Y	�+�ʼHL�D���o�?����rx��Pl�c��G��o�W�^�d�%K�&�r>��P��9�4�1vC$F|6�yk��1>?�>}!�G���B3�T/���1}��y�"Ay���d��HG��+�X��p��+PN��>���1��)��d't/��C(��+!�+�y4�jpy�
Wg˰ut��nWѰ�/������Z�٠�΀{U��y��EY�1��n���t�+�b�J�XtJ ��<�-!G��S�4E��2�=��xz�ܴ�HS�zђ�:��rqb��	�PC�	�K� QB�sb�V̥�$^E��)e̝��C�M�
S�d4JQ�}U���&�����!�����sy����S��pǠH(��:.��k�@&�F9S�)z�0�Ω��ϓd��b2��5�n�C�r����(\�_S��xj��
o�4�y�~Q��ރ��,8�O��5�ۢ�#�_�k"��qz��+r�z����lDU8�,����Ǿ���k�_l��V�;���6�q�)~,�Vs�H��v��ұ�	���������v�c���\�?�ז��y]o��]��`�A�d/�c�( `O��W&��(�X�;���K�0?/^��E����ݻ�ݾK�QReq����) ཈�D!�'R��ĥ%��EvY?����i���nf�;ݳF��0L����:���IɭY-p����ᄐE6a/z���"��0e�O��8��:Q 3�OJ�l�z)#࢓dU�Cs�
KuJ,qLz��f����$8lu�?���6��~9Vl�������2�Vh��ה�Ѯ�=X�K��N����3\��gN��泽�g�?���&4�g�3"jZ�Å8��!���H�k0J�JZ~N�Cp���K1N�������h�W�[	s��TTF^�;b[;�Z���݉���T	�wq)�ƙ_�f3$1����{�5n �l*��e�$�����p�u�OV*+�B���l+��3g�r���t`�}_��"\.t߬o)5��u1d�!x�����s��R�FYI�%�qS���:aϫ\-B7���XZ�G��+����S�W0�b!�L%,���"�}<�����k?X'1~�^�ĸS�5�8F$������}�Nv�����O�|��q�s<��*��G�p����2fV��ԨT��A����G��\l�ґj������:~>�bҐT���K���C�^O��"��߾,����sl���u����1m�E8՜����><��8�h�<��d��H�{D�{屸��mgH;(��
(��rV�-&Aי�g��Q����kʥ�C�ʦ 8��bҹ>1�g�0�cX���V�M���d� ��ggJ0hT�:��]4��!�lw`�����Tp4T�X�bXÔq/7}3'���s\�'�M�$�_�ssp4���c��m�:h��ڨ:֦�2��&�9T��H�5��i4ΫFE�4���� �����6��Ɔh�O�kTP4��q�UD|e�?�ۍb�ƛ�x��h�of�m��|S�.
�#��I���E%�͞���ؽV�8h#J&���<넀����!����'��aE��>;�%_dX��!$$���wq�Q���/
��1Tȡi�LU�w����P��ކAR�q��?y�i,�-��󈆅֣������"�8���3n�x%f�Xq�@i�;U9��@g{��t�*�p#i;��h�$\�L� 	��,ȃ�|�*�_����D�Ho���|s�{&���uvt kh���Ĭ�#�t�r<� N!�FO�~�ѰS�e:�gl>���~yq�����Jr�EBy�!��(\����i��3M��Ɔ�3��}�B�!�"7�A��>����&�ԩ�v�߸
w�|�;>��A��(ۀ��{�LwO��S9]�� ���N�hM65D�,�5�JA�JNVq�P�'|��7��7��2��~��]��Nt�ō�C�1��CܸN�e��"�\����cƤ�8�JB��1loA��'8��C1-_,p�jy��3�;�L��h������%��0�����α�es���1�ZC� 	3:�.vZ��rե$?L��Pk7�0d(�+1��M$�� �$�h��s��X��t����=���γ��KX�;!�D�$���[���D�0L(�ʮ����8�HZ��볘���1��*����Q)�Jm��n���y�0��!�����W���p�h:��-���9ǃ�{dDכx��������Q3�P�4g��j��)��a)q�����㻰���޿��+z��p�?���7!��U:)d�B����k��W���A�����;ԪPx�-��;�@mvN����W?�;_�%d��i�����g�f�_��_����m��1f^z:�$������7=J��L?f6Ҍz���s(M/�/:�K`�;B�>��p#��hT�ֻ��.���vP#���nyu�;2'��$J=}�;��F��<^*IR�n0�h�'1�k�&Y��Si[f��"E�`H��Q�T(X��y��+2�"w�:,���{����q��Q-��Zop�;(����.�����Nx��Y��ƈ��>>s�`G�o#Z���Gۃt��E�<���3?R���$�a"�p&xҁ��%)4Q(2dq�H�;�Ц�Ɯ��m�t����T�&�-���+y%�\*���*�)��b&ݨ��ɕo�����X��&�l����:2	 _P��?6��$�ϲ�1G@����J^H������!�q_~�4 
Ɯ?O7 ;#��r�v��%sW��e\�T���֊�4<�| �!ژ��bи��Ĩ߅A���)7�.�ݙ9�EB��h�;8_��:���̲���*�O[�|�w��]D��\WB�רZ��O>������]��(��C�so߅rako�9��2N���B+�9kW�������bN7w�Xoy�\x�e����0s�2l�Z��씼Ej���n"T��(�4���j�H���g��_�xj������p��i�wB�;�P�椠�W�6�(=_���$�7]{���<'~������v����s2?���t���?@�w�a�*�|ۭI�`���[7au�	����c��d�����8^�����S�F�D��e}	먨P���Q��.����jMl���q�+�T��!i��&��;f��4�x�.�AM�W?z|#r�֡K�H�;��\|�3��������$�vv{'����ĝ�٠���X��h�Cѹ�M�����g��j�DT/�=PccR�C�$N�q�{PP#���`r�2/�U��2ͨ�{'v3���A>#�DP�;�ĺ���o������ց�����2�mN��Y,�挋s�Hӥ���@0�,�f+56=�,ߘ�n`�^���S6 �y%�k��\���	��J�SOa��VnQ�۵�98:9���=��]�ه=�:�zx��1x(�ᴈ�;f	��&cO�.���>E�ݝm����tG{,��MU)B���QVq�t�g0:>���3�ty�V֘ZKM]�z�Fqc�]���i���`��M8��e%�j��K+כ�x�N�W*8
�2�t>ڌsR8'F�c�I�{ڐ��Z$���$팶b~~666����<7C���w�P���x��w�|�{*o4�B�!�� �M0�q�z��i�.�	�/>�y�Ǎm1F�H�'g����(�(q���AC4Q�W�$0�Ẏ��p`�HuRC^o2���z &�%�bIՄ��X'񴄜�;J��QIu�m묿��'
�/P��x�	�1#��Hq^{�U��7^�?�������38�����h#��;9p�pM��N�O��(e+�"���;��Yǅ��`o�|�dnT����>����;wsq�T��>�0xg���.�0�U1�����v�Јe�`ĩ��4��$,��u��p�)�u�a����vo�����&�U�g�p*�y�\U�~�|Y9�R{f�3l,��b'#vf��tqRƟOq�x�Q$Y�GMOl��<�BWd����JCB�+HM��Ts��H�*��T�)A��Lԁ�B8�6.\�kׯ�G�>�D����t�C����H�qd�i\��0���X������:N�����F���]B}<#�+Sw�oC���L���z���.]���T��Ml�Z���p�f`}u��г!8K�' z��ӴB�w�X��(�F��j)|���M�Ƚ(�d�Δ��gW�>z�!G��9U��?uk{7��L��>���JF�vC�ˋ�Q�R�gM�w͞�����*��St�+������Ch���c�wB~h���{Ov����}h�1k*��T�6��RG�A�'����&��v��E�7tf�s3s��*�U�Q�-H�G�JE�:V��H�-��i|�,��Y�b#M�e�3�9bc%�i�ls3X�_��Fʻ{k�c��_�*�Ư�&�o�����?���w��������gP�Yf��nF-�T�J#V������}��^"��25�=�� ���"5C�' �|2E�B4}�<��r�L�V�?��g���q�ǠWN�I���� �T���ON�g� �g��N׼�)���MA��$d�s��a���e@���|.ٞ/a��9oj�B�K^�g�;�"~9_}�6���cF��X��K�U6X�QN7	����^�\<	w��S1�m�����`yu	���*%c��xm�m4�'-����`"�5��c@tD�o��^��=�H��=kE�#XAAP�>�L���p��)�]޾���Up��� Je�i܂��6`~f�&ϧ�I×1Ks;��yMJXN�<�E��ֹ�B��3 �{�.//���:�#?��RJFS�1
��sQޓ�z.��#E]9s�ץ�f
y��I(Nt�s&�՟���=2-cȈ�ݏ�!�'�k>���7) ��F�������C8��,�����'��!���
`3b�x|5����Y2@$)��Ԋ�R�L9�1W���L�A),�X%QJ�鋒���⛊#Ὓk.���R|w�h���bi�Lɪ��)�.��7�y��_�<����}����k���\�q��襀ȅ\�"�n��?���}��\2	M	jΏ0�'�%��j�^iQ�p��1��|u����M�QkDS=��b,�W���-wbJ�<ҹ�� @�l�8I}��h��k�h�y���|`��,ߛ�L�|�O��4��{ޯ��/y��}i�Ċ��Z�(��s�?�z�;�&��CH,'�^�+}Ũ��Ǫ�%�nHyR�?'���;/D�5�Aa� �*
�#���s��P'1�V6q���/@eaN{C8:jqӓ��m8�?��j1����@#Qf�$�#�lM���	�d2��N ��C�l �Y�ø��9%k�U�:�+R��cyp�*��S3�"Qd�)	�}�Iח�PK`�A���b*��d&9��3�<Q�6{���:�h!�^P��� af�Q�����C7 �F]6�̉mh>#"ߤ�'O�\��y��e�/j���T�9%G#F���3x�s;{�pxt
��}5�����$��rF]p�޸*����~s�pREۂ�I��>��\�3�Qrprr���|r+�D�BB���F���0�BH��ƒ�`�R�.M$�+\�"����Ϭ�p�Σ���7��勰t�>^_[�>��h���=H���ef~�4�ń��n��vAb۴���̞s_bC��L�+b���J5�hU���e<�ǝǙQ�ӪTEpIupq����w/~�B����Ξ�Ys��yQ��`���4ϑ�D�u���X�&�s�I��X7�HC/sL��(=��3.vӰ�_���WlE>&���%�q�<�X�C����D�{≩�D|q�xLj�T���uz|̍��n�;�n<�n���,T�p㭷!��O���:�Np��8_K�J��%�x��$����"�P�&��8��2
+fぜ7�(����K�����m�(v��	w�B�΍��k!Q>t������9��W`3���J��O���I�^;����I�j��^���ט����u�Q0WXuV���G�^V�9$���:��Y0_8�O�?����L�[��ǿ���殇���������z+S�I2�]�}�ހ�S�aI!��]�阯�"Z���k9U�=����$�K�Q��*T�U��,���S���'�d�e��F�T+��̈�(��!�$�H��3U����X!��E�KL�^�?�����Tv?S��;��:��{����ܘ�A��-D/�G�>؅^c�s���)���	0�`)	��f�u����F߳p��|BG�Qҕ/>	�GC�S�3O�/�{\�! ��g�'$͓B!�]dL��b������3�Ӕ��O%�:�.���RQ�(W�K�D>���a�J�>�o�J�!�!�7,�9|�ܑp���S(���}J��DcH�8��ˮ��{dF)f �W�rp��z�e螴��������������4�U�^`���;T����b��U�맰I]�ba���2�"�n4��կ���8==���� Q~ڭSI�R� ����4T!�Fm����XbԜ��{�@)+V9~�+�2�80�귅*,.2߻��#8nT���׿�rJlAX��fx$w���5L�I7/�Ai$���F�ͷބ��Ǫy�@��?�;;�Y%����`�Q��+Ѿ�vx�7��������-�6����a����2,bN�cᄖ�m��-�I
� �K��LE�2�KgИ�{���,�/�a���.ofL]c
b�9�e��D�rZ���c-����Wn0��Ѝ��$���/=>jC�}s��n\���|����C�1o���Jt<��ɡ/	�+�i8#@p��@6�,��n�@
vL�S:�"g���ĺ"����[����l,@�%�N5�0�z0q����/EB��+[#8��;mh&��N�k;�p�Ak.����ڿ��^��֍��.c^@n�%�u��󻗪91w ��ɣ��A�3U͓)���qZ9�qBԼ����m�!�Y����5��`��2Ã��s��|�P�����c$ϵ���1"yt�an���%�+9;��S�*eW._ X^ @`r�W�(-�Ba� �v�sq�xP�'aws�%/f�:��Rc�.�n�2	#�\q��Pe�(e��r_�(!��$o$MHƑ�?��<:�)~�6A�w���k�2�&�����\��'!"l�t�Z��ҋ/�� �(CYf��tnP�%��"�躙�}pA.]�zc�<Z_.��y�~�>7�������i.Z� ՄE�]] 8nV��D��	�N4�(j"a���B�+J�j��UeB4���b�"�l�(�ދ({�F��:�a��b�F!���3(�'�>`u	ݼ�<��k4,iYr�Qj�$N�����4�y���K�S"E��&�YH���k��k���{������|���k�k�@�p��� ��ǜGF��̏��Y�u�����+.�qC�+G��IW� L���+�J'~��{D1ʒ&��M����cbE�\��>��eȌ� � #�iA��ȇ"���{���SP"
�����w�I�S����P�O��ñ\Oʄ�*w�Ű���-Қ�̐���B#o���2��S�(n�A�R���h��q9?!�!W�f,WA��V�55�Y�ON!;�0�F��W_�_�� ?�v����փ�/]�ٍ�^J/.�=�F�5bL�ۈ�k�87��[�j9��z�h`;h�O���N�t�	�'PkԘ������X�����Ǿ%�$�n�31�x6�d��=�������+�`}m����;n�RV#���������y���9K�
�$�<N�D��l�t����:�$0��g}u���䒟��`?��~�cz��36�L��5 ���1����j Ƒz���ۢ�jg��,�]D7��p�Ў�f�\��$�W�I�StD,Fܽ��V�avy��hܛ�N�h�Ũ���rp�B u�T%9�4>���h��+l\q�"��c���tK\$D�ျ�\�p^y�E���d"���D���-�ėsXC`1by�d{��=3kF;Un�r�*&���Ľs��i�N���T�&Q�͙b��%s�Q�s��q�a�p@6�\b�#0��	(��WGG��7vz-�����-��[��A�3
$��u��=ۜ3��ۘ֘j>G�!4{��_��pr��˫S�~S���ɀ��\�W`ia�V�^�]����p�ɒT !��a�}�+��Ak���_}f�.��O�_ͅ�H哤>���sQ]4���z��#�ٚTf���0CT�RV��a�#�߇��1<�|;���3B��|8D�_K��ĨX��ʬ�3�UJ��[��p��w��k���������
Go��L2%�\�W�<�.(;������畚�p��V��(fN���p��%(V�^vc2c3zҮZ1��|(��xy��f1�`�|���F�����A�K��@dDKh4�p�nԪp���U)�)��]�8PnB�9�N���ܰ�:��I��奤a	���!��=8h�!�2b�dM���b�]�Nʤ0b�Br����`Y*y���N�ˋ��"���	y�8�KH��<��^]Z�|(�*�L
�2''S5�:�m��'S�K���S] ���5���i>�ִ���X����#�|�2w�P��P�s8��`�gE��,� �ڹ�"$k�{�A Ӑ�SdO�c��q9�S�A�A?��A�ɢ���Y6�"i4��#��<ñ��'�<R�n����5tl�&�g-���+_��C���l�2���;��6��rw�xӘ'�B-���7�`� ��va��<ǝ!���_�o�$�ٱH0k
���_C	�TT�ه,9��_�G��Ɠ��E88܅�nf�����^����!M$9�>>�O~����=�3�is8
�0��ٰ�	��L8�����.{�$)2D E�ԁK�e�&�|#�6�q��Z�Rb����#�yw�_GS�t��ܽ.^dC��䉟�.��S�r1N�5R���3�{��GC#�?�~�?�Y���Ǵ�������vו�XZ<�]D⬮B��ʢ���'��p�2"�����8�|���k�F]�=jS��*!�� �ԭ��N�!�a]J�~��TN�������O�ڪO���l��r��Lu�L��]�,`��J)�DO�0����|�[߆;�w�����-�Fդ'c�a�/�{��H��͈zM�<=�Wl���:��{>���>&]O�y0@/ǽ�:�ѹ�sY����N~��i~N���	��yZ�631�b�#��힑⨗�d��\�zLf?���a"ɛ�l�ؙ�Q��ƪo^��CO�p{:�H�(ׂP�Ҽ$ު�Ef@���8������6��	��5�I¹R�Xm��ǧg0���]��=�&6J	ܽ�ܹ�14�P�������Аך3L�dhƵ	�Aw̺4��n߁��w�QA�a�	���x�[� �/� ^��ύ�^���Q�c���aO���Hf���^�;���~Ey�A��W���~�'p��*\�z^~�%�r�
'�t���T��[��jTSčam}��h��9H�t�'���O~���w��si��i�I.��Ib_���������sB'���u�a�Or�Cc0�cϲ鿙%1��cl~�&a�����2O�G[{ u 2a�D�*���O����~ ����@V,��M�G�������d��PV_�=��Č�����
|�v����h�C�'���g�����:��5Z�/r�N����kW���˰43��"ENˤc�H,�`=|�BCo�C6.�E[��1��e�Y����m2MV�:A����x̉,#f�#�_�	�9�^3�'�&8�Ri�Գi���N]�m0��kI����X�?_��c��)B��b�uI���;��DC6R-I����?�dx�R��S����]�7�\�:e���W.CsvڝN^`���2�Z�z0���)L�T��7���)�]�E�z���p��	��"|��t���D-
�����CC7�6�Pǯ��P[\DW��L[��R����]���g �}��ଈk{܇ݿ�+�!z�����<7˅Is����}D��fkP��س���ր��p��q��s(�T[���{Jdv{cx�p��s�S�>��h�--A��<"k�b5�NUB�����
4��$ϕyU(�R�7@�z1����9nqy�l����/F�����vR��9���O�W����=c�S)Ű�0鍫�����HYzZ B���a~��'���5l����_���3
J��iu���	��g�v�U��\���z����L��I��>���w*���q�X�cW-r������X���cp���D�W^�	��`����� X�1��e Ǔ5��S�/�b.�	Zߌm�,̘�s����Yl]a��"��}3��
�����mk>�>�!��r�3;y�qf,�W(�b\�KRF�M���(�l�|}$�3�x+p���ކ wE��l�"-��X�a�����{�HG���z�E��,�(|�]1?7�Zz�cR����ԥ�r\��^�ܟ�^tz��#�#ШwN�ӏރ4�m��Ѐ�F�:�Q��ϣ߅ް�Z	/aV�=�2<�6���G�~vD�5��Cm��C.N��y���Q
����������t���J�����6�\E�~�Q�eG�����۶���\�cD����t��ӧ���#D���7�b/���9�c��$w�����{$=�!x8�i��u��������M�v��}�G3���_]}��ܝf��I)J��}�k���q̰�h���5��݅��#8�887�-J'�b��?������ῆ�A�ż�,@���ǳx1�HCdޒ�svʈgc���X�>��j��%�OK��"Hщ��㉸�]�XE��T��<.*1AP�`PҸ��p�yan���Hj��d�ύ�/��1��k�I�&�G��щ@Q�F�K/�1N�I�/R��ua�$����S3�|�폼!��a�j�P�s���}��պ�f�7p�c�����ɇQ�+)�1�����gcld���c�>�k�ks��Z7}�5����3)�kH�yFI��&B@F���t���WC+1'��n���
���l�;�.�m3�z"��Ȱ��)|z�1��N��h�* �{���-��7ނ���G�����7ބ�ӂ�V�:�^i�k2�h�O�ݽ}���/!�n��hě�1��o��X��	n(���ʫ�_�̯\���G�H1{}��>��?�+�&._�_y�*�>~{{�D��:ڇ���'L���xfxYZ
d�I5���.����ސ�ı�.H*|G�8��!m
��>�t,���[�D��M4������<�������>#D���ɪ�1Z�T�L�m�.q�x0�Y�ᤨ2W�Ԙ��z��>��^{�:N`x���
&ؠhB˟RN\MF}ҰG���A�	'i�c�{���@��TG%{f#��e߃�b-smHB�{�!T�s�F$D�b�Tι��$�yG��,��<|�\YX��!2��|q}�@�=� 0L ���[6�8ss�(W3��35�̍	�����NJ1�Q�L:�,��y�1gMkH�6��K�����n�P��Jh������!E�P�cV�F��9	h���4[�|C�O����ĺ99�HX���-�:^�L�	k+�L3��e�)�Ą�!���v�;��L�J�@l��x����;�<;_��
Q��;��� �nʙ4t/@��f���:�{m8C�[_Z��C�^ ��*�]� �^���1ZV��Xk�`���&�]��P�1ҝ�Wиp���<����T���6nT���Χ���v���8��@1�v�%�����D�H
����'o����C��W^a� a�兔Nǋ+Щ�8���*C·�u@��� q��lN��JL�7���3�_���x�՞F��r��Ǐ�m�{�]�b0#֬[[^�>��B6�[����	PW�&_�?�7?��?�6���e�F���m�,���E�O�!ˋ��,��&�mΩ�� ���i<^ޓc������)[�iue����,Tb%�����Q�N'42\�V�(=�+c>��̍L�"C��8u0�"	夒�{n8.�u &i�k����&�i��W�C��7D�vn�ȝ���I�Jb��&
�0�"�qfО��I��g������{]O
xE��W8>>9��nJ.g��S��C�&S#���O�*�c�rB�$WUFv5bUjPA`P���$7����ڝ>���q	8%�F���3�&<���J����2����7`�un�A4<��څu�]]W��'�]���>��X.�-�.>��]��f�9�}�7���ޅtm������l�|�hԹƄ�_�}(!:������,�����7��G���U���{p���q#I�}(�8...p��G!ݳ3	��r_�y���D���S���|�|�&������qL���*���0�EQe��(�sC������͂����<�{�NG����-���L04�%W�����$�����"�X�s�*7��7g`~���'p�71=NN���>{���и�w���Tq��NO4έS7K]G�e��\�8�jDF��7�����!I��kӈ��PY�G���n: ������G�Ll�j,�© ��M������q�-�v$M�7;��P(!�0¾Y��*ĕMr������4�CsH=F.�|�̓Իʓ@��&ӏ�kP�S��0YP�G���PbE҉r��Щ1�p��24���/ǟ>���C.b��k1��~�p�V������,�H�Α�|"���S{g\�YC]G�LƱJ����r	;i��?����yv����߻7^~~�W~�f���������z�\l\Ec��kp���pJm qM���qP����Z�;�`WW��W�wփ�r��^��m�1C�'����R�&�=n�FP�]�ʥ+p4�փ;����Y� ��U���P���aȠ�� v���	P~�SyS��)�"a�(��Й�_�Ȍ�%�K��fI�$v�m�,n������S�v�L�0����EV�9������h���4z�+?g�<��Ĥ�F����"��0��ߐĜ��a������ݪp���?����_�W�n@mv�xS�Tқ*6�,�-I'*�� ��`gb'h>�G�B%}6g��;���Ɣƀ&�5�p�O"���d���Rdr�ȁ�2���(�L��|�{~��b����XrT6&;?I,fvjj�,�c�\B'�α�2!)qΑ�KJG�e�y	��0�@Xz�Y(�#��zWrO"%Y5��X�2��׉�	L�I�q�!T�xx& :�5t�uSP�L&	j�̂ܓ�xv��@{o=?�V�$
�q��S��Ȥ�����p��U;>��@n��]�T -�L��i<�gA��� ���"
��J1�w��]89=�+/]�7^y	����ӟ�-x��_�ڛ w�v��0���d*q8�{W���rs=���h<�hD��%�6"�6@���<89�K�`ϵ���w�P#��F0�e\�R�V��1����������;��Ce�)w[���{�țB2��[,oREo���ǉA=6�^J�	N*yo�b�V��I��f��D�5	�w�d5�c�_f'��#l�R�]�=��B���y�w��G.:�� ���	�_��
�FN�'�:+�����G��G��ԡ�_����`����?�3��;n1���F,T �����y���<_9����)�_z=Β�y9�b`��l㛿/�4g���?�@*�i����gϟ�5�����e�4�Ђ�L�d.����>A�U�'�gn���ٟ�v*	����E�üC�>V~ε�q��`�󦤏������{������9R��$2����{��}"e�FN��H]d�G�B�X���{[���:� �L���Za�����ZZ^F�^���M���TǏ�X56ܜ;�����bEz�����XY����<�ہ��_���������O>x:��z�	��o�~7���b}��#��Ϣ6��6��N9U➌8o���)n�S�m��{P���'��2��.y�h��o��/�c~��p��NqtK�W��%��x�����S\O�;�\�=�K��O\+�l O�nr���z
}-/�`emM�o��)�c��¸X=ek��-C�I���32Chc��ln�\=O�w</�_̴���e���|c3x��x�e�ɫ�:^i��a�0�ٹ:�enW����d���O��S)|�W�o���}�M�9Lb�I^��W��	m�fi� �;Ƨ����"���H̗�(�����y1!�W߸��'p��}8>=ᐁ��̋���s�u
K�MC�*g�9B�$��o��-Ƹ�K�ß'6�Pk hR?3��؇^�C��FSH5{�1�L���-y�hl>��JO��x��F*b��-�a�Ԑ�p����e��c�ʄ�Z'5�"�H)�|��rG`1u�D�2YS̼��0J��I�0�(�ƹ>3�F���?�}��fc�[e��fi�X�d�9�E,K}�:����bc8i��pV�^�U�������_�>y� ��7n��%8;9�.I��KP-&PF$N!��� �ҳ��Zd�ƛ�+e�i�B��z�u) �&@�9E��'�������~6�����`�#J�Ҍ��B).\`��
z%w�ށv��{��/�o��ܹ��P;ukZ\Z�1¿��v��ts�B�;��Z7�����gC2�3�����Ў=���w�Ph�h[�9*��	R\AC_�N�h�w��R_�ýM���������C��/����'�0�8��ܠǍ1�Mc���=��9��t����i�E���&`,	u�̔������)���p��=0ʊ�y��Q]k�8��2�� ��	��|#�L��}�G�O����=������M*V��D5������-�7~�d*ɮ��7���q0�z��fFk��y�q��{2������mltG�H6�lwԦ��&�|�!�%f�Mj7�s2޺1+�b-X������R�7404��懨B���b�$v�3�焆�2��W�5����mh�����Jb��#�M�ApJ��}�s��a�v��a�~�{߅�������g�r�*�
e(�����1�y���܄&���֓M�Rw{=��Ն�i�n�s)�O�m@�/����GP��@u�ґR�
��]�ͼ %4��b��:�?pLNOZy�9�~��*3�-�D̓FBrec9T�Ka�� IƝ�D�Iq�\�0�u��_�C��b�Y����u:�N�t�t�	���-�tr4(��� �o1;6Db4���o ����C-�j8�gȣ��Õ߆��#�����q���o�K8ƉH�5�&�����/�g�=8�)[�,b�^���+��_"�I�q�6eDA��+W��O��K��]��<�q���0<���:/�zn�Z'��'�"�_kq��Ǉ-,Co>V>?�䂋x��fg�Rb��(�9j��{f�$�r]C�΍�pk��i?nD͖(��������|�DQ��]����͵�+)��8�8����$���;^���C0FK��?㢜�nWIt=�\�8�1��"2�.�r�����l���z���Y���~����6'Pi8�b�ßy�.}6��H�ʍKpz��Z� R?89��;O���~��K߂���e�OYkogκ#8B�|?�7�<y��:�����i�,dM�#D�@Ҿ,�5RO0�"�mf��,�RÐ��A��$cH��h�TJ�8�F�&}'8�h��=�@�N̞�/���R��f��A�$�F�E�pr�ml9~]&����p3��I�n^�p�1a��}������oȂ1�v��Mb�(��I~���u�����n��p�g	or������.ZY��������]Zƛ.��ސ��R>�Pf����{�c�)�Y��N��Z�����{&P`��91'p�=4$�$��v:�ч�Z�S1o�6�9�����&�RO+�qL-a�!'���&�9ې�����鹡�<� �`��D�M&�O�ys�Y�S�gY�.��1��0�����XP6�ZH�E@��%FC����"�7Dm��� �s'7&٨h������L��Ŭ��HXH5c��ޗ����+��rR�.DÅg�z��2����:G�*���jisx�������C$\��v/t�]�U0�"����y�9�"�r�*��zƥ|>��,!B�zt�����i��:�8f��6����=�Gz�!)�3�J"�[�eQ?c
i&���u�׵)���[�~)�K�fen%\����}��\��NK?����y񞎂��/��I�����b$ɲ+���|��3"r�\j�ګ��z�^f�IqJ���`H � �$@��џ�!�@i$@�p�%�b��&{�t��]]��^�Y�K���/���鞻<3����"y��##��̞�w߹��{�[o�E��---jL���z�Ff�����o<�O�����7*�j�ciR��LS??�����n3�Qʛ��o�8���E��<b	xL�A�y�/���^4)i��?����ܧ��_���!���3�d�if�hgc��Pݧ
�R:�!^�{׈��Xp�yօYD._es+�hJ��X�3 
�݈�F���I���ߤm^H���J9iKլ:�Q���Ac�0d����rѸ�L�7H�Ѝ���ʱRy"*<@WNH���Bn��^[��Q�Pvy��X�gʴ����{������Z��)�`�NE�$w��AM���9;� h��E�T��F^�֑���c+��ªg�"2d���E(�`�3��J�k��E�~d��
���j�O�Tr�f^4b���s��c�{ホ4������Z���u�1��"�CH�c���ct{ppHg/��gj�P��w{s��_~�v6��_P�uM���KW0�dYBh���;;֟7�Q/����t=�5��j�	&J=����.��˚�=y,�e2�k��q?{��h<�y�]m_W��sZ����TH�-���_G�ZY�l�:�f*�(ɨ-�L�*�5U����q���"�#��q}M��(�o u���H��("�9N)��H���X��F�Ȃ���:�I����dۥ�w�ӵ�$)��N��Z�\�?����o����t���W�L��/�"��<O�MF50N�亻_�\�/��_/�ZZE�+�h�����HޗH�1�o�����ի?����?�{(�n�	#ЌR3���T�tT.t1�F����Kq����`�p۩��x�o�� �Y%G���\L��/���'�s�Oi��0E)�BU��9e-:�~�����E&���F��l��p<�qO��[3��HLİ[V�C���*սM�ùQdu�{c�	C����É�4��T	t�-�_�E*�r�

��vo(u˟����V[n�!5=�hnqV����kt���g5���~b��I3V��RY�,����ߢ{w����5��[���%:�	���!&�*M:�����+�һ$�L��un�%��%RئM�<~�`(D�_�~�I2���k�G�_������iE�^�=i��.����ӧ����bإ�??1�ﯭ1�$Jb�Fn^z(�3��
�kG�x���=4m,?���u�`�q�����܍ZA1���w��sp�&�>����TG��A��&ݾ{K�;`9��K�<�}��?ء��{�s�m^����_�<��6��l��T�J�ӑo�
O&L(T4m�x�
�n8p�C]��HK�փm��7�A��{�Kw6�h��}f���]��6U SU+�x��E��&�jO����Z���{�3[���aӤ�zO�Z��`Ҩ���A���\~�W�f�`���k0=��^�\f�;b�A��Vi0z�e��-�����xnt��O<����e.��-��3��'e:��۾J�/�h��q���%�E�^$�Փ�壋��������m :��5�0�A+���0������d�=�������n�Z���z�6�ަ�h�������G�A@*��C�C��{;{t���:�,����<
�Q���$�]h�4�����'�EIq�D�r��6�Pf!ya`Ȍv���vé�'�'�T0�^<洕w
s;,~���(=L1��\�"<|�[�نt-Ndl�޽G���inv�b&V%U�����E���4�|�>��b?Π;'�?Se��
�ߨDV!ܝ�$�,_�4ӴK���k���~��2�◁H)w灂4&��J�B-8)��"y�)�]x�=�	�w�W����o���EkK������>��3t������f<��*Cvc
��,�����(����5Q�+�#�WȜ�by��;�{_��r�*�򱑭�׃ȧ&5�
kP,-?�S��~�
��U ��H���/�hZ ��\h�̹[GN�*�_�(��K�TfX�}s+
� h�����	My����b��X���t�fWNRsn�QxS
lD��)iS6�FsF��T5zvP��V��$�2L�kqhR�L!ӄ�j�u'�.���]>Wo@��j���E�:W�/~W%~@��S*}�؀�*FMV�Q>��`����`�A�-:��D�JL�I�ŕT�z'5F�cDE��D�4׿���4V/78Ui��`b���ZYD��oT0���>c��B��˪h4�'6.��U�/��<I�Ǖ�-^Kh6��h,>wըV=P)`F��������W�E ���9_��nܼ!�������o��o2�k&RBT-�@I-�Tw��1h���GR1�45�A�G���q��<�*���Ŀ;�S��7�r�F�c������oU�vI���>�����$�	�)�`c!]�cMU� �A�0B��DXX�������GNх3'��|s�z�1:8�Y(����wT�#�HA�y�/̳{�����)��f���w��O��O����ޭ{t�Ǜ�	+�Q]�ߟ���M��Ga� �јc�˄7�yhhL��e�d47�x8�!?���� @3V��^U<to�D}ve�� ��{�,�zv��
؍|��E���,��5x�.>��%j�/�n7�DPf*��@�1�Ty�5�Z���8�N5sB ��e�9�R�E;u��J���[�ǧ�2l�{��@�xk<OWU`��u�8m#�J�P�[�{0�=��(����7c�`��@�t��)?C"ّ�z?6��r�ΰ'۰�z4J�3u^њ�������ˮ�Qx4�כ9(#�p�s�o�7��>�mu��	cY룑o�4Cؗ��Й��l�$P:��J��w#�$���SO�f��믳� �K����#p�8ϭ�-1�8��LcL�I$�.MJϵP;��Ә`�!F�����O+4�G�Ww>��V~{m�g�����)t>�"�����u6�
C�����r�D�Ǣ#��:�ԝCH��>��T_P3����%��FZ�������K�s3����?�'�)5���H
I�X�#������{VWy4�8�F������>�����o��
�u�}���5F
T�[�G�O��jȜ���-�p&?�m�x&冬�����1�i5h8�Ӡו���S��<�G�k��̤��\�!c���*�)D�(�ł�%���Nn�<�!����N����ϕ� �%�t�g��h�Q��z��I��cTg� �=.��,4�$�q��͛�t��|�殧f�5�.D��FS���Z����6P�h"M*(i���j�6'�f�(L�Yך�<��6���H��d�gFM��C[�A�ds�;�R��PS�,}�����u�^NKd�с؁H{<�P!�0��H�]�xNR�{�[=�P��)"�O���i��b�`N�X�s4�G9��VvJ�:�.��Ӷ�C=�UN�؀�AGAK��zrM�2��{x�R�6�":<���;wD ����Ok9�BG�
$�͞�гtZ�ɖ�d�|r��P�̃c,�Q��i��s�nV}�r�<�������/�m0VdUoi ��Jv@\@�kkҎ(��;�˰�*�ė�(�cl��7����to�>ͯ��c�hc���ߤ�����~���!/��)��y�/~/���	�d�7Z�'���M?~��t�����_|�U��g�=��L�|�G.>FK'V�򕫒�%<<�J�4�K�t��Oy��T�n�iMMX�Q�L��!��.������,j{T� �5�qzZ�
���:�+�]r�!x޹�}t��cd4ZyFCa�n��S����i d6 �C�٦�������!QԤ�D�5)T�]��R)�	R8N�"�|�>ݠ��������$Y��t�a�%�t�-qy���i�F7;����Co�=\;6����b�"�S�񉛥�^�1C��YcB�d�����9�q��T>@�l0lȵ�@uL�*5 ���aSj�w	o|6�1ޙ�>���$o��s#��k%E��h3yV0�8�B� ���p���+` �B�W�D�N��K���O�#���hB�z�l�z� ����5{bu�>��/��+�i��o�Ԟi�y]���C�V$ �;�Hy�7^S�0�Fj��nL���	���y�I���z�E�ql��9�$��>h�g��M�7J&g@�0�|���Ύ�Z�z�4�����["��3 �6?��\�~�3����7io����"md^E�I(׀�� Ƣ�*�jǔ��E����!��G���(jp����ݸI���6w�����H?�����R}�#��!#�]4�f�.���`��v��AUa)������O �75Ú�x��d��i���H����ƗO�zG�ĐfkH��� �DA��,,�4uBTs���L��wx�ԣO14���;e��\Y���	�%H��[�>t�z@�r��Z+D��d��|6���6Cj􅴚+$b!�rn��a4%P�5�ޒH78	�T	'M ��Gf|�"c5BG����ȼq�d�����
�2hT�T��k�rxeI,V&^�D
�P�$O�ju��14
��W3���K�4�.
��l��JI0Q��#B)ˀsHj�I��-\����)��:�/_S���DO]7Q�G��6Ep���x'�84  ��IDATbc>�ml��>�{��feSɍ[O�/	~�obS���ey�:�z�����oE�Ib&�
 @�c?��F�F�)0tu�J=�O{�?�D�~�c��ʙ��ˏ�>�p+���;5W(v�!*.���p���䭲�$�犀��v;��]��ݥlȓ�ތ-�l5�e8Q�s�3�!�9{�>���h�w�7�쨹�8:��h4ϥIp��7�eb\y�:���~�:3��:��WĨl�v�?.��ِ6f�?��v�fظ�6�km�隘A��@�cn�s���P��#A3&$���1��GY�p�� �h'��m��x|x17sŚ�1/��G�85����Uts��!��AFIC#�O4�o��;2��)�Jсvi�}�N5��NH���-A��$/"�/$H�c����oʦ��Vu��6���Q��h�<j�
�
�frE�²h$��4���!V��צ繁�7�&zo
z��1���MbERJI����!r}��e���c�釃C�����Մ��^�D�5�(�A)��@��&�}>�2r�˜�&�j])�g��cut2�ڬ�J֓y*8��!y] 1)rd��&xm��ӑ�.�i����^�'y��:�ݡÝmIV@rҐ�9:2��H<�\�@ �,�Y���S�����ݣ~�r�i�Lo��x|�c�=FW�^��C� �5~�#f����a4�O5������M�X�{勰�M��&���¹��x�L2;��表�Q4���Z�`d�.X�ݮ&���J)U� �4A�O�&�o��-	 ��CAk��C�+'���Sp�iMQ��7C���oUڈ�6��g�xp��M�wq6�ˋ"w��G��z��(D�yC`#�>`��F2cL��*v3��WǱ��=�gb��y�zMEw^/@'�Z��6��Cd�g�>�>�p��4){̵U�C��5�/��a/,�����ꎖ�	z�>�,�|zڐ�Bh�TE[xl�����4,�|�]բW!s��ܐs�[�����!��*9�fM�p�_�X #�K-��7�{��B9h�[u��1�X�i^f����1g�[��VE���4�@����҈'���fYa�֝᪔�'�����>?8���b��a�r�
��Ħ��/�\O�])��3kdB���\@ �� EV�� ��[�S�,ڝY<m�:b��OȦ���j�)�ix�2]�6��/>vQ��AW;���ƽnнkWE����ޠ���H�")9���e�NF�oN�<I�;�t�xV�J�,��y`�9�^|�~�g~�~�W~E� a��f/vTJ�i���#��EJ��y��}�a�8J�G��u�+�s��*�Zx~f)��Նn�,����+�<��\�V�{ݓǀoll�D�g:������S���n�DY��v�Z|��g1�TB����y�m�b\�w�&Cjluؕ��șӴ���Y.�:DÂ,(͔��1� 0]���\�~�n~p�Q�<=�Գ�L�����s=��3f�5і�qAI����f�3I*�=�c�p/���(��Hn�u�/��A�Gl�P�ͦ5'F=�x�D�}B��	�P�Z�k��v�_�(�:�y`���)�Eg!5��Xƹ5մe[Z��cA�Xh2�F9ט��<IFP�,`1v���A_E�\�ݖ��W<�`tS̭0�E��5�
���>�l$�l� �����q�E;��^�n���z\�;<�24Z���;-45QR�
ϋ�ʕ�^��-[���	>xꐶ� �T�X���gq�
MQ�"x����Dh8m�d�R��9,,Rga�N�}��<r^�(��G�H�gg�بvy=��㢹58�&���NЂ���͠I��e:��u�.R������ϿH����wߦ7�����^�.d���"n���Jڻ��w����y�t�	:�ߣ��mi��ڦX��H3`^w~�_�o~󛴹�)z5������Te��*�m���j��5��0��s�����|Q�u��Ү�e����`����z�E�r���~�:�ɏ��N�˻{�m����pD�lࡲT�`�S����`׋H|�P&.P��.-��g�Iw��i����϶[���|X�%K^� �,3C.�7h�M �[#⭭�v�4�u���ߓ�ɬ� ���� A��ޚe�1'�h2��L&�����B��<(=�a�]��̴�M��=�h����ȵ-c'vݛƩ°�!,F2�F�H�W�:�ZDj�yd,ܨ�bJ��,���gݤ"Z>2����{ŝG�}�Y�-x{u���޻K�K������<��D�K/�l�G�0��s
q<���X�]͂מz��2d/�p)�i@��i������,�Mx��&�����ua3xEi�n)�Iyo�B��̪��F!-0�����ߓ@N�G�{43�҅Y�7��#I�%^C����]�3l�
c�A#����0{�9ty�~n�:+'���Lae��s�A�s^��CJ���у�w�k��=i�g��٧��62����yڛ�g��8��j�:��EZ��n���3�������۷��ҩ5:;ۑ�F�ȳ��" %
1U� �4)����_}O�	�Qq����,�_�/Q��˿Ly"��6���Yro�Ä�$!�J����XY1�Y<(�a��sWZ����o��8�B����mu����th�˖Y�	��YM�6�ѐ6����5����RH�⛾�c��c�=RS�%ʻS�,���gCv��߀s������9C'WNP=Q%�$���%8��� 񅄇r���6�h~�Csk�������,"*��S�����#TK��:bՕ��Hب�r��TOK�HRͩ�'��H%&A�A�X ˾�+�[,���SZ�26�I�F+8
�^��1�=|�6��R˒h�'S�el)5QD�)��y�(�Bs͕Z��X��T+\�e�ϒ��@���?��;ذ����FmHN���=Y���x#n��ػQ�tH*�ȐXaߓ1Q�pKz ��q(��w{��K>'y�t�Y	�{�U��]�eM����,��dꍦ�tv��Y���+6  dF����ĸ#�H�"5eK���"
��$�Hd����i6쳴r�"���Fm32���M:��������ub�,�����Pp�Ǟ��C�:d� 8�Q��7l�}�����O��P����@�<N�ФY�[�)��۩>]��S`���=���M�v�!H_�k~|�5CK�K���9��/|��x�����5��j�����<�*�*��cOZ�S����F���C��6�w��(&FY�}>a�Ǔ��w�m���ʵ�Y� "��NM�\�ro5���J�'�>�0���x �=�ۣ��u�C�?�
�Awv��ԧ!y2�{c:(r���J�x�:w��.��,��������B���+��=^x0懻Mڣ!��Q�����D�,�;9�p���Kl��:VH3�h�높j�Q����µĉb�9�SH:�ʉd��n�;;v��n��Y�)u�|��+�@`���H�����2!U�NYF�!Ѫ��s�6�8����=�4�r��|_ni�����r���^�|?1�\�h��x�LHUA7v�2���,�2�G2oPы`%ϵ�.��G�|�%3K����Y`6Fl̡M5{#�4`/tJC�ѐ�����rO0-���#����`�fj��I鸻P����wh��'(�^�%{m�c����+�]�=ͣ��0��)d��Cg F�	6�V���'(o�����6�)�y]��0��Nhg}���:1dgԦ���������h�=i�ԝ��:G��m�>_T'�>��ݡ}��jH�(�������"U��԰vA��>� |~�9���wޡ'�|R~F�TY�J�a��q�f�tl1-��c�ԇ�b��\����EU:`�wpc�p�=9آ���~�_��D����=1�����SD0� �Թ��/,)�*���Xy���y�wud�������R�?��׋˴�� �p���]�y�ipx�OhiL���&=r�3t�����5�]K7����'�밊δ.�쐏��z�߿s�-��Ģ��T�j
M��ƙ�EɌ��L�C�t��M�df�h�*��� G��!~�_H�ɕc#�ޗ��n���^��.'k�+Pf4����	d��E4�q��9ɢ[�ƾ�YM�~�ڲ8����ZCj���2����c�"�.��P�n���̟*�V}-�+�,h�?F�Ar����!{�}��Ӯ�v#���e`��Pz?~?|��(�����(C���-� U�z�dFJ�{qϡ��E�g>����D�;�(�� h9�a3y���I�TGlԇ�<��$}�$~�k1	�K��4[ԙ_�t��:�����O�d�>O]��HUmHƋ�BH��B���^DhH��?-���5N�+R�Pkw�My(�b�ϨSu$0�#�x�����O	8ٽ{�o�i��,2�f[���zo�q ��P6U�!;�6��N�9Cw����ŋ��|��y�N�N�+9��ח����Ft
��q�t5���}���J,�za����ަ�+w���s�(����K'Vi܁�aԅ'���Ƨ�+�IT_`��ܹs4��4`s-U���.�3z�������Fy��髧V��ڒ��y��y�^��<��1$	���?<r�7F���k�^֤pG3*�|�Ip�q�k*�m@�#ޔh�7��v/J�5u��׃��m�]�P������Lr[ع�\���S<�F��m����]j�)��KM�v�g�c_+�20�}m�&F3�<�@§k�����B�xT�:U|�"+�}��G����j )��/�(�}�覠"��>�+���Y��8h֎�/�8�+�{�Ըk�z٬#5:L��-�F[������o���g�4a#�Ќ�4�����c7���	�:�_�Ә���c|�i�ը3��׉e�H�'z�LȚ�wh���JA��힋l {��.S6�5 ��FB6�F頚$��C��F'ٸ��s� '����iZ����ԫw��`G ��*�Z��TG��3kD��6��?s�f��kk4�i�w�1`CQ�Y׈��jLkX�8C/9��,:����M��A��Z��0�<`�d�W)+��ˤsҽ�����ur�ԭ }��_8O�o\��_x��@7n\{w��i��Ie��TF�QM����e3������ڌywwG. h��|Qk�A����3.F;�h0� 2�hV��Z�А�!F���W��� ,��T�&�h4}�'tM��v�;�R��Jd�$O��0tb�Mi�獠K;�4��}-F g��q��YZ[��L��R&!��K�C͸�
r�!FO�7�|��\����C�V��,6��,�h�"�����wRħ���m.��`�>�B��H��]Я�Բ��%u#`n��jXn��h[!�k^hŠ�{�c������EeB���=C"(���5(�/��#�)�f�m,H`ܗNA��.���&X
�f�$�A������������?������$���R��sR\˲������.�i��	g�9X��!3M��!D��*D�G����$P���h� �g0��L�I=ՠn�y�w��giqI�� �L�4��*K%���xԓ���A]j ��-��-��bZ3�7���1�yJf��H9�,�(m�V��T��t��S/��Z���¹3���}�,����t�ҳ�x�Q��%������)� -�nc��gr�D4��]m�v����U�{4���h�R*����l�+
�N�[c��6���<�9��:����[��k_�����=��s�ĥ'D�o�}QvKT�)�̙6���lJ���P��?�?�!�Fo��{{{����H7���M�b�.�Bq s�?�%$f�{G�E/R� �1�c���&��I-�g��*�𔾝pKy�E�j6bρoZ�ox���.���bKh���wi����������j��@��tى�F
���"�>�6ֻ{����7xC��7/Ԭr�ϻ�2�5>v#����H��EG��r�JKZ�c����"��u��М��t�#�7v���L!�VLl��u�~6�d�����T=�����T���IN0h����J_H7�
xV�-=J��<]O��E4UO��M�M'yt�c��G^�U��.�
/��M(��\�2/ >@�-�~�����:Rk벡zS�B�$y�
�2U53iZ�e��Ze*�7$��RM�{r��O2 kmb��(�vf��f�.Aw�Z�VF���$�p��X�6�ip5���6��zVg�T�\����5��Q��-���=�����������P�P{P� z"�$;��"�U�|�c�!�Ԣ-/��~�{gi��6�~�!�?cixUȺ��B ��\Ս٪�ӆ��ES���
ov�42��y_���A�3����l`(�jG��}F��yskSdﲱ����|o}�Μ>#t6^��=~�G�8bH?��W�B(ӅH^u���7$*A� Hp���~�>�H`T\@ٕ�g�)�u!�^��j�ʈGEn<�>��@?�/z���uA��A,�f-�M�ga���t��C�i��	ZYY�l����NG>�*�����'�g��n*�)q7R�ׂ��s%R����[{t��]�s���D�m� �&'���p��yq�=��*��=�`'�X�+4�W��2���c4�#�h�s.ՌF�b���D�2"oΫ�qǆ\r�k�ZS��I)�{d�a��B{�T^�SUM�H���&��e:#�`����[=�@^;���<3Y��Q�B4#���I��ԤQu�ո+�_��ق��u�g:lX
ˎ�m�I����r�B)n'�X.�3�C$�$n-|,�hv^wP'd�#�6�h���;Ǐ���ݕ�P�#g�R���{��U�\e��;��հ�8�-'kyi��f�Q1 �t����|�kS���3ϽH�=�)�d�����P���dt��X��SYXS�c�^|�:dw�@�g�MU���kYZ��f
�;ѦX�-a�{�;�]�%�������o�#ϼ٢�%6�}�^
$L9s��˓O]�Cr ��{���Ͽ@?����c�я�ci���㏋$AjAPշ/��G=�v���U�t4�'瑿} �# z��M��?�sI�Wa�����]�[t1�;�^�D�}1`AM��x"�5A>����F�f��ه�����赟�X��n�t"__�K�؄zC����~�3����կF"�"�[�L+���U: �1ycl�
�����Bc3D ԙ[�5�����8P\�
J|.�j��葐�B�{4��{�ʘ~���q?�f*y_��1�*���K�yHs�NT��:�-� 5���S�x´Q��Ӓ
qC��c�|&%ǭ��\�'����*�wd�#��!F���3M���� ���ю\�t�9������P�����\фo6q\І*�%�(�D��d�SV�v+*��/(�D�����s�!�cB��IB@��YO]�{*/�P݈���D�nݽC�;�4�tB�s��/�Q�0������"�����g8cΌ�]�]�����6`��5j7io�=�&ږf<�p�i����h�v���ޡ���Q��OCa����t�
k�k�yU�%�FX�mۛ	���6��\�ƴ}�$Ͳ�]���I��T{�����oߡ#iQ.%��kF�Õ5Jϝ��fM��}�58�"���q�ZBF���:��]�'s�����G����c t<��J����ҵ�ߗ�v ���ud�5����cV̇uC:�ph�4���Ţ%ԕ+W$8
J��)��,,� �M,�;�\ΉO^�u!wIj�����E1��W=	��͜H�kmQ�Bx;�;ltk����F�8z�dޞi��q�6���[�~M����Y0�KהA��mf	*Z�B��C��W�����S{vA�B��TEŀ&A�ň�D����E�#�1A�0�հ�a���G����G)a"ԋg!�����hKQ�h)y�/D�B<����� ��h�d�.{I�DN�TGl�W�$O��2̿����TnD�iu8R�˧�������U�h�7D�/�߄g�ܸ��,�qU^A� �_Xw<���V��:YM����k=
�0waL���Md�B�M{l��l�Q�1۞�6�u�Ǔ�H4���5�������'���o�A[�]�M#��ܠ�++4;�J�%t��F-)zF!Rwo����XuZ�Ohui�f��v6�2�ۡ���T�6y��s/��ݠ�y��z�Ҧ�"#	����_��x�*&�(Lְ��-�����������0�:��X�ݍh~�4��tI��9{[�Իs��6��>���BC%���IL-����=①:o�I_��k��+W_�i�U��{�b�-��_���6{ǣ�����"1$6^)g8����9��Z���M�t�b�B���C���ZUh�Ʉwe�6$��0���1NT��3a��$_�����~.�}r�0x�����֦<��hb��D���'�C��.�����aj��A��߿.%���?�/$�j"#���N g~?t�뭆��a�/y�Mvk�y��#��2W[#��!�-�@�d�O�I�9�XV^T2c,�Ń�~�+��Q0��a,2m=�� ����XA�K�P<�����������`�I9/�$F�s�eópIY�/�J,��ĳ<�Z8Rt*Ū#�u�K�F�.ߐB��q�u��aܢ��D^\��#f����`�j9�
��r����%Ye-������mG��Ý*@7�mC��WǨ?��6wP1�������9�kfO��A�Je�q�6���x@O^z�^~���������'B�����.��4���g4fH��R�5��~�g�p����>{��������;�gߺ*�z<n�Lg�N]|��v��ݸˠi��KGx�rT��5��K�
)z�4���~p���<n�)޻�F��b�7��Ό�w�ǧs�Uz��_��]���M6�}Z�n���D�l ����0��k٠^ʞT���x�5a�3�K�<����R�'O����z�^���/}Vb���!�/�Z����'���ղIZƌ�q_�GP��*Pz8��x�&��9a��v�z�]��'hqiYx�����Ej	��$�l�����1m�w�k>�-]03a�Qz�1��פ�F������ޡݽ=YHiM�JqgM?T�ߡ&�53����v2�sw�����3�<+���,uj-��>ל�OP��4ҎKEH$(�ͧ�Í��7ޕu	$.��к��$�TFT!��+J>#Τ���#m��G�.�����u���v1|��0���]�#W��s�#��L�S՟���(�x�Wy�F\h�d�sC�V,��W\���I�Z&בW�A��լ2����]��ʃSRz,�q�MF��6�$��-�V^��ǍD��\��5��6���7�Bs����q#���lH6d���:�E+%�kT���t��!d)�Q{��6������5嘋hP����ƭ�}�ZI�u��NȔ��M����ݛ��ӏ��_�2=��������?#�7��}6�(>��c���-���`Otg@�����oaa�����a�aocz4!c�����Z��e�i��n����D�P��`K+eG����ӕ��$����Й���ߥ�o�I��-Z`�dn�M+'�h���!Yi��ߖ�Q]��}s�`z�,Ep4�D@�Z�{~~^��"h� �z��)��+����x��c}#s.֒y���L�x(����ǡ�i5��R]��/8!/�mmm�_Ο?OgyDtZ ����9�a4R���X^�.��&�/��H��j�SdS��R)il�[}`�@_BD��Y ���B�)_f���A�F�z���͇z� ��ӫ��3������/�L�st���t��9:�v��|�'�V����OC��`��v7��lQo�H������;��Rk~Q�H�<�[E���2�"�j
:���vx�V&��<C��A�D!Ri����%�nY'X��U=*�z�Dܨp���"9�)ӥ�^���M{�S)��E�Q��H@5�j�:GG_���(�XI[�^_��v���C��qA��5��&	�~(���$zBrG)6n���JHˎ��4.-%�;�
�`��)��"�`�QC�����lm�T�����>Tl���p�`��@�8 M},
i��0B��~zF# ~m�g^����{W����ln����5�[^��/<��E��&�5�	�[�矾D�l�[�Z�J������AO���_�&ǚ���y���r^鈍���ߣ��UZj_�vRg�qH[wi�=G�>�l�:��Z����5�=CЈ �!����U����<��/�+���%:���oF�]�t�����/��L��~��^�N����Fyj�����ʼ�Mع�pDghbE^x���1������+�/�ٳg�޹{[�i��ÌiTO�y�$���~$b��R1%����-���F�����r�I+0���P��;�[r����WxC�{^����n�KjF�J���I%*?�1 �{��U1:���,��C�x����pޖk_��VX�(��?�cj�!Zk��3g��Sg/��_�ƥǩ�Сl���tru�?�P+(���������R���n��KJ䶡�$;O2v�Si��Tx��R�r+�����A�,��R0c���S�FJƸ�\S7���N����	��A���1b�%C��^!IZHR	�'�D)�f��K˝�����k߀*TP�������T^k�@����S<��:� ��u�Fj��Ք`�ֲ�4*��a.��D����xhd���ڙxJd�ꁶE�C7R#�&e��(��`W�%Z�-AEF�ـ���X:u	�i��d���&W�1�H��{?xU������$&��^D�{`;��m�X�M�d`���w�w��o�W��U�����������w��ͩKO��ݸǆ�ߥ�9ʚZ�����Ƽ,'4��]4h���Ν�T��(i�����P�ZhKF��!2��c� n����g��M��s�P����;���>C/��<��̓�� mc{���tL�D1㪚�Zę��]�e�)����{z��7�r��`����J� �!� ��9{�V�O�M��d��6�CiЫ�:Ѱ?L�LOڣ��d��O�s�.�9s�,bN1�$;�t���<^��bɀTE�`��3���m�����Y�p�d���u�b��F�V�$�=��U5^�0]�Kh����@ڠZ�B=_E��Uj�x�ٺr�n�Z�����ݧo]y�N�;K'�h���<��y3��;o�o���I�ܾîr���c��Zcd�5��C{1i��,FT+V�R-Hf��F=37�����N���V��L�Zf$ѣ��:3fE^v��ߔ��VDk�ra]2BZ�2�;
�2Д�ƴxc�}q����xN�W3��siz�N#��G!M���P�� �C/�zMS�Bx�[��Z+;)I�[�Ko�hM@�'�j�W=�k������ݽm���{�y"��L!�<d#6N�� LC��!+4bS��	�./l H��6TV��Ba�\���8���~|���k���������#�Z��Ց��������
�����'�W���t���l����0}Z x���|#�V��y���u��Ӥ�O�z�kϡ�/C�d6o c-��L�f�Vh�H����
Y ����K�����~��z~��y�/�:�k4�1�iPn�4$����|z�a�6�ŕy6��EV ��7ޠe6�i-�1���M�q_d�မ>N�b���6�E4
e&A~�Q/?SJ��� _��eA�j`aI;�9��{B�x�K�]�ȅ�6R�
�K���� �a�a��~pXu�����B����"����M�C�a�.�_� D!6%1��D�U��0o>|nPe�Bv�yG~���l҅���9�Е[7%����M�P	'�)�RќH�!0v4e�҈�AS�1
�FTH\B°��5���T2�T5���|�R��ը'6�sWdܼ�3b�mʬMR�c5���K���NM��7�4�O<��O�B���y�/^��K� ������S2��Dn�
���*��ֈIx���Z���,S)/�ɻ'ɽ����һ��O9�^P^Ed9#r	�'S]�BR8u(dny��Z�}EA���ܓ����\<��T���)��[�?����0��~�#�׿�/�K_�2#�������������t���.w�����[�-z�{�幜���<=�r���$�z�6��cG0���!�4�? ����Z��R���^�Ē����>C/}�󴽷+��v��,^Y>I/��ЙǞ�o��ѷ�����������$_�@�`|D��A��˽�=�|`�@%#����(���?�S�G���N޸q���].�1�%l�K�}x}��ǇO���>�I'�*U@Y%�=���صhwڒ^(�y��I�l(��:%�
�Y�&�	�KH(�r��$��V1^��XeAY�0Ћ�����wsݡAs���FE��l6���'ā�Ƃvc�y!��\���u���	ZW�ԫF�[<d����_��~nq���%����wx�M�`*2�A�(��'����h�fs��k���6wbY.��q>�&��Hrؕ����8e��ޔ�d���b�F��j��0������S�ʹJ��$1͕��:��D��1�Q��eYQ(J�]�g�⊹�9�_�A;�#��V��1]���"nD޺�P5C�J� ��O���;Mf�/4$�B�@C��}y�`�DjtL٥*z=��#�گW�`x>��f�:�������E�\�i�{RC,nr�V�ڽ����.s�V�F�,�#�zx>D�\.q*:1/`�����=��%�zd��`uů�.1�ڧw�ݢ�%�L���e^C���#�/�囷�+������5gZ�#��p��fyl�"����oM�o2|4s�4�����������ѽ�}����M:��B_a��� ����~��������Gi���F�CI2�y|�(X,l�NBe^�)ۡ�yb����� EV�6�گ]���Acݜ`�P�䱼�46�Փ�z�~�O�����~���˂q�  ጿ�%���D�{5��'�T���.�M1�Y���b�#�D�����ct��i�Q?<�JC�{ p�9��$�<Ң��	��}��h�L����/J��E�몛������=s�]�͔�A{�wا>v甑/�~��8� Ց$�2#�j�0>'��ao��8�9����-&`����zw�\�L/=W�^x!�k*�W�lS�D�V����E�����I�u'��X�����+��VPv�Џ ��)�Q��[~�3S#��P�ࠜ�@C ��c���Y:������e��ū�'�
�)g�雹��b�M�V�o�����F������4_ �I��P�e�͆���o��iznn�s�n��&
r��.��ԖK$p��^+`�̗rs,���qW�@3�}$����^��h�l�������싲*��3�=	 cc|��������.#�}�v�6��}Qe��6�x}�:�b(�����&������5�3�S嚏x�4]��ߢӟ�4ݣ&�N��S/�~ڦ�w��̝m:�l�ν�%���9)��x�%�p����|�������6��}Iː��~��l�g�?*��k?yM�;�	�	��㣸3��zǡ��z<ıǭ�ث���z�br�و�#�S1p1#a��P2�jᖠ�+E=�H���3*��~�R����S�<K��֯^�B6�C~���x�a�m���@�S �����,�P��X�d,Xx8_\��޾�� 
9��0C3�Q5�R��w����m�M�>u��x����Ǿ����)�P���l�)/�
�`ԑ7O"Y�(�23���"{R���SO���k�u�����h����>����R�^1���c����%������<ݏ��r�6�x� �YE?s�.�9�W�'�ܻ�ގW�3��D� 5Ȫ�ª�O�M����+���r�}- ��P��JOA�K�o��j$��?d�j:#�<�0�"�?#�VF�����^���-�� ƨ �*�TJ*~��Jt�tz-��cF��u�}��s!�����PN��_���%e��6c55����焖�X�O�@O^z�~��c���_����o�yУ��{�>͜X��;;��:�8u�]=I��;7�w�}ʐ"�ޭ4�_����i�t�S���/|�.<�y�`�W���"6is�*�c��1O/}���[X���z]��Ug8� �F>��C��Q\]%z��L�ɋ�t#憱XY]����VW��l^�Ǥ�Nl�����^�<>T���Rk���_/HK�, x�5D�wx��F
� T% $'�'#P��L��,z�L&-����X1�n�Ę����v��E�blI���z��N�I����D�Oj2�xt������F��YZE���u��U��h����B{�N�s��B}�.�fC�գ��^��� ��X+\���P��3����_a�J���0:b
R�JV��D����+a��ﰍ8��sК�h���}�i�����b5�ᩉU-C�B���]ZRc1��I*^Y峵�M��<�XI���ϯ镠�V���>ߵr�6�0�4��H)7�t��bA�	*T�t��fј�]��@�5�ݤ�lKR_]bV�<(���Тs�Ě3�6�&0n���n�1<��Ph�f�%ȍ:��+���h�b�X0�Z3�(ze�����T�Cʹ�D�>k^�b�zk��E�n0"�o���/�����]��ǯ�M�n����!��>���vƈͱ!g|���P���}�i�}��Fk�fg�f�V�6;O��F�Y[�.��!�a�Yn��UZx�A?s���@y�m�'"_\4fiROhXOMD���O�B{�j��T9bl#(vih�>�@�{'O��Lû�K�ٓ�͔,,�tC�6p�!~Ti5�я��Y1�8�����']��D�'�oM��Y�B�0�{�+��ؑ��j�M-GO���`A+u���	���=qs�[)n��'�
�KG6�����.��L/ 7�s�w������K��w��Y��5��t�w'ui����z
�u��'t���h H*�"����$�T�M1fR�˻��V��`O�Z���0wJ���t�YE��DPq�U��̐�����F (����"�_GX�sh�g���83Т����R������V:Q�k_E�!n65��E=H��I�
�.
��y�Ńk�P�ތ�R�r6j��1|3���kݻ$n�����u�c�i�s;�MK�x�l|Gv���kH����7�ڏ6T�4�:#֤�Ğ�0���s�4���?�]�r����z�*�L]���W�麧��3�J��К��qYc�~x�,sb�K�`#B��ޡ	����u��v�^z�qZ;�Lo��&]��E_�,5���z�/�2 �C�5Z>{�N�-��w4iv~�RF�j�<n�6��G�!��y�t'>����Z9I��Eڑl0Hg�y���a���f�%J�z=��-������% w�4�y�I`w@��:ۯSl�L��0W���u@���(:�K����!��(��q@�8���~[$yQ>�*1ڱ�/��G�t����^��?�ib�AR$!��&�J�i�@��<e7ȉJvMam�
m;�����k�����_�s����~o]60P<՚oɂ�����_��|ҕv�R� ��'��g�����_��d����uZ�֟Rr���/[�҄�B̭.��GIy#A����]XX�OH�:�O��;\X���뮾N3��QQ1�rW+O���(U�;5�&8<d����I���U���g�~H�2��Lv��5xi���8mB��&�&eO�PA��ҔX�t�͇�^UdL�|���i�������%��U��҂��P-�%����tzV(޼G��n\-j�L��z��n.U����r�7v��4�F�(W�w~��$_���[��}H�w�W6��,]�Jy����I1_4e��U�XI�=���_8&<zA��$��-�}�,�=�ҩ�	�{�4=��Ej��K{ِ�����Hlлhm�B'6����gy��0�G����!�z���HuȄ�z?й�bA���L�zv%(L��2��� 
@������F;�(�Ӛ����G�O�-�g@�Q���>:�e(`n`��no�й��*FQ����Y��[b�&���Æ��`��}�+O�R/�Ĩ#`��]��;������B�1v]Hx��� �J�����E`(P��hZ.>�"�)���������l'�"�n�+�\~�"n!xtqG6�<�=Y�hR�����5	�ɫj[j:5��R��e~�C�|�������N��?�6)�A��N���k��k���7Y4@.�m�vE��`���%E���TUè#���yf��p�f�3�ב��Ni6�B+K�sZAXj�*Qt*�HǮZ:���4F!j�SD|dbn���gͲMJ��FՎ�X�!)�1ٹx�Inbp5�+z�!-{��I%W��ĸ����T�!� mLU$�M8����:�#���26��]wi*9�`��^�Py%��d�XMEa��͠"�����8MDB@4>%~$��
�)݉�uܺM[��a𱷿G���o2��J���u�q~$��AFCNR� �X��S�A�6�G+!%@K��`�Q@�Q)�μ謯^|Jd��t{����hq�C����Yf��n��~�ƺޖ��ed���=��цo���`��ڔfVi��JZ|���>6�	[�ep�v됟ж��c���{W���E����,5�����.�%����,c)?"m^�@	��L��V_�x�s�=G�������%%s�졃]�M�`���n�w��g�x�4��l�[޽{����E���'���h-�bO���*s�}b�:�_�>�51��BEN(�����<�tJ,����F�=S�h��o~~A"�k�NI��to�@�m�xgmYDtM���"�F�?���Gؐ���j�m-����,(��oiV���lI�п�5AZZ���F U$#�{H��S��1��1bpi'HyݱU�V��)e!I�Т�hX*�T~�$�A�`h�P�7��rա4�e���.E�,�ڿ'��r��3����<�k+郠E?���81�=�����)��y�s�M���{�>��4mӯ�✕c�5i;:�ˏ0�ƺ:�S���B�%���}�ґ��z�����V�)7˂���DN�4Ok��c< �P͈ls�]'��	bP�ݠ�(  &x�m�Uˢ�cJ�����7E*;M�_rD-6��NZ��9�ӽ[�Ssy�Ϝ��gN	�_�O[�Ro�_�m���;|]0��jHJjhJ����{ܦ+�� U@$���`�_;M������K��$�W�V�>��n]~���f �� ��5�jQ����6̛�>D1^e#"�v;m*^K�1�30� ��Va��J�aؗ �t�{<@����U��n�}S5ĞB�E�;��Lh�`�@���=����������G��'3��{�b��"DTX����4�$cdݗA�(���ja䶊��I�Ϙ�����u��W�#vA������c��P�ڧ��ċ�#:���z��Mz
{+g�=L��M�y�˟���lGPE�9C��:L��T�I���2�
k3��ӎ-�N����F34U�˞�b��)IZ!��-nxD*7�m�?"�B�����M%�QXʞ$m#H�I,H�u8*s��pc���đz�#C�y��޻AvN�tL9�K�Y����c̋jp��©�4整U���6���*b �7^S��&�\n��WWI��[ȝ��@��`�қ�*t}�����P���̚C(�T�f��o��z��^�Đ��{����wWĬ,��
���6��FE����_]�S�0��ȼ�۴w�M�2���ϱQ��<;;����M�jm����	Zx�"%��Q�#�kv����a���dã�a�A~xw�.<v�fWt�*�βG����>�Qz�]��MdN=z�.>��PacT�����
�U&K������tE�-J� <��3��zi�A�/}�K�/�WimmM7�55������eλP�ʔc}�k��	b�T>.ƭn����e��m���4-�x*����Ȫ�~.'���A���7���\��^{M.h<ъP�I���i���i"4Ϙ���Q94(�x�;�~p��,�.Yc���:oZ�!���w�b��	Q��nާ_|���ݯ|����kT[^���>iu�a�)[�n��h+��&���*Q���l���j�<�z�ч��p��k ��.o���:;�u�oI����\GYhX� �a����Iٽ�h���NX��񶂡j�+\y�˘��^�m�iŃpٍ��:��$6h��L{̊Y*��"�A�xmi�|����wW���1���F�ڐ�9$��Zl$�#�s"��i��y&���%M��$W� ڭ�fO:7Y�</cY�pJ5ynzR͚�{�Nd<@'���!1����P��χx�v���\���b�~8���C��'��6@Wi�]J�:1ӡ:bD�����K���HL�Ƃ��=EPyaV���l�^
��`��>���}��C�/��Y��t�Kt��%:���&t|N��Rq>e�������'�xB�F�������/-�,#�Mǣ�%�$�	�5�jL����R��#�YuVq�8���#~ �J�6T��`!�cnx0�s�I0&h�5��w0��d�T�(怫�'���4|-��33ڍ\8�"���q� ��4`ה+W����w@Ǻ� ,t�y<�l���_�f�&�-h�@*����coЧ�ސQA��l`Ʋڵ�g\6��9'hh,��4t��� O��0~��B"�xET��hm
z�Q�E��� uj�����()�KEE�V�H�ŋa�e���bO�s#���_~�e�����p��g�
Ř+���1m�x�{���u�e��G15��"W
��P�gj�����1^Qm�ȏb�@���A��{��(�C�;6�"�>�6o��r�1�8GY �׏�h�'~=��6j%�d����3i�#X3�5t�)7h5��h�����hU�TM����[u��ᅐ�Y^����?C��|���WhOh��Df�fm2�͔{2
�c~��{j�Z/�@���e���Ӏ�;	�/��M4;C>��.����h0�S���VWi�ϯǛ�
���c�]�1��CQ*�l�b{]��^|TX�S���&}�ӟ����'��)��7�!�L��JC\�^�E:�y�1��b���(\�O��t����k.��N�%J|4�4
��=�F����U�7v :3v��0�<�����e6H����/�a6��P�&s�% ����)%�K	 �	9P�"*_������,x��1<yU��^�g�Z�,�k�L�hƓ�ՙc��I�Y�6��Z����UUT.�L(��'G���T�IP���*�9j7\V1�r̂�����'���ߟ��M>R&��Vޒ�P���6}�`�� �2�bP�ݦhp��v|�t�J	��d����MC�*�T�Pq#_Y��X��QE#^1� s�#V|b�U�RP�ED�̺GU?�]�P���k����gY��yH�t���������s�����p8֚��]����̫���{EZ~����/��o�1�����x�'������-=�=��Kt����f�۷�w�Ȩ�3�����=��/�F���wE���SO���Gh��'h�߻�Fr�I�{b�<~������T�غ��c�犍#��b��Y%���ݘ��w�J?��ߗk�F��_����;������gl�h�Yk{���U�������HR�J�|D34�j��K.,���,ME+ͽ(5vڒb�.-�H�h��@E��t"/~kg[���S�$#h�6��ݧB�|}��|!�����ELƬP�KP!ƽȳ|���*�%���f8�|���m�nث[�x)���Z֤�=O5K�vQDeA��+����-���&��ֺkzR��������H�Ó�t�TL�sw�A�r��?���G���֌��TI(���ޯ@!���ajIͲb�\�U���{��D������sN��,mё�o�2&DRŚ��>f��^� ^l�h�b�����r���fDe�	����m�Q3O"Wn,S�~
BR16�5"1���eʕ�l����R=��;�XR��w6��w������Wv��尫uz?E�����z4��T_n���5�Q��h~c��>��O�>h]PkI�ư�v �ٺ���|�V`�+b��>��1R$P�IECN�2�d*�j26�	�A\
����r$ޟ��B8�U5���kׯ����J�s��~���駞�M4�
[#Ścy?6��ɘ�k��ǟ.R*>�aWꥈ?{lH�~�_��$����<�ƭ'�xC�!?	�ސ4D\��q#�Έ���FS^%����u�m����e�ۊ|������
w
M��r�M
W���r��[��if("V�й�FW��k����!m�,�6n�;���bʂ�6��o��q��Lf��������:��6�jH�h��2�<��K"G���t�����K{3�����iOg�ص�r��9�U
��kӈ�ro*�)j�$�߹^{yO��n��%{�Z@��E�.vt�I�ֻRf K�'�V(�SP�iW�%G�����T�Pyũ���zd�Qa�r�h(=�F�Q)��e��	.���=J�Za�Jݣ�����Z~챋��y���)v�
�����嵋4TF�<�C6}+^SZG�+��t~:�ȶy�m"E��AY{��*Z����K��PwrJ�
]�^�xI��<qm�8����izobG&�8d�i���SY�z�D��(bl0ο��@�����׾&��K�U\~�2=�j~�pc{��E1�q�[B�4�a�
Ď׆ؾ�:)�n����Mm�I R�ܹs�	�2b��=q�P~�30d�S�~��5��O�]U~羗kUuwU���%!�0 ��a��8�3�0v������?0���������1�"�5hiI�^j�����;˽�̪��udgV�[�r�Y~�w8	IK�XL�F둎�-�Bؿz���t�X��r�|I
�B�`-�&5�i�Ek�c�MCe_�	M���Y5s���ܨ6�3�;5b.��n�T:�4���׮�m*>ᰑ�`�c$�.,�AFc��W}��
n[J��&5�.@6�lB&%���ˮԉ�4C�n�x�h�����,���Oea� �d�	�	,=��N�?��c��PY,�x��3�Y�h�-#��b)v�8�M���Q������zA���j���0�!��EP30�$@*�?��Q�0 �U����R�±"&���|�;ɏ�2���I�M������/��Y ����p�������8*�{(`m[oѵ����]����={tD��CZeA�fl�<� �I}P����$}���Lu��'Jt�h�I[qm&���w�_R��&5vʞ�^ {
Qqo�5�ހ��'�Ї�>�/�����O�b�G���^�"�?�����M���ܾ���㼈��հDN#\,�M���R`�]���&�	�V5p��f�9�G��b�6n��t�֡���3X�E���en^�!�*~��	�.�� ��1J��X�H�h�Ns�̄�w�$��k}je -F�4z,q�`D/;v�e.�F�����h��G�X�4�l;�<�bd�F|�jnG`F���=�Fig�GU����#(6W,(-0=�~E�4tcA��T����c��?"`�L+8 �R� �o*T�����u-�+p� ���	�m E0|T�Ƃ��O���oa�رcK���GrY4�T\���A��TG����v &t�JA�$EP��6՚R�Ɣ#y/��%b�
^[��2�r��W^��}��;o���-ʿ�|���*}�񥙿�Kዬ�"8+�U���K��O�����U:|�=�m2��9Z��&����:����t|7$eAcBݒ���P�R�<����K&�7_�w�
��̛�`�[o�M_�ڗ����NNO談�0?,"�ڡ�.n1FkG{�����ԇ�����'��=AP��I���/���m���č�9�CS|z�w+�4l<dR�CVLa��I���̬�/6+:^l��y���|H���0���1Z��rI���'U_�u�X� �	m[j`������)}4b���$����صR�JΊ������g��<�) h��Yȋ�H�Y����]&����E�i��g�m���O���{	J&��,��sϘ@N�*��o�j�EC�޸4�e�p�fț��^`]��{�<N1�x��1<ZUV�bЪ�X��X*,�ۣ/ }���:R�h��m8��	['�))"n�V����WPb)HYD���b��*O��\��Hv�k|��gE����y�.���Ȃ�c�sIK�T��Z{�	^-1S�:�pfl�6�PW��"Je{|L?�ۿ��w?�?��os O8n�`�}�ϪBB�y����U��d[��¢�łd�3X�� [�al$��<>;6���ʮ��}D��������mv� �!��S e@/�d��ȍ����n,�1V�������<��mW�gx2��+$����dL}��;���bq1��PQ�r�&��Sk~-Vk������G�x���f�]���5R޵u �
t)j!�gӸ��T!)��r�)���i"��8�~Gc�㍖���|dA9�f(�y2�$�E��{��2�̌+|�]�ԭ��ZAK�I�{ 'r�������)n�5�@�%�}��E�l����Ӏ-}�xeD	�>�`��d�v�$��Ga�1p�LQ+w2�sp�����C`4�'�*�鶸d���������:�2�>4����	��e��j�B3���MdH�i�\h�]B���)0��戭$F�h��#���'��{s=���8������������l��g�
����"�8~v�q�bA[1P�pQb(\rr���}B���#�iI��>�����g��+��+�=˙ۘ�QW{�ڤ�u7*�6���*�LT��x�~���������Z��9�s *J)�5@ �n�b����!�� X
�r��!حҜ���ԪJrE��[΁� ��Wj�钕b����7mO�s�_r	е������uH�E�qE�}� ��A���x�q��$j��=Y��,Pt���5���P:�K���`�|�|��(+d���.I8]A�t�7�L>��4��g?Gw^�ý��!�VJ��)p1)���YE5mҚ�`���wWA�]!���Bl<(&]�X(�?Ɗ��<I��m����Š�}Z����җQ�p���RB�[��K�y�s��P��*�	����6^AE�ᱦ4U!��l�-Y�A\����@�AąF�U�h�xx�V��PB����N�=S�)�#�>aj5d�@!o'�'����N��=I1��Zu�h��v�a��
�=؟�%'��3�6�x
j��������Y8�N�\�m�����M��g�$[���bڍ��K"�u�K<���}���4uͮ�������l��ˊ�suϖ
I����¢��!+X6�s��G?����W�'����u9��h��>D.�|g�G�ܘ�_��v��{~��������o0��/��aAۼb;�LtTN�̣�����gt��,��ȫ�*J�O��N���ۂ	�Z��r�]V+�$sw�MZ���0oǍ�y-�[�g�^1�F�����n�L� v4Y!g�n�(��9��i{� 	IȐ��)�!��b=���~�J���}�V��eڀң�s�v���f���{� 5�������>K�7�R����E~�z��[u��
��J秵����,/<���l"9��,�E��_��Tx[�O	{��@,.sY��
#�`��zld�ãY9=��H:�{�2�VmLO��RR<��.X�\-x�d�B�K,�QM��Me��
�"�����#�J��w>!Ğ=E�c�*�
�Mp��u#(��9�{�ӣ�>�W��h�����*�Ŭ+֛fu��b�VWO��+u�Qn�>h�by�B>$�abJj!��Q r�|��}��aZ�8���-�	�āb mu~~��.���)3�ʉYB��y?׷��N�}�p�f��,Ho_�(\�6�eTz&P5iY���NY�?�G��h� �j\Q2��ޅX�HH��ui�Ȏą��DX�F#��G��c��y�����ܔ;hy�����	��_��@a)Q����"�a�v~�O8cmf��Q��;��8`m,Z�x�:;�C&~ew,Zc�b���A�3�u�P�UǪƪ�ӬmP�bP5n/��2M>)l��Jn\5-�j~� q?��[`��w��s�DPa��V-��T�5����;��4�(��T�P��"����JJ�qLJ��ťq}Ćh�H�(-t�,�diV����4�0AÂ.��-�ӼXH<�����I�K�n�Z�x�1 �d���d�����(z�?-���+������ޱ�2/�2�����E��~��?���Sz��g��(���y��x��֍�.+wբ���=e4칶)[�N�˸�SCP��6X	J���������+�#��9���c��h���a�B懑M d�z���#�T#y���ٜ�|A3ق0�(�P�_����_�}Lp���-�D��u?�p�ulh��I�&��;�1mFS�R��~��T��AR ZN�҈����&������D��dJ#���g�
S��A[�\���՘��A�|���]?��섎|LLy���F)��.�dc�V��T5vd"X���;Jp~���	��)�ՐjPh8����n��K��k�rPP�"���{9�\�*�ƐI��v�BC'�.��F�5�����AM�KQ�R�PY<��E�I9�v|�>
��S\S6a���H��9* a���m�6�2E�I}���)�w���K��\�F�d�I���Q��I�pO�&&g���}J�/*փ��q��:(p�
��PKz|��6�!K�fV0���'4���ا���;˖F<~�/�=JL��
8A+��F�Eo����=�O�o�C�,N���gPBc��aWnM����4#V\z�1P�	�=��oh/��^��y���)RJ�ƙ�ŲT*
�xG\��/��2��a��)�!� �8?$K�v�H�T�!5�J���y�1&ܹo�>����*�|��U��R�}�	t��8���r#����@��\'fC�C�U
��Xr�z'�9[�$?��_���ʬULfY�θ�h��a�9�#�kr=���&U�<�ىB�ߣf��y�6�v�Y�&n���@ALr��%@��4k�lF��eH��+�64��,��Z{M��eᶋ�w6�/̊�?�[v�����}l{Y}[��l�]Ǭ��5i7>��7�O{�u�k���v������h�*<4� �UsP�]���$�KjI"H�8`��7u�� ��Q]J�}ח�����m�K>�g1�u��Z���g5@���܂Y٦�Y܊�	�"�$$��@ݼI��S��/�k�?��:���K:�
ӛYs}�_��|��$����%ŴkS�1�M�EPbTd�Z��s��Y���6��p��V�фF�N�u*i[����ˏ�����&����;���Ϙ�[���\���o�\�<��"J\U��T�f�Z�l�9wP��T �>�/����m��-_Mc<�y���@��[t}v����C+��0Had0�H� ���oX�'��6�?����&�B�,j�l:" 
!�D"�k��*���B#�h�A���sP���A�{�9���q�(ӷ`<5#^�´�b��\�]z;�򖜙��]]	�>��&V5�L��mi�Pg�7m�ܻ{�w������Lpl�깥�Su��&)�6R�Qת�T�\��ẋ�q�|ڭ��'����h�V�"��U����ĵ9��ŰO��t�Hp����d"�,}@��@�Z���z�3�,GB�e�9:썹=T��,c�9��B.�5���\��*f�Ʉ~��t��Sq�5I�È>���~�?�q��_|��fx~��LV6b VD��J��Q�(eJ5�ō���Ef��i/��,+���N��=Y<�=y�9���1
�	D�TK�;\e�'R��A����5kU�5��̥����җ1��\[ۦ�m�:չ2�'�?�	���2���/��sIT=�L���)��B.|v���<{@NWL�4Q���Bb)Փ"�*z���(x��&�z�L�����^��r%� ��ή_�	�my�����#��Hk5h��O�5��q�	�NIq �a�V�k�,����ψ���f�m�e�����d%�>hY�f�^�y�O��ZC���!1�t�~��r�Ox���~�BzBF���vi���r�G��f�u;��pV�R���\q�"p[KZ����p�,sU��R��0�'YH�H5���ZWw0uJZ��|Dn���Sm}W�@_6��̬�"�P��@J	��K�1���:������ﾙ�{�n�ЖFcQ)�mP8a����=����K�/����L���v���7����,� ۍ%=v����Qp�lB+��"���{������m���<���r��by5T}�<��3~���_����ʗ靷ߦg�}�~����Sݒ�P���_�3��P�E�s#�i�M�1��z(������$(�]y��|�y�P��'U�Jo
���11���45�,�8��|���@gI��\/���)(x�R�5�J@2_���N@��h>���c�f���q�u)�*�hjRX��!_�r��X~&t��A���8�����ܝ�y�V�bT��8 ?7^�O�Ɠ�n$��N+�{���D�\���]���z��ؽۀ����
�����J�^���*������}�ֻo�T5�D��NP��3Tm�6Kմ<Ƽ���[�(�!�J�F�5��[�B�7�i���U������-�Y�=���vк*iC�m��6+�GA胙G

�ɸ�vD�d7͂�7�2�w���gi�8c(e0�T�q����1�2��~����>���k���M��W^ᲀ�U��9�o6Kh��]�dF��f�A���zeYK����׮ѭlI@�O@����t�|ӫ<V:����UV�OK��eH���~����=�s����t��Mz��=�5���^֧AI� �P;��UV����ik�ni�^K�J�_��_��IX��V9U��� 	���|?��|?�?�&�2��'���Z2�a�`��ǒ����#C�� ؑ��=t��G�U�W�Q����n ��i>7��!�v2fB �B�>�F�k�ɚ�d�9X�뿚I2=��L>ݮ����|��,k���5}����2a/�2H��߮��z|=^���ri�.�d.�/A��"(*�K�IAy����� �~e�^�����i,�9=d�δ$m��qO�=i\��^����St��!5���tUC#�O����,��fڸo��$�X$ڞ���l�a�l�\O��Z�~*�*���^��xuN���Yhܠy�j���Q�y����׉F����r�6ϧ|<����w/k����|)�xK��H-��5�c'V/���|���l:��͛4��34��z�OY�MY����Y�[h�Qi������x�������o�O��O��?�>ڸ����O��u�"˒hd�uk7�߾s�^��˴���CV�e���;}�ۧ�ً��,��7�Y֐����<�����ܑ�u��,���7�d�;%��R:K0��T|c��7���9?x�Ek��;e��qA���f��8ҩ��h�;�kQ��H�",Q�����wd�6��Ka:��H�5�7��s�^o�ƭ�y�g�n��HR�G��}�pZ_��n=�� ����Ӻ0��|�}�V��N#���0��Ҕ����b���>��,`����Ǉz��j=��ڄ�=�Ҏ��'���R����ǖ���|5)�3=yI���� �z%��0���TYWu]rC�(=���Wi��vq��V�Pp�d'+�Z@!����v���ѽ��uS-�r/�:A&YO�g��뿤�7R�&,�YsRS�h���q�6R��$!A�5�]ی���뿠�?��?�s�O��|�`��jކ:�4�y~Oi�ޣ�j��]��=��ab1	2W+E2�;���8�@�>v�ȹ�M�K��t�-vh�V+���w��?(0Q�p�*��H	�L������=1؎����j���m�����*�dU��>o�f���c�����"�B����}�9���3��A��-WR(��A����r�?{�9�F��ݨ
x���mR5�mK;�٥����M�u����D�|����a,�}A�K�����y�T����B}�w��֬���o�⭧�ȿ�D�0r�c���زH��wX����|�.���`�P-���I.�Ag�\�zm�4R=�TYr$W.�����.6�jbSp�ȼD����w6eAM��8b�I�o�wn$8�{�wϽb�Q�9v\�7&Ѿ�@���q��t��@����_�J�6�h5��wzF�&r�iPX����9�d��pK������p���˟5�TH��/9���4\���&k�H(�E��ں�-�Y�����,�w�����믳G�<p�֮���~�z�����26u����}w�%/��~��2��̺�� Z��3C��d�����ט� c%nL�{YP��A�4�d���
�tu�0�qh������l�6�rX�ܠ�r�/p1�ܸ��}����_(��\��r%u~/�>��b��Uk 4��$>��Q�uR�li���tk��W�����s��{��
���p滽�1�hpwEqw(yQIx�4�6��Ԛh�Vࡖ�����[D�eK���q���i�u�||r,� �:�EW�H�7ޝO���;��\KPH���C����.���YUv�,&�g6o�w��� (�J�}�֞6�v�TqS��Z����5e�5ȧ����|����A�?p���"�|�1��֚'��.�3����71`�����M���7*��F��P����A�!H
��Y�Z3��� V�
��bu���,�V����U�_�r�Zvk�c(��g[�����?�G_c��͛�X;�o(J�S)����?�9���B���B	LxY?4��F����4n�]r<Ο�`���ʟ��LWBY"��`���q�nd��A��c��衘�m%�V�ᴁ���,��l���i�N�i�h��#�Qְ�Y
�TY��-�D��ѥp�i�Wm�M�$Ů7"�Q��!W�L0�H�QmU�-A)j���Ɣ��󢧊��qG_T���%��^�V"�v�g�\&�mZ�A#{� I�L,N��s�X�o:m�m���w_&pNڠ�����i>/Ł/L���%��M��u?�f����ʅ�Ɋ`�g�4iM�xt��J5e�%	�&ιi�d���j��m8�x�vz׽��L��7�|��_��A}')�!���5��l���Ә���X`h`�6b����ԧZ�M�r9^|����.�g+(�Fi~��g�d~�$*����ܜ�j���a�1?���ї���޻�
杻�h�9h��p���Ώ��I�^x!+��E�Ze8�oQ����3w�`�%�/�
�Ns�֗��hQ%e��9n\����冊Sh2-�g.��
�d�v�XWM(���\��X=s�a��@��ȱ`�;5�8Xb�Ί!�naMF�Q��5�f<e�'��@�Z��7en�H���w���ުFFůރ4J��R���|��*�LFT(�n9j`ʗ	���1����T�X���a��Ι�]��.hE���d��-��%����UwլL�wK$��Umb�X�h�8T�ɸS-�U29��; ������'auK �4#I��^e^rqˈ ��
�����4��)��!c;v_(�:�L��&���&�+�86 ��2m�VfB�/����a�'�	:�Jrahu��RmԊP�.Va�dJ��V=B	����"��,C�nJiy֚��s����(�9:z����ݗXK�B�;q�=�P7^.���4࿇P������k��ׯ�����b�"�S>�y.B�8so���CaG��,��$�D��Hg��E�-7�hF��g���-O$
S��ѪB��N��I5i$R�l�Ȃv��I�����(|�uQGm���`` 8b`մ(A�h��Kkn��&D��m��<�Te�))����Jդ�V�.�\�I3;�?���I.=��}�/8q�&�҅�5qOO�kۆT>�=軟 �4�c粲\;4�zL�x��M�[�B��ru_�x�Dޘ3�M�đTS�Ɓ��ɲ(���j1&~��X>����wѫ���|/(��\U/B%�;�p��5!�4��S�,G��>_����.�(!��y����,���˭N����e1��x��n��E�&IN ��V����}�>��9�_�s�6�-K�;U�(vz�#k�I�4q��a��Q��޽8������tp��3bK]r�`�/T�c.:.�F���GS�Ż��_��	?�+�k���;�I�@�)�:ƍ#��4�8O6�P����,�npT�ak���Ia)F�/)�.��5nY�1q0��s\�7��9u���� 1�+�\'O} i?єշLN����5����k����4�T�a�V(_[����ڣ*�����q+��W�ѳu���ha��5�N�X
:-o�~?�z��g�M��>���%?\;��m���FƄ��x��+4�}!'B[�Tج�.�m��J�!Ò�їd=@aI5KMmۧ���"��J�Q)e;�s/�ӥsԑ�Z��Q5����1��~����Kz���8�z�mҹ��!k&@����~��m��=��`��0N���whIx�t���G���e0�f�}�?~r�>]�v�5�1s��� �
P�%�9��8"!�auO�~v��DG�<�"#b,��u��E�v�����t�~/V�nO��x��M�]ǗB�$�s����kA���������f�5R˔;'	�|1BУ�?H�"�N3 Y�Os�3�	�q>�"
 �+���%�䒠��^�����
���U4�V�׈U0�kTSGf,J�q%��Q�|�����"G��\ :��
T����Щ�.l�Ak��~�� UaZ8ȃ�'3��w��{b2��e<���/B
l#wX��G�)P N��H�,��
�]S�m��o�9�m[=�F��2��n�uKPc}���jH��*Duc��)��(�V�N3�[JuL�� =dOwL_	3�`�dr�&��C����F�����٠���Z=�:N��5mɊ��q��e�uO����c��\�vT�bͰ� �������߰�� g%
\���ef��:�p����CQ"��
��.�	�<Ώ��w��E��Z���򊈹�li��s�����w	�-M���oHHh[�. �$w���2Y�q������Խd߫ ��)Wq�
���VQ���7�I�.G-���h}:)���#�&i�[����){��+} ;�;!�R�"+�KI)\uqA�!"j�N�)�I�^�A
�ݫ��3TK��t����/Z��5xZ�#�["�;�#���>�y�HAKF��逭�]JUص�����Ц�$)[���s{u��m��r	�[�F@_c���;Lp?���kpm�{R�ݤ+d@����h)"#�_o����Ia�%����(�u{�=��c�y�S�vɖ�T�(��(��c��]�h?�kby$_�J6�{Vnxa9Klj��AS������P6GS�RG�� ���\�� �f.,=�Մ���A�C��\˒� ��q2�]�
'A� ��q��|���}�>����+)1���e[��j������1�7�m�!� p��Q�czܵ� ���ɿZ.B���|G�� �}Z0W$oS�9l8Y'��!T�QX���I9�\��!zΕ�T��}E+��"{�P�/J�
�T8��YY���*�@)�Խ�B��x�����R,Bķ��
�HL-��U�Y�����tLc�����=g�«�?Il�=&1���
'
)�l��&h��\m�V��P��jPM*�B$*5��*���Ơ�uɁ�[�6�ne^�����"��4b��?�e����T��TSyD���ұ��k}�c(!Y�Xd5De�m��ŊjT 1��b���_h�ͅ����n�}{뻠"����d���#g���Vo/�I���о{U�L1��)R�K��n�Kp��nL�e��	I�S�9�:Հ�i�ɔ�$��p�lJ��b2�5��5���%�:R�*�3/)IXrEv:A��?楗^����uV�e}A�>��ndl����ps�sQ��|v7j�L�I����Yn���>@!pk�k���щ�`&=5}��Ml����}prD(n�`��U����*zC�^� �찾�YS���V�F�4��"Z˔��$~kNy��#v�g�j�f�/��I,�K�(h�C�'K>n��D��3����*�k�A��C�w�$���-�O��΄��>�x�XDh��ܘ	vkּ�пƢ��Ga�<�>	�5�)W�?U!��nB��(���&�Ĉa�Е=�9����jn��KZR��d�'��X�YиE΄���͵v�`�g�d~�"3���{͵�T��T������]4��e��}���[
b��}��x�n3�)�c�c�T��m]�,�c����{������l$!���#AІ�1l�I��Hs���E��_��7�����XēPQ���q���wYMî)}�V�;�U��4����~�!h�����uE���#Ya�髭_:S���u����p������33��B-:�&����5��I�(�,��� ���DA�����B�u�2�Ś�E�=pT���Q�bC�Bo��}��ɠ��
i���l�^�� +�3ْ�kr�Q�c�k�܎�f�ioQ����2�3*�VR0r]�D%��3!5��`C��O�^X�H��&uP&��K*��K���=w-/DwmM��/jZ}E]d��xl�~�^z�X!��Z�������?���ưS䩀ބ8[��zl�}�^KU6�;,��m^��}�,�6RH.8p��������ak���ο� ���J�)��4'ln�.���^[�s�
Z̀�.`ݎ�l�4v�^&�����`�����/SQ���rl0al�V�Z�wiƛ_�M
�Xs�%ckJ��B,E�Z�ҷ�a_:g���ޕ�HR<W\0�m�R-��_#ׅ�^�U
�`�J&��"�t��P-/o:�|ʊ�_���N^����uLq	d�齚;������PM�s�^%�-���It;a��L P�,�Y�)i�c*֠d�k��	���:��+W�J�
�Uʉ�&����ǘ��d�p�܎��>hٛ6�ݵ������}��TAܿ�����Eν�Y�k��MPƯW6�8 �:A_I6t�Z_Bi�T�p��/��O��}�#�
G��n �;E�}@�u�}�F��78w�}�Vt�yW�˶S�D���k&�dJP�m���E�.���9(���&J�)R�����F}�fj����R��4��al�Z���̉���g�mW֚7�!RMxdWL��>_����7#��d����\6�RҨ4u^�A��Z���_<�c��E��`���̪�&�V��BT�g�A4��,�4�,Ƣ�x����$��|���Vz����ȴ�e������M" ���XS��,-P�o�-m �"B޴J���T��~T�HrQW�,�����7����VF6�7܆�����(bR�B�wk)r�#�_,�5�?�lD�6��u�㧒��ӘB��}�+�oG����-U��,2U�8�\M�~�����9=],�Aя`J�^'����s���B���.���4T����K:�6
�����!Ϗ���T��v��0R�&�T�/!��q�\�UX�?�t��$�k��ʩ�7�lh�n/v[-��o4<�4�w/A�Z��y�右P?ɯeq�4\��u.[lD6��Uê�DKp�}@�
E2�	l��dP��ْ�e�ܶM����vkNU�E�9F���,?�dF��c�nʹLNc�*�I�wR���Q&�" �!�ݤ�	�c�.uܳ��(FE�vCA�K;��h|E(�����aT#��P��p\h�k�V�t�����rװ�F��4W��
�BM\�/��pѸ���F�U|/2Q`�Y	��I[��v�R�A��(a�@k��Ҫ@��8����	r�yj�$��Jᢦ���d6�l\Y�ʻPH�����eK,$�7E��_�l5�=Q��-ρ-0n<���w�g�̮�[v��7�
�u��s��o(m��J���L�<GQD���\P4Y����� 2C�s��or�<J�	*F�r�.B��0����C�7ۯh��ϠM��]�)��'�$���V�8��yŃon�٣��R	,A�����E�(>�	$�TJ���	�Z����G�r��I6��O:P����^ ��Ȍ؀`�@�V�3f�a����|��9\�@�pDoԿ��>�p��F8i�� d��[X�&�g�<�m���Z�n���$]�����M���-G��r;# �rb��]vC�L���R�����>��>���F D�cs%�e�e1R�I���6߳��H>[^���}����A���;튽]���u�V�Fx�̯�X~�����~�6$�,z�e��yK����w��Oc���9���t���g�LE±�e�G����=Z�/X��@��ࣺ�z-����Q��eP�P�Z���0uc;)��2�-��[-�KD���	an ��}���,^&��M�p���Lsc���5��L�8f���ƴ�N�᪚L#�	���}^љtJ]���*�� a��A�J�G�k�|�$��gϓwӨ�#C�Ao�H��m8��1�g�,�U�_��r�F����W�[0�3�ɞ+��{������$pN��Z�j�z�v �g�2I�<R=v"�,�X��B�˝�k/�V9/���	��f���� \B*`�Iۛ�#�YQ(#�^w�X��ؔ���f� Cq� ��Ǥ��d֧�"���V	����+Z�`c�pӃ�������ꀽ!M��e���^4��b��)�W����[*�?�������?8��d%�ѵ��k���DN@�@&9�a���X�}דn���E��v��\�:��<�`�e`�M���/��(kŌb�2�]� G�hQț��?��
��Ԛ��X?":{̅u?����E5hٻm�g�w��6�����O�`ߛ�$mل�l꫸e�B*�vu�S�6�d�}���)�>Mh)�]�:��K?{X+��:�ܨ�����"�$���W��8.=y�$�<0��H�!]B,D�hȴA�6�&�w�=n��sZ������A+k�OjAJ��8�l��=�h��ц�m��%Im���.��2��|+nq���CV�O��q��b�=ݮ�Q�]g�ݐ����
����-2��(r��|�Fk���^��-�r���ǫ�W���7fk�4э��.\1H�fsc�C���ߥ�7orɻ��{�ǜ���3�7��g��m44��Pn����A��_^呷��_`k؄�S�������C��o�EM�<(\;9ȫs�T����"A�{�X(d���j���gy�>��i/�h{�}u#U��/�V3,S�����O���$@:�("ڞ�C~��;�k�`��+��r~u��#mk�e?��@�lc���ш���h�o��a])$H�Fd�^^,�y�*ZZQ^4_�	����)���nЯ�\��mCB��8ߥi��
H�q�؅��cK�ٙ햐��>
5c�lT���*`R'�ǈ�'_Yk�I]w��G���7�oǴ\�u���ƚ�V��T�9B(�4N��JƱK-��tF7�Hƍk����0�cH����`���0�s<׭[��gXb(V��h���6��E�݊�4ۖF�t�|<���*Q������3aWL⟺�W�Q�J���jI��	�4ǁ�����f���_)k�M�Ѝɘ��<�S�Fw�`�8�&�׺��{T.�n^�AG���=O%ñTH���N�3O���u�Eg�=��j�F��j�����Iy��Ķ'�&���0tU]y�ۿ�@�?�9fy"=s�Z��RmKS7�ݑ��Ō4{1F<(��eq$��k�
���]e��{�:��]�h�m�	.P���Q:
n�	��Yp�hk���ea����7���q!h��?��ڦ���q��~�&����;f�� �V�����ۿ�9�.Bꅧ�?����t���n�t~����?0F��Fle3q_V�P		Zy��'�/_|�e�♰80��Jc��O6��dω^��a��b��s����n¡����y4��� HM:��S6��pt�4K�����4��A�D���1���@_�)���
P���^���z����Zn,�6�s�f�g����!�t(]���7�+�8��ޔ���9a�.S^��g��UkRs�H �[/Y�A#�g�^�V�ddw���)�f7z�L�����H�"�RILY&Qޑ��b���w3���%A����(��ĕ�]�/n?uQ]U��|�+��+�;�S�O��Rv�������'دp�>VMm3�%e嬙����.�l͟?�@����I�&E�t��J�}t�&'(M��m�i+�Y��n>^��WU��m��!�'̝��    IEND�B`�PK   ��xX�@M��  2�  /   images/a83bc8df-a6df-47fd-a18d-828755ca269b.png�y8�o�7|[�H�"di����Ki��-ɾe�)E�%d/bb�%����c�Qvb�c�����<���{�<|GG�q���������u^t����� A�ʵ+���h��w�'<L��{��q� =%���׊� (gP��%M��߽�����I�f�rͨ�����6G�0.��3��g_P8v��l�����+��8���O�':�ٳL#��/Kc_��\�U���wu~�4�@{\�{c�
��=j<]����˯�U;vj܃H�d�k��ghe���,�UJ������/84��!���Ϳ�˂���xiSSӊUL�G�����4q��w�ou4����7�:V���So������!u�ݻa�^�n��I�Oed��A���h�5�P`��[uG6������7بݠя�Ү����d�2��W~mcy��ˣ�a}�%DE����"+���G�'vmu�<Ƞ!���O:�G�'r����P[�<f��ׁ�'����Ms�V��iE0�?G��!��|�P7O&+]�:���h�K|DC�.��Z�,#z|{��#���u�E�O��Ĵ�H��WU�+����n�/Xo�pgC�J�8K$���b��m��
Y61X��e�_�ɫM���J�����S�>\؄=�~�޽ӏG���͉��D�t"!񕄮,+��E���h?�����"�w�ޚ�x�#�b�H��h�u ����u�K,�%��c�4�_Uuכ��Hӌ,o�f���:�T�[�����b�1~�G�/�ǟ>}b�7�e�w�Q�j�F�wO�x�ެ�_����u��d}�gL)�,XPY�R�K���<�h�)O�-��c����S$j��pHV�0'��"��}d�m��n6M���^�N�v�poi�c��m���\���Ϻ��u���Kh�{�\Y��B�����֥�~�q������K�y{���l9׶�?~|ȥ����(��얰�����}b�}����X<<��zm卑��;ʉj���S�I�@�3,X,���̳{I��O�un���Ȫ�EG�<'XK΅��Tr��j��f�}���6T3l�\��I}k��~Z@y��.����;S�PM}@;߯� �lH�IvBؖV,���1x�y�FR��ԁ�t�A<~x���.k`�̱��l�P�]k���+S��e��ꎿ�?�Bl3%a���/����=�H�i��O,H��V��z`����%�� `��`�%>V�ANZ���i�51��.=4Uvv�::E����?FXS���ZX����99] Z�OI�=w�-��}y�����ə��Hq���bȡ�<Y��>�U���*<��q�Ϯ9���o5aެ����8�@�x]�K+ 	��%#�`����iy��y�B�o��R���'�X�y��d���$���v�Tݛ?ћ��=�xps��g���ʐ�w�1�\Q�呣w*H��j��g��d\���9���t7�����J�/���{���L�G[��bL���3��27��x�v�}G룆�\�/p���Ő1������ N�#���f� ���Y#�$� �˒t�S�s��LX:���,�(�5��OHl�c�u��;��������GF�y��G;�]��x�bf�}�bځ����g%Lnn��s��ߨH<�@p<��%^���΀������^�~L��v�U���y566�M�	����G���qX�� P�j'�9�v��6�W���Ivy%��,7����aڟK�l��X�(H�Y*��L��1�S���CP�8D<}�`��|k����A+ڴ���T��Փ�6Ω�b��>�Lק�����V�K{�̐����RܫнHc��K]]�xtJ��;�,���4p���#K�+�����W�O��|1k=Ǚ(�Z+�f�x��)))�XHĆ�a�w���t�^s񈏒J[����0Jl���\��{+�\��Y�[A�+��8Ų�J6ES�j`sK�ðڗ/_L����v�`��OgɊ�c�i�s����[���ߘ�##�����RZ�X�����c����������Ą4�~���2�{qq�E
6YYJL��Hl��`L�pp���w�ڦ�J��ϱ8�SM�5^ͮ�G٣�.��u��0�X(����ٴ>��:�Y��)���EH�����>k3uh�UYx�a��I*^�=����(š��������ރ�>>>�
��Պg�E�Y� .ZI�N��\B�}�p'ҿVMIb���j�]�!��9+ǵcb!K~y0��b���:��o���fQ�nn7펲�\�e��c�l������������3a�+���s�%e�9,j�ֱD{{�'{��5Үē$���<K�#�;�eH�vwrr��_�Ԕ�⯽.�F5eU�(���H=v����e�Lo%���k�����/8�<�%�����[�s8�WR^m#���R4T��&u�	�����xx�
OW.Wlt���'o���󣛾k��}�n����>�m�Ԑ�4�&�k	�Hi��*2�_���1I�s��D:�L�N6�Yc���5VRW8���Ȫ�������N�sl^ ��Fc&������z�q���g��	��4nw�$���sMiU2:��z8)��$��D���;����y�Z�zlr��mps1��
j�Y���#���4�Y۾.e�{D詁�I�Z���H��GH�������ĢJ�e~�)��c-����)��7攔F..F�� ���$�Of_7=_5�,� �ߢ�r��iI�W/�������n �R_/^�7������o�8���<�.���RF��W>	�>�x�=�(_����E��O��M�pMs��/s����N��0�1�vDBJ*�._�5/�|���ي/�U�I^��HkOsKKCM͕��{��{O��/w*$nR��d�ͦ	���A�n"���t�$��>OTߺ�5'�[�lI����&b[L�F�A�<�ҧO����K����%�ɱ z6[��8�y�Q�V��`�f1raK4ɏJ�8�DwQ����Uz_�Dvk�Dh�.s�Hd��|^�Hx����(��!*��/_:����GP�ٷ��b[���!B6�E!&''�E]�v��}� ��I�DD�ڎ�S��?FGGp�t�te>nС�q� ?�8g�&�k4c��p��#��F,��EN��;=HW�>q��������K�����Q���Z�X��]�e;ƌ�y�z6��y��Zx1	L�)��j�>�����ז8�npkgV��	,�m���Z����I�"`�TD2!6=@�A(��v�n��ZZ�O^p"�\U\�P���@��[}��[\�|¨��e�u���=3�Т��XZ?�0�����[e�f�ܮ5�,�y{��ي �Vvs`����k:&ff;��F I�����LD������?~�uf�b���?��֦]�����w�`������Z�N�S�V�v��y�wA�Ǒ� W}o��H�L�PA�Qcc�<V�|�`,�}��y?]�b(
�W����N�مL���略E��ظV���n` ��Պ��5e��;�Ji�s��4Q������������O�����B<:�+Hao����@���hg���z�d����A�#�@�N]	��� �.�9�<t,���(��I��F������A�Lٙ���#��n��x�~G������/��s056���r>��2�;d��K�SE����s��CYIR�S�wOq�YAv�j��ާ^��D�4�)rs�Y���L���R�i�o�ؘ�lB���VK�*���(5�;,gb�v����$���떺�H�}n�{gL�v�Jp��PR��!g�O2s����` .}��!؄�4S��i��*X�!�=s_�=��W���� >����ֺt��_K�%��h���~�5\Ʒ=�ЀΩ��l��脄ȴ��9�!��3tVx�~q���;���C�Fک���{������ i�cɝՂDjȡ+(�5�]i � g"��K���nF�>Ȭ���Xk^tČ�8'Ѿ{c�c��ĜhF�`��7	w�ݿI�{.�"�R����A`ҶAG����8��g���&���5I%;V2���[�291��S���ɬ/��Zeڷ����kڕ�8�E��)�J!�H���zʫ�|�`�m/��U&���[������La��U�օ�>�i��8Aߞ�<�(�l�׋��I���BCB�So��B�Q�&I~�7��}Z���1�Pj?V�p��V�* {���`�n:�c"��s��n=����&1��~Z23�[6,L�X@���JFFF� *H��V���@#/^�x�3�(�<F��9sR�gy���p�O3�s�hR0l��Ҥ����뢓���]~�ctf0�xק�555��V�c/��N�홲�&2� +��g�{x�<��s)�v5�U��^�{o[���ii.���V��i� �q7��"�AU��t�A��� [�G!	���'�z߿�l$~}�2����?{�[{V�W!���I�(�"�� /���<��d�������V�}�����t�~2ٍ������ܜ_|��w%���{��D�(�K|ͦ���4m#��ͪG��|��C�B~���Ƞ�=u���)xy�N�u�Kf��p����f�V��oF$U�G
�(hj��BV�Y�W.Vԁ�l�#S���&cC��Q��oe8�x��*�������y��I###��El��	�勥7��׎�w��S�`bb����8�Է�\��l��"�Z�	����ݓ_�|@Hu���j�(~�~z��I��)|~��@�q�~�MzUr�>�-;TG	J�=��o�&��$%
�#W�����7sss�b�]���݁�� ���fJ*6`j``��t�i!�R�M%����]�yy�l"�������nڧ��m&~�њ���Z��-�����-4�Ikv�����;(�����z�(3U��6���A�@Dn�3/K5���߹���Ձ��\9S+,���	C�,�=ǽ�}�r�Vtpy$1lJ �EA�*!ː�W��,5$R���S���z�
�[F��������z�x֓�FTގ��$/e��^�w�����̒qA���&F~��`�iy�gs��5�l5��M����.�R��C�I�	la��(dD�[uݗ?�{�J�+�)��ӯ���Ӗq�
ٿ"�����ˣc�y��5$�����ﳂOl���;�7��K��]���Z��L���S�����ח�F�EC�m�f���C
���񊊊SO\k?���p,a�n��W����p}��{�+(��Ⱦ�r}��!�rm��I�]�!e\;�4�*��aC]����ÄӤu����ULMMzlY�Qq�фn�����`�ɳ�2+}�s������--��q�=8FG���D�m,�E�.,6��ܖ���2�)���'�9�k캡��o]�܇Ji�	j��s�*��D��{���ߟ_<�{θy;�gǲd�.d�R�\��nƍO�>7GuA�y��V��b���4������������i��)A�f�����bוui0�D3�)�:O���V�c������˯v���S^���R��	�޽;
�W����xuy�nC�D��|+{=�p�X���9GG�Y
��жbٔ�/?I�Goۘe�h������x�H]~�})e �J�Fl�W]�_�WG�Z�|/�[�4i��N\�(�Dǫ7�(����!`���a���ȕ��C&�35��r�H�Xb�:��!�V.�>�f��h�O��F�|b�Oj(�mZ�2�J,���'��K}�Q	D�	����-��Ve�������أ��٨檱H���e�<��˵���Q��������G�
 �\z���v&�v0M+W�L�۠�t�5��=~v/9����x�ƍ3+s��Nx�ʜ1�6c�2���׻�Y-`�P=6%`W�3 ���w_���a�u��zwj7���������I)�>zZ]F���硍c�~t�W�.6a1���ዓY ׃7Z~8�}9�ĵ�8O��j<�TE9�g��X��t]���MIV����}Kŋ?���S��l�]�+��/˫tؙ�׃,O(�ȸ��;�4�|@����6¥�WI�VV��9B���H�[<
����m�E�������[�����<��l٪έX�2��M�'n|��8Z�2�;0he�ڝ�)�g��PI�(e0X�b	|�XXy��ץ'��
��3ÂZ�d������)�P� ��>�-=�^�\L�]�/\yk�}kk����'��b_afSU���Uc��w���Y��Y���SK��Rd�����L�h�s׃�� ��3�,�U].�]-Ԧ�!���8�Y�%l�Ĺ����e(��6���1��l�B�dB�I�CE��`�W��b��N<����p��Tk2�,��{=6�$o�g��������}�C����y�����APra���w��YM�U����[��U�},Rr���9�@��ZldL�2Bz͵�����Nא�}6Yq����e�/� -\wJn/�������h��ĕ$)��|Refb��ా<�lW�9�T����`��b'x��}elLu^DvH�4��HՓ�����B]Y�����ò�~��?�z����O�o�d�'�d��(�R"q��AxG�d�#e����U.��i�r�j�_D����,!Sh�6cB�����Ǯ��+4ؓ"���kVsIY 0��}�g��=T�6�7�&��ey�@c��t�*2�����d�0����P�>�ȶ�)�Wa����S{S�,��_��a�?X�Ļ�����O�M�k㊑�\�yf3A�I���仱:$d���W2km�4�U?����c
7I�,����
���F�X~M�,�=��{M�ϯ.��_�W�b.<٘	�&n���j�X@O�88^�K�J����o��'���av��\A.��s1�6��'�s��Qe�jO��K23ղ�+Io5���Hhoui��W�%���j��m)Q��+�~��]3��F�-�����vo���E��mo��T^�0����R_s�U�.�̘���.j{4���9�J�$�O��U=j��|���=����&&��Ls�qzo]������ole�Z�ck��/g�����8�g�H՘�W��E�X���G9\*$���Mb�o;���g5!?����x@�(�Ñ	����L<���4���p���ㄡ���j������g�p���t������#=��g������e?w#��Ka�y�5'���WN��4w��32PL;�֫n���|ã���KҴz�0e�E�IH��ڠqa�^�P�$K�}-���^;q Qm�ʧ4�G&����p�ƽ{�~�	�����Ync��Zs2��c���LoK=M�M�<��k��ﱚ�L���tL�s�S=���Ǖ0��G�����C���0���u��j�዆~��.J
�Z��ү~��QƧ��,�w>�P�+�]��H~cm�u�W���݂�S��zK����*a�ONu�����ui������'�e6^N+���z��d#~���1��^�}nf`v�~݉�{��i�ML�Q�L��ӗ]��Jr��}pP�Dֶ�׭.E1BP̾�:�Cvə���`��w�j�t���n~�����%��i��dTOx��:�V�k���XE�3f�W�U�Xm�I�uNZ�޽�C���V�	��6R�F�ʂ�V�0?� �+ԠQ5e!#�sڠ܀�3�4un����S��@�a��-�w��Q4Bu6��˧!\wD�{�T'̾)F��~�P�ǖ�j��)��)��dg�5�
�+��<SP�g���尟J���%^Z�c������5_'bo,��@#CW��|��'1ʌ������@H5��p��4rxF�^$H��T^S���D��ҥ��W&�M�a���[\��]55%.w�ܗ��,?�أ�؞�u�v��v�wi`�'��1��&)*0i�ʳ�t���	������x������ܧ��-lm�D���^�<t'�S�0��q�J��l"�С��!٧�@�B��i��^um���|^԰t&���n:�߿���Ʋ���q���܌ׇWן��a��b��Ģ����>NY�_i����J8BG�����O�r�ј�/�i,�jxX�쵅�޾L`��PXn���K,^_�|~��xD�-[c���Ox�)����+�>�Ś�^���]�"^���}��5�� �Y߾�U����� V�jh==~�[�DCNK;-�H�&�C�?W�g�:�Ww�+�~]�%k�XEKll�����LK��]ŉ�a��Yd��_��O�JH���:%��'p��մ�@r%�v}¥��P)"U�&�|�/��Q���ø�:�������ZQe�����ӑf����訇�랏��n!�[����Լ���GZ��?̦����' ��
�Y��νZ�s+7k	 ��K(���b��&d���V3�N_<�Y2c�4cKe�kv�b9ܟn�y����sÍ�Do��ʖ¬
]���Ҭ#��XR�n�������iu��'k��k��������]��P*~�s��<��T�9a�i����w���T2lZY�}��Gqs�,4sL��P���#�<7�KO�� \\��Kcm�������D���j�:��^?�5T���~*�1N��Mş|]�\����m�B�">[׏~+tP�~10�����ݫ�p|x��G�y��N9�i��ӵ.88=L�X}Z���\e�M욵�Ϋ�) ��$$�����{ս�H�%ֿ<����ңA�V:*��|)y��$��c������y�.��ERT�{|�(�����j�~����L�܏?�7�c����*k�|�~|����E֬,|�uFr]Ϸ\�マ���WO ��9s#f�lb�?H�����n��9���A�p��E�����ʩ����@<�'�o�W�M�RT�F&^z��N�T��~��O�K!x�~L�M]��x঳φ���~��w_�j������
9K�k���0'�3*�Q��`��p9It�@Q$7\`G�h�1mM$�r5q�'s˜�A�zp�9�M�b�]i�r]��R�Q��;���}�aF�UK=Kӷ��LgaQW�C)�򓳔A��`J�|=Z7�!��d=`��Um!(��v�<[%+��t�f�w�Na����WeE�E}'�Y�W}ks�&�J6=T?���+�U%�[b��EC_|�'\���r��< ��T\�j�!�\�"QOEjrl�bߣ�RT������I ��QG�ˎ� �H�.�u>��/����1�Y:�x<����3��\v��r��4��"/̷�@�Kʟ��璴}�[ꪌ'��.^�ny�>6λ��}���SQ���:��TG�.��I���=������d��K��7�J&���ȕ�c�����N�+���BϾ��a�T�GZo��n��
��e�܇�����>XP1�Th�WB�+S3�
-=F��F���<�}Ƌ<�8d��$�;�� \�}��Tԃ��3�L�WX�F�߹۸��j&tvv�|��^�Ƶ2��t�@r����g�V6����,X[oMvhՈ��W���{V��H�N�>��M��n�vT�2�H��z�A�x�AhO���?�&�-�ŧv0˃k��s oB�ƭ�Y[�gk�%w������f�12��	-:	�1	o���ݡ��Tb���� ����b<������a2�� rk`q���Z ����a�T�éOQ�)��x񚝍M�I�h�F���<�q�fϧ6n	I{��%�ߊ������ɂ#��^3W?��=Aw4û��FC'��5�ܤ(S�����m�2Dz��u�?�)�e�zx|`���g�#���$i}%/�
�WI]r��t̾M��	��N!�s/����񉉹��&b����>cs��4O�63L���gq�3��~�<;$
wF��6o@���{]���'r�����}CR���/��Y

sR9��KV�d�z����"�p�P�HDK��'Y��H�ƭ�b4������s����[J�)�9M�D�?y�c���,��7�t|�:v��O$�����b|���n�gu`��Q	��b��4Z9�f!�@s�Ҋh�X��Z�q/c���xo,��K]L����*��~�w�����T@�.Ү�-�du%#֣�q�F�o�6����H����-����sL8B5!�$��93�9u!K%ޅ��!����ϯ����?�ʱ����[��'��#Ezm�;7���vp}�Ϡc�y�'f�9V���p�ḫ�7�*=�lNm(mi�Q����6Oi�z��O.�m�iT�*[ed��1�Y��w�p��}2�ߒz�Ӊ��P�a��}�Hz���@�8`kkR�}���/B����M�'#+JΒ	%LAe!^����샴ӑ@�Ŧ���W�9�?��b�J�p��_�R�����p݆�ۨ��̓�(~�Z���B7�>ĥ�0���]:��n�{����ٱ���I��E�?��>z���lg��L9r$��͊�d��Vq�&�f�K��*Aa.�2�2��
���[r�������>����٨�E��)����0�ơ�ڧ�auڵ�9+z��C{QT^a\<<rY��D;�y;60$�X�*���!b�F���M�P-W��U�����>��o��%$�~��[̘vK�ya�=A��?<I�=�5��E�j���Ɯ�G�Y����w0�����䢋������x�����f�БdIS�3A+@��Rڴ^�<�`N�k�8t��v"o�WK��aA�c�,��Τ��~E�����z��j��! ����������1�|4�SD5]�v���m!�n���{��*�P������?J�0�]FFF���{�������S0��G��o�_��贲�r@Wz@�;�c�<a�G��
/XP�66Ff�Ú~�-��5��vsJ�L�X��;���T|G�UĮ/mm|�
�:؜x��G9��g2��y�~8���ҫ�E<5��
|ܕ�)M�'�6I[0"��N�E�T7h����oq��u�~H��;�}�X��gx�$���j�h5%.,�8#P-/BB������J����[�,⑀��;Ԑ�3d�<��c�Ζ�}E*EvQK|��*¬=�Zj�k�=�Yj5�����[��U�/I�%���M3���wI��q�ԅ5��=}�~~@bF&+�'�l#$e*�^�]dɞ�G���H� �;�$�@�x�
����ٚ�S�2ngc�wY��Y	���q�9M�uV\k�]���l�t�h�1�-b��I� ��O�e�ӟa�nO�z�Ɠ_�M���Sҕ�!�r�#��4����q�%����%��j��T�ii�M��	��'�%$�U�N�L�O�|5椫����E��ˋ$;�.�D|������M���ˏ����1Qݳid�Ш[�{�d�u:�Q%
��\�*dfM���1�z��ߕM?�"8~�!�����>�9���80�����lUy�ؘc���oi�Qڧ����B Aj޺�� �<_�a���?�^L�Tl�\���Y����(�K��)I$Kï��_[)	X���`�ّ߿�*���m��}��C���w�b=��૮�1Jp����*��Cg+� �T�P�l��>.ƃ��%�.����]���7I��a�����ؿ��37}7�;���
H�|�����z�}S���2��8���W��c��洹44B,U��_�^����� P����b����[�	'�z� c��x
��H,�V��R���5���+��wQ� 9�U����}`�P9���Z�i�p�	g&�8^��)h�'B#�ԋ�Z�+�x�� D���*T֗!�H�%A�ǥMO'D�Ơ8���z�q}�M�3>tR��d���vV�V��j�(d}�e�d�Z��=�|�f|ֆ�A���{~�}�����@l�C��R�G�s�i�0j�_U��H��d�x����
v5N�..�9  ]A�mC>����l ����ۤ�Z�ѕ��ڡ�|5�x�x�s/}*��7CaiL�x̛_H;`�u���Z��3����P�h�������/�<�5v�v�����dL ]��
h���+Ԯ�1��fE���� fm����]evw�}4�zoү��*a"TO�x�xW��l�7MS0.��f�ڀ�z��c¢�̱�g�Z%��*��ޠ+I�DbbːrDzs�r�&�P���!�����5\�v2���q�p-���	!'CQl\��q����IUWi������v��3[G���fe��9u�MD�e�g����g���80�_���tP�MOO�O���]�;N�&��XS}f����\��f��4�v�J��rr�P\J)w��nDw��+��G��&<���zW�<d)�|��)��+髧ix��f�S?W����� ��j�����jp���h5�"o/{�Je/��4��;���>X!p`��h7�®c���D+�>��U��5 [��=���7C��h<����E[SS����=n����h��Y�v�;B����ǿW3�[��6&mװ"��#�۾R�Cx��zo�8���!�lY?}��^�^hr^^�����R����
?U�Μd�h5�/q�/��n�r �F�2q"�1�?��cW@ +7˽C�ob�mgdH��w�P��6/��#�D�|�ؕۤ?�\�M��h��ߍ���R(��s2L}��^}��-�q��Q.�g�bR�Sy���� ���~:��^r4�ۍ��+5~Ǐi�թ�VN����/~��j��	���/���4g����"|�,����ڴ8���n�guq�?6�����Pl���"��+Q�I�~�^��A�E�6ϕ�5��o7�z��e��l�ף:��S}�:R5%�!���u-�z����N1!0�h`r8����?5^Q�����ԣ\������J�z��xC�0� E��߿3��%C�@vӺu8�����T�˾��k�BnվT!�0n)?��9��K���zHX_��a;����*��۽{�U��"�{����Y���^~�bS�
r/Y��Պ�:���*�?B����N��b����t�Wy�
R<��}��� ���5tt���Y;�I��tl�T�/˭R�|�˱�:X�IQ}�t��d�ӧ�z�4����&)c��J����[K��b�Ch�����~��H_�)�\vc�D.�BIs��XP�K�Y���3ͥ6z�u�H���|uuY	����9|��h���
r33�Z��%��v�*]<0o@L�͚nmC����j�4���F���*�I���f	��ق?����8��{�ȏ����Cn��{C��Y�Ə9�v�y;E<F�O` �6�ƍH&�÷��w��AnW�e�nP�|ޟbZ����b
QNg���Jئvn���_JѨv(��*�(�. ��5��ojL��pa>��~1�q��ߋ�����G$tAB�J�h�Gp�F��&�~�<�7}w|/��Z�f&�e� ��2�)20V��iOs�o��wpJ�*�;�����R=�(���&�ݓ,���t~w"��*[��%�vZQQ��h[(oe0J��dTV��������G����u[�fꗪ���w�O:����0a���v,���KC4
s�@� C�)��Q�N'Vo�V&5�G���w���|�������\;Z�@u��k��Mcu͟P[����S������pᇿm_�}�!���iȣ�kZ��w�E���Mc���J���q�}�f�
��������Jf��ع�8��^��A�����9iq{+�4��F����l�K��� Uޯ]79��Ḣ�3�Y|(+ �w��6�f��u''~���t�/�ݲ����_ׂ��Pr~��~d�V4�B��l ]���ֆ��D5n|*˖��9�}���j��p#��饉�������'�L(g���.�0��~::�,@�Wep�?W%��D@�7VB�?@��S*��7n	�ӎ*ۓ�5Ҝ�t�X��������2�H��2B_�Y��)�SC�ɱ��?����eڻW��iP`ŗX�,�I\OѸ5��}�֯��P��e˻n���$�H�ʳ"�#~J�t�1�> ,9��F�t�����(�s!�Wh�U�[�F+�~9((:�#:..��Ai+���8�^ �js��_.)
�P�Ɖ9��ޛ�Zb���v1��K��>�]#{��0� �/w�RMAnɺ���%j[|�y��N�����Z}�m(�����m@AȌ��?�h.���u k�����A��S���n�{��#蝻5�=�1���[��E�T���qT��!��v�g6�� ?�y�'���ύ�o��ǝ�n5�P׉T$��X��y�L��v>nyy����;�TMA��������`���Ӧ1���No=�3�"�˺�W�@.��G߿}�w��//o�q���ڙHUL[	6>�܁�>b ���Wm�D�a3$X͍#s E���K7�Y�����Ի���U���^_�8�y��]^O�Wk��NA[XX����}�`R3
��=�N�:�[��&�����ML�����ѝ	����b/�g���>4[ �};2�(�,���?b�+�P���
��Ǿ�xG@$�C�v|�&11LЬ{��3sGU�?�A8�9(I궃|�_�亜����/o��HzpwjH��Έ�I�g�-��>8�P�d��D��[b{���~_"��C��@�:'k�����`rٖ;��G����B��K�Ɉ2��w�옝��1�;<	�N�H���y+TԶ�u۟8x����95T�g��1 O�'��T��ظV�䏺+O�>�&�>���Y�s��~��w����G�>~�� �3;ʹ�y��X�_a4���&�
�\�1�shn�|��I���
F�AT��Rxa1�������y��P]�%�����/�\��rJrH�H���=�����ii�<\i�A�-xGP�&��"��훦���)d�ó=���n�!�����!��[�֍�.-5�p��[��U��d�F�wF݇��UTUl;�B�BPh4�6��C��׆뀫|��ԙ7��w�&���a�6��&�$')c1 �"�m}TQ�#��PO8ؓ������ u������u<�~]A,�w7�q(V�	�G&�_���C��%��A�'�*bJu��6�B~BX欼����]ʬ���]�D������[���&��jz�N���;�6R��Z��*e�n���/��ǵ�|W��*��Y뵴ҥn����.[�Wb;|7��T���t^�ء:���5��r�~nt�-uP�I�ۯ�菞x�M.Q_�s���t5N��E�V�h�{@�%�V�n��$u[^K[����Mo�%C�B�F��t%�3/.h����J��R�8����|�8�����J����3CR�a�ҝ�Y0��_�D���t[(k�J�����L�Ȼ(�l���w�U��<k [�S��]�4ӛ��b��,��t���/8i����S?��ڳi��&+�c��|`3�|�ji���.��v��<����j��	����ͣXMC��7��6�X(�B�wf9j�R10a��!�缵]��&��!yZ��j�zl>t2�s�X��H:��O!8�6:�%���P% S�^�L�?qq�\���v_v�df��F�pI�`ie/��ΘA�n��Sa�%f��5�zz��}.���W��|?J#f����9�|����(1Ӄ��V�Q��y���+��V�C:�ĭqî\�pj��p���2�t@2�8���$q.��8^]^�hX�ѧ��W�F�����]�-�θ�k����z����Y��4�~C����)��ު�-\�G�F��r�AȦW@���[�G̈́����X�8Χѷ%�4��d��m�p	���=!���^�^�,�oE(X��_V7	���2-9v*�����{�o'�㨾�¹�[Ӽ�a�e;��?�}������
<���:��>��ޯ�:,�8�D� ��b��u»;�b��W,�;u?״Y^�wB.Nnu�Q���l^�ZA�33mҹ���C�k��ZA���֝��xȷ�{�߃�����_���!q�Ǯһ�'ۘt5���S���]�� �4|	�j�*� �>õ����8?h����Be�b��Vp��eg��Y��_��3�R929T*�:��	�c)db�$C�T��:\����R�g�r�m�/ɋ�0�,	S���g�K����aÊ2�������*?)֪B���;C�$w��@x	��x��%�R̋W�J��P��H�v�{]����>�?v���͵%R~�56K�������o��W�K矐�Wg� e�t��m��Ʌz��������]:����x*�;L~�LiU�Q���C���6�c�L�o����6���� ���#>_8��}�Y��ȡ��ag���T~%,U��Qz�E��`�xT?��,�-�v��Y�x�MZ��5��T�	�M��+@��y�]6���Ҿ��[1�6���ݽX���x�:,G�.��x ��P�Sn�9����Yt�>�`�yăW���|XO���.�����o��g�b�1��,wm��y�|�C_�Xj,�ʋ'K�۴-����l��񭝫xJ����t��v"�g;��G���DE����Z�0K����"���� A�=��_�zWT���o�u`�jC~?��_��=����{�߃���� �MK��i"w�ʝ����ɷԺS���N���8�0mzs˥י�q(�n䙂Τ�8D�Z�6ð�"�Nn�����'�rv�y��-5n��XQ6Oʸ�x�WM��<Z����
�[ا�໾\�x���(d�3{=��k�k(�s��&�2�Ѥ��Q�!Lk����o����`(���C��KW��ޏ>.�Z��X���W(��~3��;�]f��ϲ�?�`���	ʚ���>������`�Z=xD�4YN�+UK���{S��=ie(���n֕}O��3�幑��5��|�:�2�����F�J=��g���a�(��~fU�I$ ��]��r|�e�t�()�o�d��e�|m���ú��s�m�rNi�����fR���WH��b�����Bf��(�Y��C�[�z�N�}~�%�.Rj��G��6A�RY�Ae�N��¥� .�S�M�什~�?pa��&�7�I�̥;ϻ�l��d���]��/vc�K'�3W��~7	CJO^8�[�ላ(%U�z-7�Z�Q���9^Ct�����Y�:�Js%���܌O�\��v�s����Åǩ�/V���Syq���d<�yN��[�_OfЪ�*s���vU������(�µ[��S��~E�!~�ɒt�����:^�2A�gbL\W�VZw}�������3������]
��7&`sO�Q"E��o	��Fh�yO�m��k ��D�J�����<�+��rK�����+���$3�M�Q��w۶l�K6 c�H,��+9gk�Q1��v�(�M4d�᯷�p�>'���P��Z�i;��&;7�.W�wc��b�C�$3C���|��	�v�(Cw��h������i�Z=�ɝ(��L�l4��T��h�]�+p�$W<z<�*$�:2�/P^~&/��
n�/Z�0<\��/��?˼1ͬ������ J�T)ɀMX���bʩaB�@�����H���hY�E�J	�
�EW�x�FJV��m�~8��h�=�1�J=*=u��R��p��\.N���._��[���IPS9G�{��O��h��q}�0P����V;U������{�5���� 8��6�� EA��X(J��� ҋt$��Rt����P�I*����W�% - ��I��s������ˋd��S�羟��vg����+Y�����F=��!^t�ߖ3��A��S3~�FFد65~,r�)�O��O	1Đ��q%+�U~���G��ǻ&i)��²,�+rX\�{���oTX�\~U~g�M�3�lM���r�At�{�7{��wDȄA���G��GђS~�S���]���mq;�]H9�A�8v	f9^I�1�WO^RZ�<�bs��\���\��?e���� ��:b�S�YB���wO�k�◉=�)0���n�K�Q��S��̉�J"��YI��C-S��6�Q��D��z'���Y�������,6*EN@m�g"����N�os�N1�]w��yY��օ��ܯ{1�a`YR��d!�]�R����	�~�V�ｇd-���_uLl��+1��A�x?P���E7�kװe������g����w�k]�A^���)˻a]�����h�fo�Ж}���&����h���W��-eT�rN��0+ߟ9^#��1r���vCo�B�]���T���&����:�f���K��ߨ�����K�~2G��>�"w\�~��㕡���ܨ���G�$�t�7?��g#%r/��+-G1j�=��f1��B7��E���#�Eϴv�&_ύ���XHm;�/T�čs_s>�1 MkTt�l�-��y�lta�\��\ ��q28�1Ja^��V���l��c-��1AoB��9�9��{���I ��.��q/�ιj3��Fol�|�)�y.B���P�է��.!p��xSc�ZĘ�¯�g0k�J�����n����[�Sw��<�Tk��f�W��y;"l#'���h �W���$�J��nƐb�S;��H��DSBɯ�_��C!J+˞�W��:�E����	���*r:���<k�༦&�w�y���Ǯ+�!�O�%�m��U��k4)�D�.�1
�b��3��ϵ�'}Zλ��I��c�&?�t%M���bD�3�2�}%{2��ʰjsi��y��S��eՊ�Q-�<����Q���a�X����>�O�]���..V��� �������m�A�9߅��,f�}Km\%ѵL��'�"���z1bw��ظ�둟n�uO��d�!	�7�[���۴3��������핪�ɫ�T�=�ZQ�G�kU�a�غ�ۃ�לB�J�l������:�M�JsH������<!��5$ka�<vc}�k}iBU��U���:��Q: �O��);%�k���a^ZŲ�'ri���}g��=M:�d|���~��	�G��q%���!�N�m���e�4ks}�LVRS��jֵ�F�x%zfﰖw�p��}�Ő8�!x�8z9�C���)��H���<,�N5_���}�U���Z�{f�1_��Y=��Kм�(�Ŝ�؏���"!��~_��9�`ۃ�;���z>�K�J�v���~�UFEԅ�Y+v��Z�e�X�;����4��$�/�ߝ��1���`{���E���Ыv��~���&Ԍ�4*m�?�pBz)����
M�*$�!���0����/-H�tۛߋ3j����ƞ�Zۦ�5���ݧa������?x߆��ٿ7"Y#�t�WZ �TFX��������;\f��mB�i��ά�}eg�}1�?�L�>��P{x��n7��M�#K:5f�qB��m����xr"� &8{g�L��i�e���{�u@0宁���jGƐD���֧'T��'ϴ�J�?�=�{9LJ�jԀ�a�T�> ��g�C�L�WN�;^ñ0��J���L��ĸU&�W�K�Q�ta�
)�Z�s�C��3[�G{�9�9#R�6lZ���~��s��ٵ��c��{�T���W9C8����ɛ��z���bo�(I$c h�,��YmS .�90�d����9>g��j�k�3�N�^�N������ʩ;���٣&m�F��t�G���j�6���'���n�U�G���q���'rșLǶ��"��O���;la�j�b��F4��An��Թ��p8�poq���e`����}�Op��*q#�?�6���wP6ZOJN�Yj`��L�V��H��6�����˞8v|y٬�>'��p��ed�i����f�P��Y0�:��¸⎠�3�����ϗ=����J:�
��a��w���eh�������aʲv)e�3Y�Nt�]y'�ʩK�\�rىB�tC=�4r:O_hUY�)�xJ(pE&Pj��8�U�z'b0��V �C����p��%��~@��l�Q�]1�o|u�1�?��j{>(�@�D����e������|��ayT����/z���U����zc�L�L����F]<�;X���xt��a������"3]y"|*-��%Cr����'p0�H��MkiP��%А���"���y���\ۊ���U�/�.��|=���5��J�CS��j���q�]�q�k>m��%i�<L~^�ȼ����/��L��w�'z4��r21@�lMV�w����#s�}����:R3�D���*�ڵ��ڱm��N�1�on��~��.Rv7��)�;�[<���r��D�	�+s%ش�_�&r2"��H j��d��\���^"y���Q�8�b���F�ԟ��[�y���˾=\8R(��AvM!MU
���K#�5��K���9YiE함�tf�}�K��,�F�@���O�Y
�R���T	�4�Ijs�	�u~�)<i[k�^\���P�������n�2���a���.
Q��V�Z�Yk^gč�M����C���N���p[]y7���}N�_���������b[-��\qK}��2Q����s�]���<����yW�[�es ��i7�GM��i��@�'��(O_�CN�n���K��T�Y<�����}��]Ŷ�<�=�&�R�"w�4�,�c��wN>9���40+��S��WY�m���٧V�5?�ޢ�0��.��₞+Gc��Y���V���*s[ɥӬ����X�&�^�1�J ,<}@�Y����П��&>�u^�5�G�zo�<�]8ϩV^�4���`^�aEP7������mR�����M��������[OM74�V�eq�q�w��3PI�[���l�~k�m��p��+v��͸�ɹS����������ͬ�A���@��n/?��=O��ݣ��A����K�����Xk�F��/�I�=V9���.���p/��y���7.�)Ё��u8�3��Jf`��������_����C$��1T�3/����0�\C� j��u�}���p�	>�w(�"}��&'f-��H�`�*�\�_�|�?񽁒�W�y�d��*&6��?�!��#�d��f��έ�h�Տ��\�����=�ִ��1��Y�X��C&F�U��&�>�/���x�	\z�o���U֑��u�'���O2��^�yo*�W�FP{<mz�n��͘2&Þ������������}�{y�?�{�n?�u����2���x�zU̿oV/��(�#W@������Z.���k�xPp���&ɸ�ԡ��`b`�~��Z\�f��G�9_�����ư³�R&�*��iκE�6��JY�D�\J/�-���o�)W�Ǉ�~㱳F(_�?S�8.qi�a���É/�K�=�6�x0����m=��}�|�T���(&<��N$8�/�"��{�!�7�BI�
��_m�h�N�s�0����J��ª��*$x#I��2��~�T��s������n������2�g�,�œ�I�C�b�TVK	�b���fL��A��/�s�Od"}A��A.W�9�)=l���_9@��P�8���^s��C~�sF)��ԽC���ϧKg��5��<=yɰ�����9E����[�%Uo�︜���Nt�?�v�<'�m����+J��웤!�|{ƌ+z=�\R�`�=�mʫy���}]�rȑ�����F� ����ض&��q��GXg�y���
���N�0p����t��9�X��E������'�9tx<P�}1*�7���S���]uٹ��4H�p�����]�N�Jr��Gm�D��&�J�bn|�@�c�ɾ=������Ơ3f���%�!f�E�%�i����xM ��z7�f�k������R-�
{��XP�*��dnO8Y�$B���}��?E0����f�"N���&�?���XX}�[3L���v.�k`�lND^�nL�B�V��-�:������u-Ruو�f �J,1ї�ced`�������{6�,ّ�%��P>�P�G���;�b׾���&�@#Ha���(�.L�xzۛg|"�fn3G��=���h��| ��V����%3E˹�I�$'a23��;�w���󂣖ɥri,��}�T�ln���J�[�BY׵�=�+�ϷD���y�в�5��G]Gy��X�ȱ�����w���E�vW����Զ�
??�����}@P��=��C�e���]&Et ���]��an�ݓ�Aq��:c.r"C���b��P��w�d��٢���.g�]�RV�+�
�{�黍g��6�8��7�j�D��-N�c�+��9��>q�2�:�ߝ�7A��Y�|7��s�^����˵�l�����IY�@�.� {��Kr�������`�{�+F��M�{�>��'}�+�Pàn`�f`�h�
(����77=��$���'\���*�D�����M�ۡ�u��G�H��(͌���r���LL�rHa��o�w�l�;ڦ����mj��v��^�k�	=��=&�b�IS��S��h��~�ș��J�?���mH�Wu�U��~���gp3h/�����a?6�Fk牳����{Z鈳i0 �����H�9����-�n�u���7��`���R4�ٍvQ4ٻԲ�Nw<!T�_o�P9Հk;���l0���۵<>�71�R��P�� [��BD���ͳ[-�u��7�)���Ώ6	�	�S�2�W��2��o~Uk�ho=V��?Fd�0ݥ�;_���� l�Wa�vzX!��\�����"�A��n�̤�:�-�s`��/'��'��\N��'pJX(����w�t�;�'X���M�,���*.�1=iUn~n�Z��?)X}a�|s+��i|}�1[,Ho	�
����-������"QR��Ak�W��a�s�{1�e+�)�p�g�mC�[C}Axt��$8K��V2p�Y�������a6���0��}�9�V��t)?#rl��ն�V����Qe�T� ��G� �_9͘�M��g�Wٶ$ήR��Е�LJ�Z&�l��	\���SW%���= p���~8߆�aaPس��4N̴��g�@���h$ȡ'w��8Ə.<;jwT�BK��|a[��H	׌dK��J|�c�ů�Ծ��+i��u����I��Z�e`H \_x�4|�k^���.>b�S��-����|��W�Ƒ��0���LÝ,�J��5C���u�\n��s�T����=��h4��Z�Y���Ч��}<쳪�ֶ7W0#����?�ڟz�b&�,���&�ڗ/_�
��<P:5�%��i�O��?�(��lK��ox
�/��t)S��@�U4mj���ާ�P`�8�Z����g���ÿ������+�^�Y�\ؘ7��Qf��"c��=���O����v���]a����N�~]���n�l^�Bk��Pdd
�#���qU�99��M�#.��̯�|�z��+�}���R���D��&^�Ŗ�9LU���L��X��5u��|� �����H�AW��"�ԩS�)Ĺ9�USl����_�i�P�iFGG'U� (k����gt�RR�J�EQ�mmmZ�V�\`�Z�lyg`�l����7��yF~��d������ΘĮ�������b]jj`����v�l�_o��]YU�gddt��_/>t\�����']`��Q���M�=�L��oD4_���p'W�} �W����m1^E�B?�����_�F6��c/�2�/KKg�U�<�[\��6��Hn�@��s�\r~})�w)ʯ�L�]���������ݵ��x�l��
�ui��)��K�o��T��^xD�M%���r��602/u���*@�� �[ifv>>>Q���L6}�c���}�h�N��R4>榩8sKG~5�9\ Bq�,�2���шZޚ+�!��f�5p��G�W��^��Z��e����]�=Z���oB�=����Q�S,�F�7-����G�.p����Iex�I�;,���@{"�NM�	�Ƈ�L�f������d�$vga�XwZ���i5����gCCC�ee�sz-��1f$&%��/�9�h:���(9ݏ���!ʤۮ �0��kdA���������T��,&RN���lf�+%��Б�2�����mu�[+P���b�_�>�e�f�{m�c�pb�J���Jt���[��/A��T�­+�=v�T2��o�`�\Y7�� �v��@�Sݏ�����,�[s��9}�a܎��>%��q��C-�kR���yӶ��X��J�Dm �<�	�e�����[Ri�ߣ�KyF5y~����E"�g�R%y�'�o�A��Y`���� �0���۲���������<+�Sݪ�uK��I(�KKA���l���*��ќ�2�� H��C��!'. �z}�S)����h�v6�5kWf�۳�g��� 5�
zB��7�O.҈�k��<��T�^�s����O]5#h��|���>4]'
�4	�iA���9 p���h�����q�'\��Û,����}��X�,ɡ:�,/��F��Gi��Zp��]Se"���Y�)]�ņ5���>w{��p��w$�D��ޜhn���G���`�f�f?%_���۰]1�����?�r˩?Vɛ���lW�;/��5X�A:�r�L��˨��Jk��|��ڍo�5�%�s̖2�R�n���'cM]��*�B��[�H�wzJ���͔@9,�>Q��ͨf�3�z�a��u��w%�I~W���Sc�6��~8h����� ��`�*/��t����=f ���c��M�~�}������x�����һQ�n<����[O�L�n�	�ǒ�?���vU�4g�b��K�)�\2��ތR�$3w����=>�D=��J�D���iM�-�iv7C�%�fU�e���v��?�.���-��������҅.�hw�s�:c@uE�E��RGGF<k^W�Ǹ�`�� //�B�5�!���۪��H���P��pS��gо���Q(�83�[E$/)+F'_ߍ��7n�஌�*����w~��� ��p���)B���j��R�+��k�.% L�<�Q),eN]�uD��-�kR�Vc8`h2�?r�.��&�0�9��D!EQ����t���5��"ŏ�Y����%�������M���;��	H؜�'l�P������l%n�	g�:$�=�Sd �kg���B�Tm<r*M D�y,�Y#����>ϥ���%�0��
�ݥg�Y�������sa2j�J��U.�@�ֹ�cz�s�S������m<z�T�ұ�3��u������-�E��h�Oc
�j��X?�1�|�.�� ��$v��ڙw��(	vHT/}��,6��Ʉ"}��-ݚ�ҪP�W���lF(�x\ڋ o�{��k�$��-��5uxX�{T��o}��L)�]A��Y���;G�G��(�Ӈ�w�?4�����͆w�^:m1j��������K-�Εԍjo��F�f���t@���F��?gW7^�E�s��D8(�=:U��[I�}���G"��#@�ν+n�CP���μ�z~�jW����ڭ��=S�s������gE]�6��q�����T�������쮈�Zl�qqI_��;�)�J�Վ�������2C� ����݉�����	�{���M*)�*y�M�[?�)��[��E@-�7wŨ��5�:�]���%�QC�V����ms��� e
e���Q�;~|c��O�y�9o:b�A7�'9�A@�6a��S *�ox4�<�'��mʾT;v����5܉��7��פ����ռ3695�5>>.���J"�o�n��qRq#{��V�q��*u�N��Z�XDH׬�u���+	x3�ت|�L~�`������/'U�EsH%�VW�����@/��I�J;8��~�Ў0x�-b| ��:Ǯ���	@�*ǔ��H�$n�j��{Fyi�3KjQY)��ȏ?n.s�D�Me��������ڝ-�i��%Ƚ�������Q�8
�IB�72x�+ng}5��:3���cW�-V�W����ȋ�yȴ/6%� �ِ?9�<��ߨhۻ�hX����6�|Z�R�2nW������0��i%D����O��L&��s���������.�Cp���WZ�О�2��h�ll�n|+��i��E�'�Y�Y5��\T^�m�zK���*��n�B����;�&���p�G�f�
��ᨆ�S�#�f]�M=�{��O��k��4�,^TTL��ai��*cr�ߕO�X�eɊ[�C*�n6"���l<v�a�v��c����~o�]��Լ
�zp�ޡ��~g,3C�����R=�7��
��k>Ԭ����Oi�h�F׬R��3y��_�n�Ta?�5f #��L	��Y��GCFF�
����	���F��bT�z�^�� 
�BJˡB�*紂�.�F\��UJ]�?�`��[���`��GO�
�\Qjj<��9�}e���f ��G�`�B���\}��l�\TTt<.'_0�jv�{Cv삙��a�Fnt����Z�;�i����U�B��\���VӅ�KQ	Pפb�.�a��gv���l��:���zi&�'��]��4�t��m�܁�\�
��{��;����\��sEQ(g����K��{�(!?��И}V ��0�Z;0s&�j5�������v{��+�@�{�W�䝕@�h���opD/��I�wft: ]7�kdǍ�W��-!�)�.�&�wĔ�G�ݜ� @���jݡ}Sl����ޛJ�S�6xr� 8B]u�P���������i`�ܩ_]9/��:�t(!j��9/Be�/�6g::�������5/�+b.]W�,��T�?pojLRf�Ϻ/${걺�$����=�ӡy�� ?A��e��z��W�ה��8!,d�]�A��,u�2R>yM���#��P���0HL��K�Ml��S���wܱѭ;��ԩ4x���f�-yH�r�3�n����+=m9w�x?@�JGgPP~���n蟥>w�-�+&yQ<��$����s�z�_�PfX�z2�N\�kg�1�WD��Eyq�T��!7Y��`��
��ܣ����
¯i5�<lJ�G|�UH��	�&*�n�(� j��ChK5�_�5]����VWB��Q�ą��/���o�[�A�����%ƩD!;3ڡ���E_�Wb�tn`�]��Ǐ�>�###�8;+�.Ι��������·[� �j��S�=!�U@���_�f������V+��8��j}Q;��T�cP��)י]�S�	+��,�@� 7&; *�
ei���9v�
���j꣔g�;���ęJ�H�R�\Ks�1�ąM`�Dhʽ)+� ��F&�;lƿ�|�o�
%ˎM�ߧ|���t����W��w���3�jˢ�g~F��<;�5����|�� :,^�7�~\���F�5��p�&���.{���f�3�a�-Qqs+
�H�d��5�j��
�>��`c��m�+o_�0	ʨ��ni�K/S�?sE ����:7UͺƳjj����y1)���V�,��Y��٨�RRR{�ϨE�{PAz�?�<��P���D�X�#�(��q��;QMI���v�� �X�ڂv��� -��j��w�-�җ?���K����rF�sY���_i��n�\�ڷ���u7�w?��I��[�~���t��1���݅�v�V;��P�?�_�ԹT����M&�(�E,�"y��w��E��U6�� 4�ȱk�{0k8Q����V#�����WεE�5Z��W3R��ڛ��_�^�
7n:u�/ �R>2"lj|k��쨤h���b� ؜QSb?�v5 ��>��;&����x�~A;ِ	�S�~4�}�C���@�sG;��э�PcGǝ���35�]-����ӻg��я��a�;��{����ƚ7�<� �#��m��fo��tDTTvEE�PHbé�����h�C�e��掑���;���2��ўZX�2�7����ٳ@�NL�q�6��rU5���c]x�~�2�'���l�b��镋ўk9�M<2-5�bMr��e���Jƛ�>������˒���y�J����9O�Y��ȞW`��!��Q����Z��_��;�ʁ4/�S5L����{�1mȷu�8��]�"�S


/���%����>��m?G��5�}o��Js�H�SƮ���:���?��ey��̦�.0~���I\�����ɩ�����78b����hk+����F"��*��cV���HRRa���?���%�� ���t��h���$�:��H�������Z$9wWJ/��\{�G�+j	v�d�� ���*g�غv鞿j��*�h����V�@�8Ea*ٳ�gu��?6�n�O�O�;::�f�e��w7��6b
�Y-��G���C��	��v����x��K�n��UU�vɯoN$����kG��~� A� �Ĕ1;[[�;��;�T��ʤn��'����ʺr�F�X׫:���x���tΟd�������.��~�{l��l�=��$�����ҿ]I�U���&�̉~��V�9���^������`R1uS\�����x����fff�Ǯ���L���"18y��4"��.M������%���ˁ����)f�X_�ߪ���9PZR���<?����[���YS�4
o���;;?���q�M�8�̧׋T�y$;8:�?;̫���P��h�ԥ5�F������|��w{?��������՚)9�\������Lܕ���EFR��/��z�鎂"v�H�����z{{��mm'��2.;ű�D?���TSS�a��ID�FNrh���0��_&�3�)�����9�[T��\~�~e�A�������ճ�6�<�X\�� ��������~��+++*�^�S����k����b���]����[���dx{{g����`�����/_ڧ��E��ʿ211�E���}�c������"��! m��;����&��I�Y\��ot\eP�����\Gg�+��x�G;x06�aø������Zz&_�&V�Ԩ���H�;��S�H������1���%�����]�Ȉ岴����h��c��ס�\���Y��㳓!�Ԩ1�����f�/jd��>��N pE�NqswX�O���.LMoz�|,v$�	m�A��"v ��YI�P薔�f֨��M��I�!�
���Y�m}�"'�$���������ynq���ak�Q�_���p��WLe�����hhh4�s�u�UL�NPH����O�P��ˠ6v���FS� �;������I
�K�`���x���mY�hSɃj7m��7o�\��R<��;���NO�`�LC��
����e _�D��S��h�-��Q�y�NIRA!�}��*RSS���j��aB|��3g�8��9!*?�1�C����F`��Й �9�:9P���|�PҠ���.�2�� z���O���p&�u	�o��k�������������
�-�@�ONN�Y����cgg�+b��5�u�1��\���������;��AR�	�A���ZZZ��`�F0>���5%9�Bw�a0�\�⨧בI��_������`��~� ���x�,�XzJ��";�\jw�P���!z��ӕ�(��"oaA�X�򢉟��'ii4��8=Y��f>{���&sy�%KG{����>د-�~��TQK8�2ޟ�VqE�.�m�&t�(�߳5����_U�$��` �%��Ɋ�8A�5t���S����z��������;0��a��f��pC��a��� ��l5�F�>�3/�� ��,A�D?��S�W� �����H8V��<��� ��CI�U�������YM	mO�'����ǐi������[��qq,�9�۟�Ė��e�(��k�7<����Q�,g���|�+Ն�����{����ERJJ�_d<���秅@S�r�T��1�2�&45��&4A^���i��qE|���#P"/_��*++��b___T�$7�`���6-��� ��(b�Q+�JK�, �c�F��cK���2����;r�K��F��B�_��'6_���� R����I�UU�����EA�ei�ȭ|4����Y�봋���tZr� P�M�<�&�r.l~&�"���)���&&�v�/��Y��3�
���_�x߿�1=�0!M	��������|�xh]�Ǳ�.�x�v�'qtO?mJ�-�|rH����9�RuQ��)�!�+PM=�����1���h�kl��4��uS� ��#�\\���q�c�y:�Yԡv9����B����e��`0��JO�|�Q�����+���k H��O�@�h5܄�+��Ç0�?��NHK���jS9Li��)�Oq��Y���w�q|a���p��R�{sNP�i����� �g|���:�CE�\Md�g��]���0{Q���V��)�s�da���vU���u'� �XF=?5%�����+�侥�A� ��MZ����
:k�=�i���!t���H�R

��5qo<� a|��4 &n�@$J��w�Ґ7莰ބ&����ؒ��� \�;���6�6����X���ل������ƺ���'$$X��j'�=�#k�_���*y0�cZ�ӧO�����D��uv�~q*�Y�-ѡ��$J��sss�-���;�yM�Q2�BM�FFF�>���q��b��u�-���n	xp;(�M榦�� ����~��3!���.>,�ԧNA��b��=��W�X��'< ȫ-����a�!�
�
�"���Է�xyy_��l���䢣���> � @귾�Zd_��/x�˩�j����vJJqN����mG���~b�X}��R{o��ϸHuk㧮���r��B&�i�����(�4:#���=ҺR������~'����3l��b1H l`�b��c�^��s�:Н¾���ﻎ��TF��^��Q����m͚r@�@����<��h�eē����.����*�~�aB@A��EM�4����p��*9ɀ���D�Sp�83�A�r�Y:v�lo\�s.�ڲ��7.���Z�V��IP�='�6!*�ӕ���M��*s@8�W%@��Y������\d)�5d=��jVu���ŋK+�����\�j�(B��^__�z�uĊ��|��['}B�����w:`���
��Q �\��L a_�-�*��]bR�ޤ�� ݀Y���QO04^�V�z����XZ�������K������P��O#�?��%4%�~�ɼ� \㯱NɣBw
��~��v����X���m����F��m���;�Φq����� ��K�ݤ���oV
.�z�-%�߯^�� �.J�ռ߮OVi�n5��j\��J�,���&�ӪDB���}�	�d�U;!~�3�x�E�#q�kk���� {�}��fT� Tt�N����g�DMZ�ݞW��ߋ��M�6�]��
�P���њ�[��6`��K�ѿEoU�QŔ�]�c(�b�iaT������{[EM��iS���^�����U0�ʗ�Z �`;�N?�����^��ɓ�j=�su� lTy�ed��靉p��ē���e���L�Nk�DW�ŷ�j&�Љ�3�)Obo���N%{�F|������I$��N�WC����-ܐ��)��^0�o���MP]�6�s�hR��4��-j �`��4���;FO�N�n�3����(�3��D���53�wjJ���۫*�AhAEɚK��-Pb���Ф��"�������!@DjHLLL\���~I*�(IK�@b �D���iy��^�]:���A�T~UUUN򷻥&;f��+D�u1����qj��/	������"ٳU�@�N�T�vV W���PB����<�;�Trg�����?�3/]���qF���o_�|9I�� Ǟ��@_6-iJ���Mk��;��L"�5��(Oh��m��\9;� �.@�hKx<�Uմ�V\��j����<t�P���\��Gy��#��}kft�+'�������
D-+v���uc�9(�s�,O߇���2����f=G���.0&
��� �����_gń�%�=��D�^�<CήM��t�h)Խ\����G��<H<��������"k0�#��T�޼݁�����x`�̼��E��#=Ӓ����k�Y�6 �@-��ń�j�T�	vw��8%ew�ƹ�dPO���N������K�Ɛ)�mN@�UH`x�����zx�^)���4G_��X1%Ya�	��ۜ��C�L�R�a.7��)�T�����P����u�D*,�|QUQQa��	um�X�?��C�n�z
���z-e����H��P����T��({�z�MW.<��}i�2@�3�-�3c�Ы �Z�"�}��y:/����#��ʊ
���t��мV����������ԫ�F�[�	>=m�R�7�����sL!z�{k`J)�T��p��X �R�����������;���`s�a�E�^�+�]䕽������L����1)g����I���k�j��Ih@'E.�ZZ�Z�+��x���1�.)]9�.���?�LRڨ�OP�HyG�+�w�~C��@ *Gh0��
d{2	�Y�HV���t�N��V�|�^A֪��K��G&����W�̀��|�v��{����44rY7�a(x߉q�~���O�)�?�T2I�����.{TH�S�x����[[�&��XGʯUg<��)b�� *şj�.*�4a?Z��/���ʙ*�������������m�
dP�����p��y>"2�!�ѱ��r�l i�~��y`HEU��6�������]�}��vJp8�������#��3� ZЦMD�&1�NY����d�~k�Q��t�v���U��k!�A��x���nB*rR��xd��
���s"��V��Տp�f�>����D�u�� ������J����67�}�U�e��)gbV�l��(�M/ٖ66g#��C� ��c���x���n���9���ꛌ�>�q��G�vvh/+I$c.����

�}�:C��0;� �n�	��?��m��SKM���y� �[W�׳ �zu&�PX��r���`N"�詩��..��zZဏ$i덅n���ɨx�(Z��x2E�s֚I^�h�&�I;#����ј�Ud/M����͍��)�E�^�F���K�GKS�r.`wKY���Q�z�h{��?ۛ�@&��줜Q�ܖ��D+¯���fg�
�}*SRZ� �"1M	<wK���~v�6�7u������џ}U���СL@_U�iv�/<���j�|Dp�-j<]�>s {(
6@e��)R(�

�*��@�����B���j�,0ߡ��H`y������)(�v\||�:|���R�� �R �6�=ڴ9�y�����'$X�]�j5�	���јN��2]��Ӫ�s*pp=���8
i��H z⛣�iK���?���hV������<8i*
���Ot��ݤ/�	�m��d�FT�7�|#�ٙ�@�`v��Y9�	Í=��oۻrѢ&O�h	\���tM]������NHS�42-9Y��ԅO��C��D"N�єf	K@ ��T��0l�����mq�ͥJ�t�A��	TolG+(���q�`��p�Q��=.	���&� ^.��vJi-��@�����u՜n�K���ъ���J���c��U��q������c���Rv���?��ݸd�M�\Ԣ��vŦ9�⊻�[d2.>��f�׮M��F�ܧ�n津���鎶��v	�s.�*(�*�oo|~Ɔ�	�5�-�U�I�z$M-�<)1 ��W)2VѴn]Yh��4��������u�pÿ�h���	����n��'�	E�)-��{i��m��<9�]�->ƭM�0�@]�򰵷?�Xw7��A�����wT^����A�L@��j�٢��y��6X���{Y�8;���2h9�����	P־>���;�w#T
�"�%遦��xW�S��x6�?�{w2�l�w4�V����H�=JBE����3��S$���S���כ�ii:r�4�*e�&bC��u�"v��U�Ϛ���]coӢ���q�ߝ�)c9p�+:\�?z�YC���z� J��e߼����|��0�v�3)�O�PO#����[Z&p��P�SR�kH��?L�h=�Z�ftr�"�������V��:m"���x<W�a���n�QO�ɹ"/��+)�
j�����PC�s�zfN����f��x&u)��<��	%vo)�������H<�
]��q���ǿq���&Q��l R)���������\��Y��K��)�A(A�}��Q�����ed����B��=��a�� �K�P�m���!j��=���#��_+C�!oB�����If�٠��6֐[UUU]W������T67��m����$��߄�E�qvIU�MO��0h��b�@͡/���:����w0	[�4����~Aql)u��\��_�
hh�H������P�9;kV�b2b�i�%I�m%K�([U1��쫮V����^8�hB�l3�E=��!0���K��A�4�����D!����c�T#���kk;D�Bm:�*g����Q�VI�<U`�ڔnӺ�d+;�aN.��Ɔi�~g���l�'�f�;U"��{�G�);3�i�������E5�.@Y�ZF�!����+>�Ua���\!�����.�t���n�:�#w�`�U[�T�5�J�
���y�0��
y����w���#n��׷�sS���(C��Wa�k
w,��x"Q0C$R������e}��a��t�U��a��0)���r3A=���p� ���������3%���ǽ��r �����
�Hs�f�����j���{V��F��&{}��1+pG�%���)j���i�f󈊛������hhf�'�î(���Kç��j͟�'����D|ᬋu���JjJp,�/Z2�#6�u|��u�>� ����3!B|�s�R���o
���:�4� �ՋG�-*�����ҩ�ɵM�P�Vx�E��=�ǖ5::��������tZGzד�_���f�ץ?\����KEc�3���>���t���~?�@]�gG�% {�ڄL(G�����ͩ�/S�>J��B�P?�(����g����>���*����H ��K5�eZH.TRCI<��?� es�6�T�h=x��O=-`���P�$;���"�ZGh& Vq>:krr�3����4�5%�`��漦�r����E����r%�gX_��Bo>�	�[����utosD ��=r�E�����8��l���O05M�UK�!���� )IH������@\}�Dгo���W�Sk�5DP��̅�&[�8�X������f?�< �x�~�ኴt��t� ��/g����:�䰣�s�O�$��h���BB�fP��� a��s���>�7����9��Ik�J���A�9��Ki0:gڞ� ��)�C�����u�c���/����`�w,ꯆ�އ��a���8|�.C��\{�ਛR|#�Ro�fNP�MZ�?��FYk\�:����p,�=�ʹx����|ؘ��qK�Ԉr�bŮ�(���'���u�o]b_����g�� �8�%�/r0Q+�p���i�����غY�?��\�L���a��������Y�{���o�kE�����.؈��rZ�!#�DV^^��0�$a�7�[���F�d�$ K�;$N:B�R�Vοn���PK   qyX�u�Q�"  &  /   images/bf545c77-008e-432a-b90b-35b3da31b275.png�zwXS۶/ҋ��RC�H�@���DJ� !�^BQ�I�*E��H�� E @�)
��}������{�{����oe�5�o�9�o�9֘I��(ə����(u�5Lp�-��HJ��d��r�]ȼ��|��(��kxY97���v�K?K���H���L��»:UP^PG�� s�{(��t p'%�������:���36�8#AN@e�"J� 	�PHw_y�����+�(���T�j X��=}` YqaG111�,H�A�Y�H�I���K��KK��KHˋK�<���|���M4��9�I	����%/*(()���"*�D�$D%$�qa� ?(J�×�/0_G����p�u���S�T�w�O��2��L��ET\DL�/(�o�W-�ű�_#QP�:9�����q��%'GQ�;	����a���z�z�y��z�7��n�wK���g[�ȿѾ~�~�3��5��z��8�4pfrWdɫ{"�|`��8����
�����Q���C�A���H�	1���)������W23���+���(�����?�����&�j�����K^���i�N^+b���	IyiYyi��br�bb���{:����K����ؿ@q�8A���G�������s����D�<\���'G���n`���먫�x:��qZ0�C����+���u<|���0% N"�;�KJ�88�ʈ��de���` a&#,�9�9��KJ���_����*�������7�4u�_�J.h҆��y���tMa�޹���<��Q��9��������+�����|=���>05���8��& !)"�ׇ:�=�$ust�z��p�U(�sG�?=�w�E�-a�%�e�?�%`���)�S�KЃk����8>�h�AP9����>��u���e�@��Rf�v���qe�N��iƎ�7y[$W�>�p������It��F���MX��\!ȧ��7B=��#%p,�c�Fs����'
1���~f���NZ&��H�s�� �	u0O���R��`���	L�پ3�Y��z���o@��tr&31�m�Ĺ�oAX�V�0(TμtL?6)����oM0)����F����G�1�M�g�0ؚ�گ/��,2���؎*���<tQ�܈�vC3�]_ָ��Wn<ٙVJ�ҥ������a||�}_]��SV�Y
�	ܥ���ʿ- @�{"r�~3�N��,��m��m%ry,�|:��V��))G��w|���e#,��xM�ᯠ�בu�T�8K��-!'ߢ>g�
��A	ԡg��b�0��l�.ވ�"���:�8�m('���x{����qQ�~��j;��2�!no��CU�O�	<m�~�)\�U���ƾ�w��C�� �F���B.��ڽ5.��߼{]p|��W���m�`�H�������;jfv��4�[�������T�$g(��OX^�4QG'��LK�bP�
�g�Q�s�
����B�][�~{LEv��W���t�y�V,�)�8��1M]��PM7�y������+#�ݴƙn��=�&['1��-r����C�G��ޫq��ö������c�g�aq8�k�}��
���F%�`{ycF�8D�ԧ	FR�����-�3]ي9�ׇ���W��j2�컑�ґ�����u���&&F�-:M��N����wB"'�w}Osp*(���$K����?F���<�c&NӢj���n%@��w�b��ڎ�Rj`y�L����Z<�L4��,���֐��Ţmy�V?
N܀�&Q�����Xqj��+�:�r+��`A0.@��1�w�"��)���X��7	�v<f���S�h��i�V��J=}�����d�uin8}�掳��췹+ݨ�!^�N��4�����Y��&E}I��˸Rr��wӣt��1�����72�����ҡ,����_)H�$V܌Npɧ�'�tw�a}C�:>`_��j�?0���(�#�bzr!�X��F�P��bD�|�ݣ��MT�r�Oњ������ߴ�k�o"]!��A�tE�ʱ���~��i�8|g5ܑ�D$ �trZ'؂=����3��O�����2��-vn�r���^׿ҳ����	������B�R�!y��o)P=TQ�c����*M��N�<k��EMDT���}��~S�( �Kms��j�2����8��F,�G,V���j�Хld���H1�+d���`8o��������:�)K
�a^[�XT۶uO��D��1�v����*��7��Fg�{��k��"Z�4��
p{�D^6�t>;U���3������r�%r�UU)s���J[YY]���
�&�\��T?gY� p>������64ܶxs��p̰�)��V�L#�=gzbb"*g.@k*�uq!�]��B� �k��ZKwD.V��A�ì�CzY�sVi�l�8ã��4<L�w?,E�Z|�����z��4��.1G$Ǒ{Ě�M��b����B�I��4��?n�5�+���(v����al��I�^�����4�Hr\~��.9���3�#]���/.r���^i����5d�/r{Tbd�� C�n����KǍ�U��9kC�z��Ç�^}
�l'���I�[��q�ڂ��^0?1I����hͿ�,��	�m�6-�����w��W{�R���1C�dtO틥��UUO>���.�|�'XP��5�}�&?AA�FB11����%+[�tla�������S?MZs�}���R����-�i��$S����4ת��P (����-�c�A}�\�Y��ݷ;�CZZZ��\I�!�詼#��%����=;吝�%��Y��S�l�SVèF��e�>������u��ZJ�$g�;��Ԍ�<��X�ԷDv�yWd����(&�9���i����}8�!|�̦p��Y���r�A(��:��d0� ����"��Rq+u\W*��=NE6A����|��X�sm����r���M%3�yx5�h�u���������vYn����T<���|�(�kb�7P?�`}�C�ϳ���®��_|��ќ��Ei���R.C��CY+tܐ����V�+Vֶ���/<�9��T��񽙏�E��˳XlD� ^S�F�~6ӽ&�d֛����z��u�>C��a;�ikR��� ^q�CNF0�L���V���/��-PF [ ����9N�G��M_)� ׾h���A����[*���u��f�I����s��{��^�J�vU��U���Ѫ3g�`y�b�#`f��a����P�Q������.���HH,ԅX෼�|�u�\�Is+��؞�E����4��\��]A��r9z:7 OW�Tz��Vx��Y5�ύ�f�.����P�b���1���P��M��qZ[�\����5�gkEZ���[�A4L�������h$���$�IA"��;��B7�Z���<��������ý`�F8[�����֡*��>��l"n*�T4�3��\�(V��L��ԇG�~�/9���T��{�a,e��,��<7r�s�ҟ��5PGj`$g��3\=#y�6B����C�(����x��Ҭ���X���*P.����#n( ��M\�zL������L���qcZ,3����7B����f�ucXd��)���
��S@�}�*1/���'�<"�W��08]��B�4>~i0I��*�h�Z�ҧ�+wcΖb$��j7I��.���p&ବ]�`��w��и{�@G9�[����Ac
ڌ�BdҐ��17����mk�+�I|�iB��	��ڰ��K�[�)覘x
��]U���^0r�ׂ"j�)A�����E��^�|b����e�8�wf���UL<��VR��Z*�[mCS�������{%��9�Hqڇ�D�es�l�e�WD�[ʘ�6i%��.�"�B[h}i+�u�P~��/��(:d��������ϞZ�7�}[c��>f�΍��6�!"z��y��+��u��9���V�p��;�����y����\	����מ!`����B;����_���Qi�t#y$���I�rަ�4%�kt���:���')6���h�a��*ǽ�>i�������j��:od��*�q�D���
@XM>&v��0�!�)��%��׾�wAޮ�̎���**����hkB�Ѧ)�x��/9e..�,D����~"3;<�d�O������F?W�8�����'T�(t0L3��[~Ov2*JMIӸ�̈́�>cy��bj�Iy**�`�Us[Y�|��ME��Ô_��B�<
���c��7XB�㊨x��$n��Z�㖧Hv��",ܻ��˿��0�#f����l�k��(L�Y�W�ѫ��cޮ���\�q����T��VONŭ�6�T*������w�֭}Y���:98
=�!~h�I �� }9v�)�����̩��c3Fހ���߳�'��h��b���9�y���Y�V	+0eO�!�y�»����l�<氌����f��>VJB�-��A�V`�h.s�r�f�|{�u��r4[�+�#�şͣ���zVI8�6?��� �U�[����uj������G,R�'�vp0ܷ"s<_����W�͜��B�;#�a�aw��k2Ebg�ƻ/$�����{]�<|��c����|a�N`"�\�]��O�\�2#�o��/²���$�����x�30�#lB\kw�W�O�LG�~�I?��g>��k���7����jM�ȩ���Q_�.d�r�x��������5=�vY�%�����]�Qשd3N]0c���` �s��C2����/U� F�)��]Tf�~��b4���ȱ����pȒ���_�;c4��xB��sB�oL�Z��*o�C��I�.3g��2�e���"�{�9/�� V��&:�M$3�[���"�G�+����Q�n^��Lk��uܞ�:~���h˯��J�d�יɉ���[g��ׇ8�mT�%�I�hE������|�N�J8�#�Scc/��'��M�Q�=���n����އ�oo�r��#��ϲBO?D���+/�\J�]k�U�7ڔ|ů^H�v��.�W*�H�NY��T�t�һqN�VO+�Gi.nk�Է��V����si�44,]�[߀[oI�y�i���qF��
�%��y.��>��I��̃�2�d��Qt�+tX�7d�7��5=\2��q�;�[�[����m�ǒ�˵�PIV:��YWz����C6�\�f�������U�E\�苋���-�l�Nl�T^�'��ƗD�����#�H���J���,I{���7 ���g����]�rŗE�7���O�;��JKK+8��<ѡq��Z������^6�!m:QKT|�m����s������I5��6Sa)a �R����� �xI��q��8
y� j1���F�.U*�f���\�1��%Fޤ+kk���I!�O��7Q.�����D�Q\�����z��J�2���]9t�3�,mHN�:r�ź!t��'�� 	l��)�RN?Q�׍�s����WS������y�OϾ?�T��)N�S1�M��>;�
�dW�y���C��^���ާ��ΐРWj$�5,�'�2��[(/u��)02� �Il'-�!�j� �7�w!۝�h�۷;���O/Q4���v�"��]U�ƍ��j:N´��6dӶ]�F�F�51t�\�jM�4�����G�3�6(���pB���lf�����U>whӽ\�B����+ܗX��j�3cg� ������֍�)%�K�D�3�Do,��ҋ�x�	��d�I�x���b��|�+�����V~������Ri�j}���Y#B+�,s�9JPH=]㝊����2Y����_'/�Z�HBIH;a�Fj1�Y��T9���'�{����#w��E%޴g<d�� ��w56ʾ�����2�&�<?�ɜ��64���?��~��z<0���}DMfތ?s,L��$�#���;�5Ǿ�W�&6��#M�%Ƙ	Z'�Įn��z����F��BL�����|��$ �\�t��Y9�! \r��� �Wٶޔ����R���!���`��5ns��"��:/���3�O�CE��5q��T�Ѝ�
���T�3��*~��K8Y���	]>��7���X\�l���=غ�3�6`���X8��$.nI��ۤ+7Ӵ��j��Ȳ2��#fD�z��&�����:��ɗM�tK����<��}'/�zq�Q'��_>��_�W��}ͤ�����AP�F���=<����]Fȉ�����T#�#K>�ҥ�W�^���}`�(�1�HK��u��_�*&��O��x5���N3�8l��h�a��FK5���֓��;g��I���MY���B-�䨐�����&�@<x/v
zǑ��C�Pu�z�:�϶�'[#E�n�D?t�W�n���é�"E	�c�0�ց۫t&�k�o3�)L��8�]��z��#|��ߌ��\�3�`C���v���%��E���G�/��ށF�g?'*l_/���z=�"�L���[�S��_�]M�O5xj���W�4'L�\
�|'YՐ2ۂ���Rl'^���{p�6�8z�At2jb��h�|N��+((�2�ۺvQS�デ=�Ͼ7��tŔ�yW��q��%�sk[�Bf-�>Q�=&qif�u�=�����U��:A���]d���m(�RD{��z��g6�9��R]QyWϬQ�U)��p��pÂj3)�d�W�8�}r��N��Ni���(��oM����� K}�M��Y���a$����P}���0q*��� ��|��A���R��=�d�'�������Eo��F�fSe����̹	-�����ɍ̲l�n�RT<2���E��2io�x�6/��?q�f{*}�bU>bD� ������� �G��K�)��6�S�֩�����Ln��z��
M��s��^�&d)]}�L 9�u��S�T
?���ӳ�|.ݳh��$�tr����Ȥ�?�گ��E�=��˝���S|����Ɇ82X%�TƳhlG����	�;�}$N${�ӧP^P��&� 9��c-贠����3Ao����e�g���PEƼP�I�i`Da�����:���a_q1H������xS0���E
	w]�~�O�8��Vu��h�?�i�)���H����_��ԭ�C�+}��H�Ѿ�DXd�`�>��&*�_a��ި[_�؛��iO-ڤ4no�o9����u��f���-�Ǣ[.2O�"3�iA2�򛙯�γ:�)P�4���G�YB�#�8<���?�	��.�n�E�%�i��Xۮ��ҷZ&���v?b�~uI����90���eb�ԛ�ٖ�Ơ�)���t�{�̽�64��w�O�[Af7� ����>&p�8���ڿ<]� ���X���;Y�E�U�'�}F�>��2c�>m+�a��닅�ݡ����1�h�n�w�U�"6~�@�00"d��Df/��p!���V�z�b��x�}C��Bzg���\8�G��ϰ��%�){]*�p�@�4X*��C�˾�t&�?W-�E��Λ�N�OXh9�~8�;{h~�����Y4/��Aa���w��B���9��o{E�H�XЦ��m~��=؆�PjuI�.���u��{RSn����~j}�iAh��u��?c�ēõ������E},���h�Kjfn�g�mKDqO���I��kA�K(wNL�Z	-�R�^��
6���G/a��HG�������ٍ�/E/�^��[3��N�Xb �ڼ�g�tqR�y+���>���X���E�#���1����ӞD�J,x�s�����(S�U�{Hp�����:����M]�E2�����e�[
s׉�F�آ�/����wb��nNW*��u�$Hh�S;O2���dp�����ರ�뤃�����~+�w�����r��FRI�a�8�)��Pr�����[�}k'�3������U�?NX2�Xï�v��'��H{V�VV�Vz>��J�]鶵S��T�zWQ/�&u��I��&]4�xe�rT�53�.�Mh0�� �o*�}�|���d̬0��]h�p`���վ�ܻR!DRU����!b�F�������I[|��D���e�����h��Tч�`q�*�^hP�1T�|�S��H<ق��$u��Zj�l�+����f�ɶX>�Ņ&�~۞청��ZM������ڠ}[���Y%v��_��o/lx�8v;�{Q��cKQi]fA��Y;�IE�ֲL�������j���!�����U���55Ɇ&r4�?�u����L�ro�!H�V����~�G�ʴ����ajjM���C���Y���ީ�K���ׄaaa�$6�k�x�q���R��S_��L=�w��������ӵS�|.��W�ɉI�"[�@l�'|=�VԦ�q��Y�?X�(����Ti���ÃDM�Ɨ�?h��q톸��������C�T:���*�K��Ξ)�?����ښ�|�"�>��el�}rt��Gn�� tQ�eU&e?ol=�2�{sdn���8?���8�^����/QA��W��L{?n���D...?��to����}�/kF�UWW�l��
D�)�%iUn��o�/\.�˭�f)���%!���)� ���۞%������vHa�E_a���3��Y]�|��KM5+��p�r4SZ�Ǝz��r�	�6��Ӱ���,��){5g�r�	��0��w�ј��?�.�M�ύ�Y�1��NҎ�Y�~S�9Ufj���]�gKG�@��>�? PK   t~�Xp>r�  �  /   images/c13bb491-011f-4ad1-adfa-58d33d2d83a5.png��PNG

   IHDR   d   1   ,�   	pHYs  .#  .#x�?v  �IDATx��|{�dWy��޾�~NO�L�L���<w�v���$#a�mDJC�P1��!N��ʉ���RvL���*Ɗ�`L��Y���Xi%����~?�{���}���힝׮fK�5)��ݾs�=���}�;�������O\��ͦ�o��&X�z]�д,��ʊ\|�WW�ihȍ���f?�y�Ѵ�a�t�6wձ��Ӥ7���}��5F��֩�ٕ�e�k5���0�4�U��|��;���|��ݨ5Lk�g�����\7�k�wBZ�K^����60eT�@���àۅ���fs{�R����é9�o���-�	o0�b>_ �j�, աNT�E�X�����V�����b�PD����h4갚M�<^�s[h^���c�~�jQ��՛�6���C�4Jyд�HLr��N�vw �÷���Z<_~���YM�K�	���)�v;͡��GWu��A�,��'hhfGnkT݁�_{���{�é�/D_�$6�f�r�X��O.\����+��!Ē��AAHoȏr�!T)��r:F�"�ȗ�Dm%Oɵ��W�3Ff����H�͢G~+�$n7<��=r��Yt%�omA����AdWV::������(
0�Qd����P�5��9?���1LNNbhh�TJ)caac��p�d�\>/�m����33�������A�]�ő��ҙg0v�8�����٩֞�d0 k`_c��X\ZB(�a�����ѣ8/s���*Bd��[����~�a�5�r��w-Lk�jqY���y8�=������}�r�C&�����I��N��jRM^״�M>�ԍg����(?X�	��X��	�¢�auy�,�а$u�#'�D�Úb���&t,כ�K]�\�f]�o���!%�7�-ܲd���O`�T=d*1�t8��A�yz�aS7Zo�{xO`I�wI����J���M �ǲ�w�u�	�(Ε�+�G0q��:a\�b��=�����cM~u�.�Wם�����(=-�(=,ck���H(�Ǣ�!����%Otw�+�S�)WED�X���E��R��S_�oL��	�h�Q#W����Hw�쒱���_"@�Zǲ�@Ƕ����Ւ�D:G��p,����#A@�4
Eda!��"��k��qJ̮򙴙�6��g!�+�:|��e�_�Z�)�隅��7��H�\�HG���.����~/���MIT�5�㽘ns�dG�"���
Uge�>�`9�����;�_NB("�]��$�/ͣ�;�� ��ea�Ӊn:`t��?�+�a#� �y��:���T������.�`w}8���� L]*��BT��^GY�n�(�J"�I&̺L�lH�ti�/�Pgy\�w�B�A/2�\���܆R��+��h*u�CC!>]*#�b]�u� �&J1�>+�?&<���%�9�]$�.D�C�n*=��Um¥GEĮ)��ǿ4Bd�Sɬ�X���"���ґRr� �VQ5Bm^4u�b�Ʌ<La�卢m�5�\zt%�A�[K)+����ҥ�B�k�糪, ݬ�QS�g䠔P5������S�H��Z�"�oʪ�69��]�r
�F`r�T�"\��#��(
���� 6"�ź��Y!�\���cT���-"*�O�HwXʐ�!T�9��B,�H6�b<7/�r���]��˹$���ɪ'�ůu�����k��R��w!�K�VW@b�ȑ7� 7ʈvxQ�6�zj�+��b�}[ܽ������BiM�%Y<�m	�P��v�ŏ{�eۨ�~�]�������7�C^�#�Mnl)b��.�����<r�q^>��f�,ȭ+1U��wMY#/�N�|.C"�%��-���K����1d������0ot��#9���=E4�\���LY��7�Z5[�SS�Bqz��l9P�Gm���s��(����^Dؔ.��P��G��"�2�gfWq~=�L���;-6�u�5ҏ�>��Q�k"��D�h"�SĒ��K��|#����dr��b�H4�%ѭ�K���(b"�'��-!N/�����|�{�_,X��"�\.;D��h��p�T�A���qE��tZ &|{�Ĵ�3�6����H�IM��fڢÒ�'E�5ſ��_��\��	c0��B��>(��/��U+-?����D��Y*"Iٖ�E��pA�����*Wip��Ҏ�2Y()C�����R9�m�p���"�0��*"+�J�J=����l�Cd����]���b�|QL@q�j&����+�p��f:���,E�,�b��17��/އ����΢�t(1�]�ؽK��hÃ��N�ΐP�[�5Zh$���j'կ�J�>���t�R�`�7�i�?ԫ�֒��h�i�z���l)u:}��ᑖ�k5��ۧ���C�ug��KMkY���Y�W�R�"?���U<1�Al�L�80s�
�h�Z"uGD��NQȤn�{�/��b�~"�H��|��e[�+���
�!ѣA�\���D��.ie]�¥P��8���Q�RH2���;i��)�V�{{n�������"\�.��B�N���C��bn-�����('b��|�4�+\�oD�}�!�~���2��v�R��!T�y��N_X���FS�Qr��2DDquC*�$����p�ًaKqP�P��2��UAC�ԪR��Q��]>����Fw+e���0�CN�3���];�p�Dφ\���؀\�����0K���$�?��$R�m���Y��h����ex�������w�Ƹ�>���Fb��E&�.0`}�Q���{����������|E(�D�X�Xҡ��Ԅr���sgyI�w�E��gr���ƺnᶁN���1�:�8���Ȥ���8���yg5W@SD�߸Z�փ�P&�Y����$��iM��'�)�ծ�!C������m��CMGQ����:)�˵ֺ{�%�-��s���xj&g;}�(D-���'���.�wee�1��ư�ɪP��Ӌ�5	�Y�B'�P�ni�T���4�e���q̊����&>���_�G��uEB��o�#:V���cZ�coC9�#�!�,��3�Ю�ZADR4��ٲ=W��i���7{GGF�$�/-��4�J��L�yPG�笋�,�v!��!��V j\�p�GS�9:tY�+*��̨�-�t|��wQ�����ĕ"1�:��)
�n/����0��_����=Jw��k�wcp�%
ZEz9W"�q�h0���~�ד8���tFE�a��b����8[�G^(9��{h���ͤe��H��Nn�"f��fE������;fz��=A��r����ZΥ��ٻ]d\W�o!��@"1��X{��Xz���_?�B�TU���ۏ���B�CH	
c���jc�����s&�EMĘ������;;x���um���\Q&j�x�j]��5Ok��ɺ�P������T���&y���{@D�p�6�vw�60��Gw�妎'��P�+xO����ps�I�D�q!���@�܏�?}�P����ٛ�c�&U�ײ-0!�r͂��|fWLr��"i�Kٱ�.J�p����c�i-5���%�uu$�5T�oˠ��H����Z���y�a����
��K���r"��f/��	ȶ"����_�"����R��-T�4������J����/a��3�'��s�����sO鲥�����Ṅ��=�n^e����B"H�D�AK�&z���^UO����"?=�Ӊ��2J�+h��=�D$��H�����u��{�@7ַ�j��g!%o�3�j�f+(�"0];2-�.����8�_��_�ן@����)��!���٭�%�^�ήؖ��3�!�b
c	?�s艉�0��3��(�D=N:j8�яb����cڏ�~*��'��t ��`��h�o�nLtca3�D��,B����I6`uD�ٰPsy�����Eyg�TCI��)qdoL����&F�!��+�w��l��ld���GQU��~�u�\8�l�w�s�i�t�|f5�G^\���k�����3p�8�?�t�h���V��� ���T9
�$d�+G=dk;y���k��فB��V�3j���johT�-k�R�P۸V˄"u��K���?8��ׯ��V�t�զ=�J�ڈ�\N1{˰�G{�Ss+����x%@�{ؘ��RP5���QR��f�f�g5�E�x�62�\ �r��������N!�3R*�j{�~%V�U�zl���w�������%��'��3��Af�t6�̨|�JD�K�q�C���yԅ�F�r=�v��2_�b��k�xS�0HX��Ⰵ����c����RNcL���x�ٗ񫷾�x��s�G����-�".�9��A����<4ػ�*����"\���Ԣ�lq׸l7�ہ�߇�D{=���C��^�TɁ�BH]fq{��w��W�XJ:���k%����5뚋-4�8L!�:�~�����x�,��I�����p|H���_�����b���݉}�[
O�.�t�T�,��WIps�J�!��x=�B�ob[��j���1����&��f/�-�Ft3&�!�nx�`�fY&4��u���ģ,�9~J=�v�f��'^��>p7�ϹY|�k����|����8��;nƽ_~�r�8�K����p�/�ŲP/s�j"��N��%#\��D����xV�8n10�]�!�{�px�������e�n��-��>��m;D�̕-��ב�_{��B�ܩ��_��������o��ď��z�Gg��g2C�p#�]z�B��i�NzA�S��R��D���r��$U�v@���]Iؼ]�W/V��;�콰��b�rx!�_͛��fْ	'���,�������?����?~��ދ�gV�Ȣ���K_���v<��ϫ���~�x�sxaa����#	�[M�	̹�Wn4�)����Na9�)�[-�R�PW��S�s����ѦL�V)R�Y���Ĳ�ƀ��;l��j>4s�̟na���ȓ/�)A���.��K�
1g���R��G;����_S��4-.&Q��>h�������ž��>��*�O")������Q4}����%WV+��6BFGG���>���U�R�v�p�L�z���Tc� �ɪ�+��`23�#`|���M�w�x<�+�P�=�kT�T��)S=��F�SO�,H8=��R|�@���Q���9(�n�޹E��xw�2}��B��c���B��$�����zJ�8Pdu���`%w�Z�1����@�eǌ��ۨ4�D�k�����wu�pa
���na��
�=:N����yL�����{'�VR!)��N`�[@��%=�ɍ���=�Y��'�vּ$�䍩�dm{ϝ
����P����f�w��XIe��q1�W:y��G�����6��M��tv]v��Xˉ�<��J,ߘ���>��8.>
�|��_=�WX�D��~'�ٯ~�H�|���xdjf��>Ni��:LQ^w[�Xv۽�gD�������'�l �^�}��JK��6s�9ж׏�8���,E{�5r'���~���uյ&�guwv�:�p\\<��c�j`u�E<�O��N���6�ʶL�����-<����S}�puA�?�'����W�X�=DH۟Tl�j�۩ ��]��@�L�ǽ�\�������m��I}�q�cv�U��C�N2{P��$N�N����;�<U��4p����[7���(�Q]C����alb�Z}�}l�F���au@��	�D���S�[h�Evg��X�k;^�^h���V���g�-��l�5���<o��3�e�>b�,vZE������C��+����7���9s�i봕�%
��B8UG".��P���JU��fg͖x!P��*Ң���ZU��#��"��Ib�����e�E�im ���X�u�p9�9z��c"��
��ф�:cC�D�`GH�!x��f$��iJ�ch��b��m)hM��Ʒ~�[>4+>�3s+eC���}j�-��$��u����Xm���1������ut��^�BY����7~7�����{���+����9@��9Ãe#�O��?��֖pPC(Ɖ�x^Cѷ�7�;�%\��i�l��:�H�sH���::@��0�G���Pg1��b���BŚB<�M ���c����`��˧_PQ\"�ͥ�9����_�
8�o�)�k��?�Q?��3�U�\2�4�,�x�u�����s�>t�B�erPv"���:yD��{Q��DlY.��ݨ4�0B�B��ya��0�=xy�������BIwb��B.G��h�x�R���G�\Q�W���nLt�{���Xr���S���ʨ��J�0��y�I)~��� 
b��Eɦq�/���g�j��2���Y�C����s�!ļ��,ƺT�J8�}.r�UǓR.r.$"k��;X�xW3�
w?�<��������8�=��Zωǿ!��K���Mv����� kn�d���g��Z&L�����$4� �?�a�6�ؠ��,S#/�V��z����Xb���i��>��#X�[E�j���E���\�����1��Ry��|��re|~�k���L=�`�k� �{Q�)v�2�a�X8�tY�/���@P�s��5�)8�K.>��yq���fϟ���)�(�|���3�#��x��C~+� *�]9{�,z{{7�B�V0,z��#��5ܘD����׿��:1�(�n�XvY�-eZ65���7E��=�Μ�	⚁�|C>~���~Y���$�g�U�~lȽ?:�B0o9׫g�&�v�n� �����
�צ4$H��v_�i��H0�؄Lq}�!Y{�F����9�N7e:V�ί;�wM��*�y}2Nv����d�E�땺��R�����`#z?����
�-?=��d�x�r�umy�_]} ��'7;�����o�F�[��Kr������l#�`0�B����pH9K5��z��133���qL�o\X��)�1��߯"	bũo����9gRI�~��ȅ{୉�|����p��������a�$򻾾����H���e�����o���j��K����4"wߏtt .���a��2����oJ�7�g~[���)�_G�Mw!;J�~E���Z��wO��$a�O�8�t�9r2�jY���K�o�5"ױ7~�N(��1w��v��0��h\��@�1��C �DL�����[�E��:�N�(u=�a1��� ���f�e����(�&n��*��qՎ���G�J����N4�.�W&2���8Rސꓙ�������/q����R/sxk'J�n�$�1Gd������/ɵ.�{��F1���*�\��%�����u�\"����lQG��	�:�0�ힵ���j����rw����i���s��#�8��wn�~�Ĵv��m�s�:M��םb���M�o�8J����n�p�Q���:j�i�*�    IEND�B`�PK   ��xX�Rr5�  5 /   images/c34e957b-2bab-4628-9db9-846c7013e8bf.png�gXSY�6@���c!��cE&�;l���ҕ�*EzO�(�t,�����
J�*5Ajh	5��Cq�yH��~|��o�./=g��ֺ�{����g�_����)�	����9}Bc��`�>q������ ��f��W]`0�S�o���a�=�3'�/yƎ�pe�00ٿ�ڴ��E�=��͏;����1SV6�[��`���9��w~�K�*�%�6׈�Ǚ#Q#�˿�Mi~?���u�Y}��!�+�~"|P���%�1[�ߊ{��}�z�|�/�?�X�~W�@z�3f����jC�?m����q�9���?h�lĻ�;x{/��YBS�"f�uF����C�<���p_�y'7|ÝWj��x���3M��#t�R��s����W&�j�0�pKb`��/{\y�T������;�g^u/��*Z�~��n��M��JH �h{�;*"�t9d
9\�fMϚ�ċ��#��.�]'o�&&E�F���MܓꝨ������8�➣�ϟ��X�g>�1��W"b�������9��p��ut"���xx�+w���ȳ��!S�|��r,�����ʫ��Fp&���B���R���!F�$�}��K���!��N�����ӷ�U�$^f*�=;�	��n�X�w��r�ܟ�@ԅ�kW��O�ީA9���D'ԋ/����W�}�H]���ǉ�3�P"n���t��j8��ܕ�l���eȔ�ћ����=��L�6b�E�h%9���Þ��3w{������1�I-�v��,?�+&Fp�g��؊z
?|��AT���{v���!�*%����زkAf��ΛsK�f��*���-��O=�BRO���'�^�Iy�y��_�1K�/�6����`nkk��1�	���Έ�8��8		��U$�1�hk��v6�M���9׆�<TI�歈4���ѹnNZRQQ�v��V�k}�T�ӥ����،����y��+��:B�JO4�4d
]\PX~m��v���ޗ�W<2w��@ʯ��E�3tJ]b��3 <BnDv�L���QVA�*?��mV��oߜ�ܤ��7iL֗��bV�������O>�A� ����ۋg�����C(�����[�I-���
�a��=[��������=FVfO������l�R�e�F����2�^l|��W��\ �N��KOx+��M|�������C�Z��n�G�������-9�C`>�:ឰ[��q�a #;�233���C�s+��0���?��M�^�VV�ec�>��
)��sޥBR��.���8�Ԥ;�����魶y�9hu����<���=)�r}�ֆL��J���M�ܹ���3�����|)����3!�1�Qi&3#cpk���C�,B��`��!Khǫ�W��\�|�}=D'D���~�i���R2�H�r��"�Qc��D ��W)Y��O	�8O��$�8Drqq:C`P>싄T��c� �H���C���J�֬��zhxh�9����Ǥ��J�$Y���t��"|�]}���A����XoI�� QG*m�^'f�;�e��/V��2��у���
^(+I�|ǿ[*�\�	�)�<l"�����x%�*���,���Xߊ^�(����}�L�'o"�M�n��[1!U�����n��*>�eQ�U�o�-C�e�K�t5:Ӵ�3R��n-�.,�+�{X�ݐ����Xh��!i��-mH�G�9�q{#���s�K_���G �+��oQR� y�P<Y�4<<��<d�2��N�ݩ1rS$�wcfg]'<J�޽��q���鷅�s���(AQ���ǰ���q�X��/�ÇoR���UmV�zh�2L�6�iF
�`[��}�f�}"�d	�@w#������}w��&s�u��?E�]�����!�Jg#XU����48�Ю��o]��~m�"C�8���o�>����f��M+�#>~~�����J��n�j6H���#�hP��F����[��|<Mo~ u��;1�Z�����r�㵮�H�C��Q�J�zb�O��4\qr
b̥6���@����[�?�U���ë���[���i��S�����C�D�W�I-��]*�ADS��q-����ܛ���ɱ�3�4
�P�F@y�o��f��i���q��*�痨i���ϟ?�	���rV{�6��b�/�A�\��&����
6�J�[�)�<tOH���t_�n���t!Js��H��;AiD�*ixk�C6!y��ґ��j;�H�A���C�i�WIt�B���h;�+�W�#�#��<�;U%�^پ}�p�������KM���������l�M�gS���/���@jR��뮃tE���rvl9��Ձ�;w�<2���J�Z������} �I8�}���a���Jp�Uapz�y�S
�YgK���]Y;�I���U!�~� $��b�������$~u"��L�(�QM���@*^ �@%�|���VO�E�{q�K�&q�peUU�.1+�eH��ׯ�S[^�A����4a0��Ѷ�3Isss��I�����n�U��L��dû�O�K`
0�[~��Ͻ������Z\����3�J�C��ի߄cy^�a���5hp�v/$�һ���o1����3>~S̽4Kv�kHK��<����u�*��K{A��#U�,q�A��F�p_��/_�<b��)��yqG���l*7��!S9�|�3��M�Syyy��١�6y�Z�l�aY-p�9��(�c�Pu/P���a����o���:>�Y)5��+�����Ӭwi����{Q��7'v��:+
�`��e��I����h;���q���bR���ה8��h�8��Zx�2#;�@{VR�|L�TJ���ϰ��;�`����/�,(ƓwNӅe���.�������zw'��F�@�]����&�п�E��K��bYk�m�=o$~�v����Z���|	̙_4(l��]P�gzf(�5O��]sp�<A��_+޿`y��mb[�Ļ@�H������1?�Y��xC�T�8I�{����j���V|jii��"p�Am-����`�73�e�M�5Gr�k��)װC�(q�AZ(���IF��X?�����ڦ���ߛ�znF��|�T�jm)/݅(��oPRk�ǹR�)��-�.�m.�N[��0
����3�}�3��SS�S���sR������������Ġ��x...�q|暰|�m���b��� i�@�ZE�$��T\�}m&�յ~`�/��؎��[K��HB�����6I)O����[a� �fW�9X֥��?�K-�0��(voKB�C�fa�R�¢"�Q����X4-��/�AFs&d������Oi,N�����q0vA�[S�A7@��������p����T�Յ�'>��<�%����	�5G����@�^��簠�Ck��R�ხ{qϩ/�&��ri��A��A����o��Z��A�����e���t��U�Ty7}]"�d���%E�S$�%�� ��ڦ2{ %pC��y��d�ɓt��x�q .��L0�sw���>�I��ܥ!��2���s_�{����Z���!y
��c��d��v�TO!�(#�?~���q�ѭI�[�6�L�ي��x�[�2���fп�)�y��(|*ۼohx8�A�{k��B�H�3 ���ݢ��^>mJ-���n*�O�����!	u �&�8�ꪑQ�nkF3�Oy��bV��|���w)��]!$^W��_�ے�x�Sm�����ʈw:h[�q��-�d���4�c�ǌ+��XI>v6 s�>	��S�!��,?��B��'� 'ȴ�@W�3����?¨W�"ˎ-a3�6^��i/��+M��O ߟ�,��^��A`�&@{�d���]/��*$�����z$D<*y��Y�]ւӭH(qy#�)8'M�`&s�,��s8����ȐY�?텽�cz�@�T�'�PO?�N���da肝��Ŵ����SS]t�L���,�_u�ЏԳ����e������rM��f�!"����L�~dd�{��ٱ�լ�N- �gK�Ր�$v?|���ݔߤJmVUn�9���T�j٘	�7�n���c��~�[x=�����P���0{�g\�niS{$<�e��|Vv0~L�����Q���]^ᯥ��:�Ra�T��5��2x�"n���9�LU�cuʦ�eQR��(��?�J]ȗ8B��Q��]mZe�nVQ�F��ֺNj7�c�!��,$�4��H��ߕ�0òw�2{&�)	Ԏ�`��T�J7D��������A���(���G��HH��f�ڙ�/*DxvԘ� 7G���B`�w�^ñ#��ުQ�QȞ1S�=Ȇ��.������t�t����|���)��2��݈� ��8�8oEi!ߞ�q~c��g����:�EJl�}���~I
w{���٬����F5�E�T���ʐ:8dԬW*�c�j���j{�3��'��M�j`�cY!e`��|��L����y��ל���Z��U���VnOCc�:��p~����4hֳV�@��{��Mf��& :��h�Ε��B║a������O#x<��O�w���TZ�������p(yf�l�P�X϶��`���A�3U�I ��:NX;���W�k���f�̓��Ntip��(�/��<���S-(�
��>`�N����R\xo��US�T_���d����FPd<�-��zA������e�Dv�O�N>�/���iS����O?�aV[
�Oŗ��DY��Y�_6�1���O�<�E��ւ��ؠ2�[���4ogI�ߖW3Q4U�O�;�-�����b�t��Hp��r��Q3RQ�3
�]9虙�%Z��*p��3�B��S�
��@����!aaR�q�0K�&_��f�׳}��|!V�K��M���1�K��!�HR�VL�f��̯�(&�ίS�eJG����JFNJ�R'=x\U��M<n$�9��ms��N��N<ם��S$�Rh-aI��xb[���:�+�� �za�����ê��*���i�ղ�x-f��w��t��MX�$�`�L�Թ*?�(wJ�,R���s;$�e�qr������
Y�^�s��Y����G�=�]"���2e�]�j��������z��.��@��p�l&��SC����q�
M���V�g��I��� �^�E��jF����#[aV�*Z^�l��8��v&}�I��	�� Z&p�f��L�\��̖��7m�h^O5Ͱ�Ɨ���M�Sq�G���Ŭ� y:4�ߘ���En7�������FIkf�l�<������\�;�Bv]��[������G7|^���J`g�.	K�ӟD��8q�x���T�-��w+:��-+K̊��D �J�J�|��0�@ufP�,�?ڈO(\�,��Zȧ�c�gT��ʖ��^��[w�a�K�{dvB��u��E�Y�O�X��\Di�:�n:w�ɗ��ʞ���֖����O��H�/���
�|y�b?��J�hp��Hh�@?����,��>ګJrQ5�7;H�w����9.'S��hs��1g�"T(�q/�Ka#�e�I�֬@��@� �ݫ���n2ȇ&A%��v��]��f~�i-ٞ?�d����x˱)����G�����D�9T�i2U��l��9�Ւ��^ \3m�4�'�7=�2��\�R^���6Z�,o�*9P���1���Hq���y�^�d3_D�'Ee�kQ��㚜�.���:��v��8�M����Vh�B��R�M)���;�U�W���u�9���]�l�=g�IɎXD/�Ӽ[Xi�"�DX����5G�\�!s��K��:@�$�fޢ�Σv`��y�!rӋl�{c��o�t�c2+1m[ޑ 'I�U-�k��6���wM����iR1�гFUI�MXC��5P��N3Q �}>/U���X4K��K��	�h��&�� ��v뢀ڲ��@�]�Y8��0)��-f�Z�V�����E#i��&g�{_�]Y��Rq�z�{l"����!�d����ʈ�~c	�i���oIO��`e�Yy2�ɪ�n7n����̳_�
?O�T��5(7��?�2��X��E�ٌ�a��]���93� oS��(���ń!)�̞��u���Cm���%V
:v���&=��%7����'y `f�1�z[j��e�}FscЛ��M}�����V\��Դ������d���˚&%f�ӑ���a䲎H��b��w.�̯�F�$�q�$�yϔuQ��b(4��C��dU"��
�b��R�����sr�q��V��7��?W'���s�ϟ�'Q��Bc�bckU��fkkCV��u��wx��XA`:���Q5����gEbM)?�"�&]¼��]]��PVmE_��i&Eh�n�"a[V���'%�/zU	yD���I�CIn�\YG����Ls	�49{Gc{h�E��2��(��n����x�����!�5���.��s{/��n���p"cϪ��͐~����C��
B���<?��~�kW�x���ny=\+�r�(zxM}s�CP:�ϛ�������KK��2��b!�O9ҏ�p-�AξQ͹��|t���j�<�tF�q ?�.q����a-�sJT������kB�͟g�}��K��A��[�3���J�
H5,����M�=J��4�$N\��L����rT�w������zj��2�)�r�/u���eg7�u�1��ng��\7�`U	'|+%[#�
aD�]W�,#���K C�;09�~k^�����>Lc��H�n���ޙj�������Q��1�EV��7	y�Hl��x�W�i$�}x��՚�$����TeÊ/��M�!K�n�:ơ���"�
���Jm��#�1�~�p�@�b��cR�X�X8��._ҡ|։Y&�% ��|k������lǄ{��};Zm���疨��YV���x%`ɘ�f��BI˞r�,��/Jξ̤TӆX���e��q"T���B��u���[��o���D���Es���~V��k�ۦ@��>���Di�����	G��bl\���j�J�[픙�
�04�I�k���~��hX���x�|�i�ϒ�V	U��Ɂ`B0Y��X���Q��h���	%3��5�w�>57E9����j��B��S�cs��0T\t�P����˪|{=D�3�LҖ��c�0vZ{�߽!>i�8QLX��s�S[0�VH�����z���?knn�E��ץ�9�;��$�o�c�I����9�5��G��xצ3yx�z��������#y�Ǿ�y�n����kQr0+\������,���=�@9�z����_��r�l�6W��2?�ӻ0	W��ߪ�3}�***��y�w`|x���Ws�������hj�æo���\�:�����A!�SLm��;,BcmF�.]��!�/p>�dԚ?�#M��S��'�T���a��(O�g%{�'�S����U^���q蹅P9TsS53����ؒ���=b+�0�n�#T�$�*U�Q����Ȯv�n��ǜ)��Kh��r���P�����ٷ,��U�4n0Q,�	"=�_����&�������Z�U�a�3���-��_�og���3! �ǻQ���x���*w�?m+��=��v��҄�R�_d���Z'�2��q��T��m0ٝ�OJ�|���\�퓇"�4!�V@�-~���8ʅ*K��v�m�:�fl�7����6�PZ��|:2
G�I�.��Jrݚ�#Z�#��H��a������i�q�N-��z��e�$X�)�r_K�W�@�"�dz੎�����?�O�>W%�n��+�WL��=��q����%���Zʻ�BY��M?��ϙ�ϯ�O��m���t`J���p4��a�*�7ә�#�ݞ�<��1>�F�ULY�<�(+�� W.G��4��񚩓i�����=L�Z��287E'�Fhow/M�صkׇ=>`z4H�
A�/k�����X��i��#��b&#�,�Ͼ��-S�������~V���}6P�U�4(�w�ﺥz��֐sZs��֗��]!�%� �rrru��+P��	To[A�����\Z=�[A�D	�b�uW���(�6�O��md֋x����lմ��a�g�� $dp!r`wS$_����P*ݔ=.��?���y�w��w=�8��O
�ɩf�w�9����|��#Z#�Iw�k����m���J�I�-D�>(9M����Ip�S^��T�irz<�A�g�� <���_eJ�ٿi+�B`2��?��{����EgQR�l(�?��I_{�#VI�Xu4?P�奙	U��,���
��x,�d�<b���K�ӡ��D���1��;|ϻ�E�|����J������N��>smF�=-P�iKjvl�ó�>���G��4�q�̏S������ts2j��{Ks��N߉μ���~��
ٚ0�7"���+��o~�΋����^^���:��=��p��pyQ����^�ޢ��,�e��0Gi�]���N��� �_��M��&LG�D�;�4�`^�P�Y������h�[8���$��tx�2���YB���ԍ��f��U��<`�xt1��$ߣ?<i?�)�Xtn.~�7^c*�;N�Ñ)��Ս#�@P5~�6�X~���h�h�3b[��i����!RH�ZPB�{����lu��T�l�^C���R��9��+s��o��hYA�`�`��
:��}5��5G���C^7��J~�ی�(�ݞ^�>Ѕ%Ш���\q_/���`
9�. ��&�Wρr+Lq��o�މCS�Ķo��j�x��*#���a˥_�M��¤���/�fef!=�C��/sI��s�G{���s�s��{#���[a]?J�.��$l�a=�o��_����afg;����P>�4�1��g�Q	�]�ʳ�����F�{�8��`gg��Oȉ�,\0���Rv���wg����K�j�!D����-α��2Q��vg'!�������g�|�Iw�]w�[����7�|v��>c���\�f������h��Oފ�Ut���gNK[%(?y}ՙ�(�9aWCs�>h4-[J{�Sm�U�}N��f\{����p����	���a��L@h��j�uT��-'�W��,�y$��*���_��.S���x�lykq���d�b�X�4�V�?�'DF���|xA���c���H{�� �:�kb�"���{�[y^��;	��zXݬ�h_H�f����?�(�+vظ?��ך���Dn|��m���b��JRrE����4���S�������A�|�Ҭ��#2����T������*+�E۫f&^��
B�XVr�m\�L�*ѿ ay6%���K�bUg{�Vqn�^��QVfT�Zs&��9z�[gU�����é��c���S�J����
jw�uJ=�-Sfjt�}��~"�M�w�0�S�r��X�r�t���U����\5]�aJ��){TY��oN�n".`�+4p7e]��!$�����0���3��$���}bm��EϪtU`vF�.Wn���9ӎV��`�;{�﯅�?P��
��^]��4x��T#�>�L�U�c]��o�w&	�G*z�A�I�B�����bWt�XO8��9�,?��*WMU�Ȓ��'߾F�z�{U�N�����A����s��۸ڹW�Y@��jy��*m���d��������YXC�d�v�Bs�r7B���:b@���}��I"��?-���Mޟz��,���ݱc[q!��󷽃��A��&K�:~�^y��0��zT��cx�&�<a�i%�+qc�.�m�-e��|<	b֕�@yDAg�
X�_~OqM��p�t�N��c?���_�����!�eW����̯_�[���lpX��n��Y� +�z7E؝U�*�V�ʷk�Lh�7��:�E�&���"x+�&b��T%U�Rbx-��Br�?�p_���K��,$�|@���1�0F�=�Χlا�y�/��Q�g��5���d*�~���O�J:�ޥ�ث��S���ga���4�#���� �J�]�*	�����gj�1e~�;���e�����P-�������NE���ϟ�"8q�Z���
q��##���F�C�y��T�8��"D���Kw�����ذ��b{��O۷9|[8s,u�[۔	�P�Vib����Z;�;?um;��B!A���=#Y�*7�0c�E�2���{��d&�&գ����Y٭l��F�<C4Ԃ�!�gt9�׻|@���K�{�|�>nZ���FZ�ު�<��M����S������HN|���S:ZZ�����J��D�m�������X��%��Zh�(-��[� �$�,L��q��a�Eno�'M�A����r%�/_�Pa�����X��,���14�z�L��_	3�
GBc�9�}�2���S���؉y䠗��/0P'��YS�y�@�΋��W�����b��qc0�*>
R�3n��S�W���%?�{�o��	�p`��|dlaa��V�Ԭ�)E��t��_]��P(-hڊr��S��7.��i^�*9�:%�2��N�"nmSn�58躻����ܺ����.&�-�Țz@�e�^Nl�=vâuv6ׄ�S���	����n�;��ϲ��I�����3����O,~�r�"�#�ڮ��N`��}�I����8�*<u�L���U7�S^�j-���9a�2�A�����si�Ж�T%�jֵW��
��������֛lWf��9�T#����%�$���za��)֊OG�\�h끌n�>�r4M���W�׻5�c�l��u[���w>�}-����=(GX¤O�������W��ڜ������<�S��ڌ|���Z�����#�B#o�e������v�k��7S��|]XȂ�%�,R2H��r�@��^[���l�� T�����n���b��U�y�7����O�q�
�׷�+q��aD�w��^��C�w-�	��9�X��§4�����s6L�&v����[Aj�u0�w�eV	��ʆ�.��X0d8/FV��,�<��L��E�.w}�ڜ,f�k�!fM1�_�܃�2��Ҋ�fQ��t�5��d�ن�s2��.T�5M
4�m� �6�RP��Ջ{��llR����ŗ>n��� ��;���f���-�1��K������|�y1�(�����z�31�S���1b}��|�@�����V`���ֺ��`�KG�o�@(�X�F�I�U�Y�)F��F<��`BX�j.Xq��>�B��f��=�<��Ԋ�_@����i�L�uK��6���p�]ߝs��՛��7�x��i�!'�RjJx��%����Zg�2&��.g������VffZ���}lBB��_oaw�4�^xg�Tb��Eh�I���E�Ů&���cZ���C�i��\��+R��+��p�����h�����i�}�J�Z��C~a�D�����R�N��A�����Χ4�=,,,:������]^���1e����D�v�ι����=�α���%�����`;�=��V��5C�V�m�oo�Wi��ko�f%CW� `�P�B�r(���I�o�a�ݿ>g�"0|�s��d��Fd[W���V.m/�]�wh4Rt��R�����A��ެ�r��l�߯�U3-a	�'�B����RSS���������}��uQ�^���cc&���ס�4 .�.Y֝w�����(X�!���L�5�����Ֆنd��w]
 ��?��f���,t���R ��}=/+�Ɖ3#��I	����k/����q�Y���Vݜ�5��X�D�RN��|g����|�_�'k���1K�F0�zi)���i�ӻ����J��xv�eO��M���[ <�S���!�M�ϸ�f��)�M�����=+oy�}�$���9#���γ,^�]ap3�1�ݔQ&�t�q�_>�: 6%L%f��<#�c U���\��`#��CkA�lV�x̲8��%7������"�/��mϦ%�հ������}�.���\� 0d3����'?tp�%P�hk�=��7[K�S���,��O�R��RpO�
����� ��˥�|~9X���;;��$�����R9H���z�{@;B�\����<���P�up�O� _�,��v�Sܻ�&��5��LL�fH�n�� \#�)���y#��n�@���gIY�z1��|I_���ye�h�}(ZǾ�w����y˯#D��H#E�A�&�%z�k��''�l�2歐2�	��&���-8ǒ�Jg��Kc�~a�c5
�o1k�7���!����%��?js�*�n�����I/[āMD#��۷?]y��~Lk�D��q7Z�R��$q�׷Ma�@pM@��U�����!���xJ�~���,��;j���:�����PM��MS8k� ����ۅV��Y��x8qm��E*FN� �(d� p�h��vG4�P���J��S�Rq���yUx���UV��Y0�r�`�~�5>h�\L� �~��� �1��5H�A���h��J�P[��\����L�B��3�+4ӱg�o�+���d\hKt`I���~q�z�u55�e��-��8�J �����:V"���?ȍA&��2�v��i/6��Mh�E�pU ��_9��do�i�Un<�n��	��؈� n��*����V�L<�B�G���NǗ�=��[��v��Պ�!;���p�:�Pٟ�P(x�l��K�7<�����i�
0���:�֞�}�{���h�7G_�l�Hg��?�dE��Ç��6o;��qs�k%�Uj��Jom}~�-�]ɱ��69%ki���º��Ɵ�.z1�(�_Uç���>�F�Z�W�#��T�G�UXqa�Ǩ�����͠�r=�8FxT"YZZ
�n������?&������Y=�A��	9��던��:�ʬ��/ �:�q߰�5;ui��g���5w�����&��UI���w|�"�n�&u?|��,���)++KV��5��v��g�{+�(��a��[�M��r����I�_���CP����M��|��"�3UC!�$v�^i�5��7.v�(�SI�c<�����$���rb�A��w7Re5`hi�`|1��O��V^�pl\��Õs)�n@R���:��<��B�QD�̪K�?mt�G�k�oq���65��C�vJ6p���+�x :;8+[mr��C�3P$<B�_	��r�MD�Jha39a/C �[�b���
敞�$�*@�v�nn��bC�}�������s����8�Ř���<Z��q�R�]݃�� E��脘A��d1æ�G������8�W�U9В��vv(���Q�@RI/d�w����>m���Mp�$��֦0�_e�1�Yx�jk)=r�ު���[�J#�Bk��ur?�Ņ�Y=IT�'�`C7�s�]||U���[u�hk�T��ֆ�g�c"���Zn"���[�0`j�/2Z+_��uE8�fx�&+@H��d'��u��M�y�����8#�z�N��SM���'�L��E���0_ ��Q�3I;���Ҟ]�ګ���,���U�χ�T�V��ŋ9V7�s�W-4���w>��	���L�Nq���-�1*�k��614x�B@*z�hY�`;�j �砉�4� �Y4��U"����NtHKéu�o��i"�?v0RCr1��)q�{�ެѱ�b��.���2%U�3�0�#��f����5M.���S� �v�}�.Ũ_��_�E���B���� �W�h,͛U#;t�xW�> '���nD���V.���jj���_�EQJ>|���ʜ�
(��|\v��2H�'�2�PV�0&�f`KO3��s�K綗����A^����_CϦ�N>�Ry��>-[m��nݚ2��Qz�	��/��E|",��:T�	���}(�|q�$}��f��U����aЁ�<��	��gϞ�F���1��,d{� P�ak����B�`/�8�"��o��������:V�� h�d<Њ~���8�zl�"�ZLh0�e�Mo����{ȈW EDGE-����������>}�F��J��E0[�ѐ��w�tGH���)[K�i=��p;
J�~6���#A<Zɱ!��~��6��Br�fC����G��<Zꘓ��@�?�͐)#F�7g����S�r��� Lʒ2�r2P�	I8n�����N5�E�O�%
���D(�=#sm��%h��O���ww>!�9�Jg�h<�9�YU��Q����-����m�>pW���,M�bt2)�����T�AVV$��I"���H��y�� �����~'�NWd~\B-����A
c�.p��onbԤJ`˯�6��ʮT��`�ʊ����nm�׽ks;r�Uc�wQȝ��eQ�R�^� �a��@mZ�Ǐ22 ���f�4%�����9���s.Dg,�IjW=�498B��|gy��/gv����}�%$iuׄĻw�@Ƽc���O��#�v�*¹w|�)���O8�|�2**���^���� ��9L2	����s�'ԗb�[������L ��t���m�Ɋ[�;~S��E�h���!�}�����JY�Pk�z�/����Y[D)g8��t�0jJ���a���B�<��#9�]�~�2���q��G��U�gQN��~���I
P����V�s��=�h�b`��Z-�*��'�)�0p暫��;1��P���gc&w�����k�������p��Y9<�g��ۆ�i$ZOo%�� ٩:))	�a��(���;�Èn6~��C_m����Nw��Y��8�����!�&��]�G$$d��F>�cM�pd{��^F�W����5�zԞ�cd�>̞Ԁ�y1�e���P���Ǐ�N�ǭ՜@�3@�R(���|5r�W\96�����>��;g@�����b���z��.Z�����!�J#hR���^:1i��ō����kA$g׫H��YD6�
��p�D��=*�ZD^��N'�0�ݲ[�`�_�Ɂ����6o%wtt@ (j{�����KX�{ 1�f�V&_�hG���ȩ�m�]�~�c�0[�Mr���������Z��r��i���_��vHLc���/|!z�1��+�1!R�S�1�M�
x�`q��<�������h���j��l���uQ@+:�ʛf|Ĺs�V��������[��ϝ@U��:�YP�M�m�������P�pR	����C��*�%?�m���AKG��0N|-�;8wlHj�[8q�mm2��� 	JII�mLUKL�l�al�>6"(ʹ��M���\�`h�Q���-��C@+1̀����.f���)KM���:P;0�e � *}I2����9`��n����xP��Y�\��:r�c���	���.��<9��M�
���0��얕��cW���՝s gmሥ���6���-���� 1���V"�/�mY���_�Í@�&�w<U��ܳ�/���b�3c{"a�7n$��Crઐ����tƞ��'+��1������O�lW�v���q�P54G�CƁz�B�>��1����a�o"�m��,��
�BJ�N�Z��JS���|�T<Dֆ�:�'$<�μ�{7tl�wz\Mۅ�Nw������5cD�J�Jb�62� `�f�ՠ���J�*�2��R��m�f��Ӷ:)�2.��s�	�D�=� �OA�?PO�6ܰE�I	�O�t�f���w<F����e�e=J{�`	��2�geiY=7�V��{��V����SV��y�ӌY�_�|95���5�4���{3��x�N�6���!�#5j{@%ܭ�³!)����5u^��wE�~�+_��������C�9��9}��J�(�z�S�����q���*�j�W���\�#X�;��˿�l}w?4�}� A�nSt>5">{#Ѻz+y,�xr�����,ݏQR�KHDf�C~������n������n�-y���F�&�����ˮ%�����daR��ųsO@�	���\���_�8_4A��0L����!ن����E�����? e�=�{b#�=X������P!���ǰ��,��I�ٿ]��XT�fgg?�T�<��a�ʠ� �.}Y�r�6��R[������CI �z�^=/=�������h��$���߭첲x?�#�ːWz�lT�,���y^v��(���\���SyI��9�ak�-�4W5���G,d@����Es��'�y�ůQ��ړ��@��p�N�&w�~.-�=a��.ʊ�&`&.u�쇈f�+���(�?~��U�Y�t�@;IF�����UǾ�e��I8�L�Hܦӈ����n.55�p���oXƀZ����2�:��܌
p�=W��o���I����𫃱܁	3sm��X���IVsgY��cS�R72g���j0� �O�p�]��ҫ�]XRR�g�iQT0Fc�����Hmmm�3dee�v���+`ԓ���쾬���|O`�"�"��^ۼ�/����LJ�v1o\�����������ԕ�'|� Uo3]�¯�@��ެY�.+˥�E �lލ}w���	�[��}�&��+����/�ۀ������I�=s��K��%f���<op˵k}$��>2��+C��v�c����i�BKY��R����>��	�9����8N�F5��8�?Ź�(6Ѭ�$x ���˱�
�>�XˣtJ?|��7�����J�^)Ֆ �ĉ���G�1������CI54��	q�������������B���o%�8�,T
:�S^@�t|f���8��w(V��Q��D\my �9�R��ح������k�OX����hK5���Β?1j�l�j]&��Kr�0�����v���ZĊQ���'4��8��=t�����2�L�ؼ�ƂN�tڤ5ϫ��o�{,f}�~�LW�Z˩G�:Tol�q�w*��+��tm�ݓ�Qۛ�������Sǜ�n;������|�ϯ�"�|������5) �gP�|�C�F�ǳ�V��Ro	�pDso�L���ZaR��!�ύ��P�/�_0�=�-�'�MY{z�|h�7�
��J[v;o�b=z�n��|`僉I�^�-������$�Z��A+�g��12t:G&�ƿx�@!϶U�v23�:�e��-Ӆn�'�l�l����jR/k�� �G�Yv�uX�w��<L��[�+�j�vT;��Pw׫܀%�Lv�B %X����ɏ6�	�`۱��r�����㡉����Wr�o@NV��~޲��|9��|I�u��Kw��rͅk!؁y�@�;�D�9qO��x�]_О���ej�>��^�f��Ce�Y��uZ�Y�N�z�~ {�1��D�!�m��OT�:�0�-�O}�:��`�*+�](���
�ﾔU{�a|�t���:�w����)g�oD������U(Z�5Q�����Ui��)?��G��k�~� !`;Q���F�K��d&�YAb�Ԗ��ă8Q���_�MD�2�X�}�՗�4`6{�ܤ�{x�A� �x�fkи��K_�fW5��'�_tI�y��i?�p�J�?ҁ=wJܺi�7ϳ�[sz2P,�U	`*a�@���	�8�<�pb�e颃������+�/�й���ZS�G�^�z�vb^�t�_��`߼���eq�ѳ+�/ج6��,�@����p����}���"a>�I5/�X��W���M�;�}��Y�1I���1�Ţ�vp>�7O<�Ϧ��1�ژi0��z���?��G���������c�l�/��G�����S��vڟ�⎯����Q��������9d���D^;�J�������|������<�o�kZ&�������_�/��K7�6B)�A[�/h讠����@�P���}��g�J- �^�B�6~͜�P�X�`9C�i���q3p��'þ�	e&�xb��2�߱37�p�Qt����كI�Џh�?e�j���Mm���ل���I_<�`�3saoV�h�e{�ɼ��]-O-W�����հ�0	ߝeb���vU	_>�]�2��8YL��:Z�G�gD�w'�� �c�o<�G�`a�u�xV���n�cYhe��s��r�:ߕ�|t3�וo:���U�wa���d~o�-���.ly���gWT��z.ݷ���6%��Lɇ|o��°)*3���Gc�iP9װ��#S	�2���V&QJ���Ut��kv`�[�����2ye����
�>q�>frYn3a�7���ٵgΖ$�sjM�)��2�u�늹����bK���yE�Y�-M*��^�*-�����k�/w����G���?_\�j��W�9�+#�k^s�:��K�Ŏ������#�]o��wP�e�����x����H��H�
]��u�k�|���#(�2N3 ��0�������Ҡ�����L��{�x���oܒ�rJ%���J5e��TR)�b�(��3�E%�i�u*E*[�)�mB�uƖ���e�>�g�,Α~�����������i�������z_�}���G���)��d���$10h���|�мM��v��9A!��Q�i���(V�7�^��ϣvYN�<��mڸ	!��s��4�.�	E�\<�dA��^H8�o�%�$P;۾Џ�OP��2L_�Oh.L���DJ{��c-���m)�+��f�)l���\�/k=��&P�P�W_aV��F~��K_�N(��´P�˸7�A����&)Y����6 �(��ͫ ��H�}��
ӹm2,�Y��9��H�}M`E ?TeZ(b��h������J�s)H�������p�b��X:p1�b�S˯\8��w��"	`�&ȸ2�q˧�o��P���Q�7�!�
�jQ�B����J?��B�N���ݤ�ϖ&�����X��/D[��y����:��ꍖ� �,�҇);%��%8`�;�����g�>}I�`�'9����N�ǀT���C�|�%��i2��@2m��3�ˎ S�f���&��G�B�	]I���k���mOd���S��3>�~��b�5���oTo�^8%S-����Ya�ԫ����D(2�~�
`������7���@I�G�Y�6}��`%��V*Ӟ�h>�(�=��P�N1�	_�A�ΐ����g�,L��]`��S��s|򣊸yH�eqA ���S;��~!�a�����29��0k�Zim�Ef���S�4 ��%����%~ZP$�b��T`��~5VZ�o�O|Ԏ��*0hC   ��ڝS̾�`q��hq�{K;���~�wp~�wp�o�'i�_�|�w����������������������������������������������������{��m
���s%�k�~Y���5�?���HCW!E���p�Q^4B6��������uGV~�@Q[<kUf�4G�3��s��6��iD�O~}�B���C�VJ7�H�bx��+P6�Sc#��C9�ъ(̋�Lg�t�h��FЇײ��^�����J�ݏa��\�Ջ�I$K�������TJg8��� ��=]9rY��^��x�@��N6���2Dxh����t�bΡ��v��xy�I�"Ngxe3��z�57�ч���>V��q���_?�41.����M��o�_���DD]V�tȶ���m$R_#c��¿l}bA �Y:���,�k��5���7��S��mo��(���5J��Y�U9�yb�*JR2�͜�,�p�~����س�dϽ�L�`��;HV�)L���SD=L�)u�\z���Ǯ�La_�H��%�ӑ�TZ��|)UPĥ�6w	��wiQ2.w���f|��X���$;��^��p�z�h'�?Xjϴ���D|�	�j�~~m��pL�a>���jė>�{��d��]3� ��|�6ᐇUX�2�9������-ԑD�S.��&c�B�43��GOM��̡w9�y��.P�p_�2)v�~��rťe���1�h����S��_<�߸�B�	��zǇ�rG�́�m�Xť��TN�E��q��D�$��R;��<2������	y���]7���K+m��# ~�5Ц�����%��>��[f�[w]W��~6k�s�O��n:S0_=�����N�2;'�˲�\���a�5��Hx|6��3��;+OmN�B�s yu>X�.1'j�]^|�ΰޯ,��8�����4�<�s�c�nw��(�ۺ�t� ���H���>-�4�L�sZ�I^������m�u�v��y�4���үc��^��x�na7g�sr8��T�w���������#5U:#vS�q�v��fAL���J�	� ���#6HN���m��ə�ϫNڕ�6��<}�mO;�_�����"���W���ե��h�p��٬�i�N0K��Oy�U(^
ao��h���k�|���T��ې-Kt���r����u���M��iYa���Æ�v�����X�Y����jrS�W��7̦��<

_���_�s��D�Y͆w ͜Μ���K�&S�!��۸L�{�i�����L�a��]���;V���	sl�=��4�u�9��Qng��2�����6�X�ι6�~
9Z?��j�ŚAt*�����6"���J��0XQ�c��'����������"���c�]gƻHb��ױo5O���o�5h�I�OIh�0*�����ϡ-<�~��	��2�o7t�$�nz��P�����EȊ��Lu����S#=�a{�j����L.1x%�J�����cǸ�z�j��>���1n���>p�&�UGU�~)�s���ʄ�u�Hq��M�@8����w��7uk1Z[ʵ��818 FY彌2��s�������j.�"u[[ͦA�%.�+�G@�;�+^���)������"O��рI��3\x=,��~5u��t�*DW�ϑ�=/��t�(�]����E׳��CJ�'�׃�c}L��ȿ"��3��ׇ����<�ZVH�ͪv_HvjŎ�*����I��Tck�}�� R��H��"7�qe`��x��S-�?�$:�a�Y������橫_�X�1ӶZ�g�OA�� ���9=�b}�Ž����ӿ��8~3`L�>�[A�0��e,���렞n���4�|C`��7.c�����4gNU.����b�V@5���%��?8�!S��$�@�D����~�Z��������^[P�$���Ϗ�o�w�G�ȫ�7�\~lԥ����/3�"|E�(�����K��@=� �׆�u�����=3�3'(��BE��)�d�m�S 6$�Ћ�M)# ����v�G�	_���:3��<_	q1k�_��8��P���#���S0���z��:J�j#�P�f�]$��r�ـ���ˡܠRfTZ'�_Dz�'v_��?�+���o�o̎��9�<*�˰/�B�uʸ���t:�H�V�i�FZR~p.hi��k�d�9�[����e�EA�ňA�p*\s���ݰ5�|�V5�J��K�|�8����"��#��B�Ǜ���a�4BsGoP�����"��_J�vm�@���N^-ř������<<T��}|�*˂^�@�9���vA>��ee�r�ELtF�fN|���Q& ��:��,�ǿ�DA~S ���Q�+��iw�ŉ���9�s}Į9%	s��]<l���� �B�E��/��$��*�q�-�9��a�� �ĥ��?T�@Wd&�����-�z!����X�chҙڄz�E�5@Ĥ�}p��ȋR����@
w�b�`웒�j�e�17�S��4��p��wegHF-f����*�@��o 5��@���`�*�o˻~x�n��5d�]�/d�.���i�X��ߣ���"
���jIWM;��K�O\ ���k*�T�K�sj:�p�,�%1v0R!�\�h��c�%��!�-�(mW�o��?A_SHṞ]���)�٥�/:>G�RP����rۆ6��=:|���x�U뵽h�jʫ��d��R4��ޗ�r��w�d4����Rr�;�zqQ�h���ה���T���Y5V��g&�=���qB�)��)|�i�j��8�Z�У���I�j �G�k/��v��ig6H��`�"3J��<��s�z݂��K���Ik�Z�I-=��,����]�!�����íq���`Y��F��Y�z}�ǽ���m�8O�gX�y�k���wf٠�=�II�,?�3
X\��˹�����H��$;tȰR^�vט�7!bbF�m=����囲�x@=o�	b#f�s�/+/ۖ����YC���E�w@�-"�*D��IǍ�і�>����6���qc7���Y���}�	�m��9���)���(D�5T��ܿ��6(�sT.�yB���ΩjY��~���#ƙ��Wp_5Yb��O��x�bL�������m�v7y)�; -�E���t��=��bEE{hi�
�]hDl�c%@��
D��1p��>����;cđ�M}��H}��'OL��~���AtGp���. ��w��{�\���)��(�b�����X���t<�������4��uF���%{�M�4�4}���>�M�:I +my��L�w_]g���f(,���ݏ�KNNb4�B��zg�a	���[�KS�/�)�
,����h��o�S�����������:w�Z�Y�ET3�n�YKl@!ˇ9��/)Z�gݺ9��\���E[�����:���"B81��AS�H�CN�vD��V��gsKqN�Rȋýge�:2��N�_����9�H�*4����Zc��$���$�69[�^h��÷a(�>�dN����O�!��"�g�a�+n�,Zn$�e_Vۦ^�v�A'�o��i��_�[z]�Tq�|�O����.U�~��z���e"��-w�}E�q*�'�J�_��2Rl�ðq�B��GU�sΒ|�$���
�a�(���iU����e���A�,�L��/<��c��ayJ"��J��/3Н�i�3T��]��8ǘ1LF��]�w��3'�H����PA�@"�ɬ���51�'֥TX:v%Kq=��ڵ-�B���$;l��&U1&�2�qx�������M���"=.���p*.]�	�bw
�$�jċڧ���<%7UqtB�;��»�@�R�츽-;KQ5T�hw1��VIy�8�-�c(F��_��2H:�Ŧ¸��dp�l�$�7"�I�W���/�d�-���^wc	(���ަ�1�n-A�^���A���o��f��!9omKC0�ӆ/�a���.F3UC���\�U���i�)ͧf�U�\�iZ����I�g�p�]��Lݼ;.����ʣ�T1�������	����4�� ��!���z�9�%�5��0/$�R*Y#-�e�����F4�BP}s��~�?5jԾ��5Y�U��M�LuOdl�&�a�*��x��O���T�:m[��j�~�J�e(=K��g�i�\P���h��z��g�d&�s�&U��hH޽E���?yaQ��P���[q�-��� (ǜ�?�������n��XzME�{u�J�ؠI9��1	�����D��>���Ɏ��NB�N-�0c��x���ƒc6�*���| ���j� w������n-P6�G���
ɣ�O��8�ml�a@i��Q����ī���^B/�)�9YG[Ǹ�;Y2��m^�ɦ�'Ҫ݃�N@ �TV�l'�'"2C��uM�Y :�m�<����3���sQӂ�r�C�<�q1�`o���0l�5��{�k�VFJ��b(�5�����[�yy��< \)�v/��'�pLǆkiDnҙ���ܳ��(j� U�ޒݓ��&��jS�q�T0�<&��nq{��΋�Ĕ��W�B���e�L/F}���,	2�Xk��v���������L�9Uw"��Δ��n�J���.g��b}�|H@X�B�Nُ&����(�u���-���;�hB��iZ�9������⥖l�/`�GU������v�����e!s��*��H�H��/Fsr����T'EF0 �*�j�;���Q^qO��ф
��ײ�"6���{�K�§���������WxA�"je ,O��Ս8q����|N3�I|1�s��l�o�2�|���v����;Ыb+];�n���;��®�;�
tl���9����{u�j{s��\�397�004�p���:#r-+6{/�ŌL]V��!�^_��Q��m~���:\�2jpR�{��Qo��L[�i; ���u�@�0�g��=�.hF�?ba����P��CuQ�.J�������g�%H�yM�@��:ř��o�/!md�p8)Q�������*3�/%��yۤh!�s�y%�/���y;sNB�㬉�<`�W���-%����� �y��F�+���z�G����@�Yo"i	�.�����
Ԕ��S$�<����/";.�rކo���ګ�{j�X�Y�1)�J���g���(��+�洭�u�'b�:L#��X������Q|��h)ë�9��Ԫ��2/,K�;Կ-H��/���%px�J����w�5��:K��'W��&��X���N��g�	������N�����):)�褫d�F ��<ɸ���`�AKE&��:ܗNNm	o��}����������.���k���r�W�R��������p�A����$�p�.��\f�Z�r��|D�w�(��'����4Ru.#5�;ʤ�Y�O�|Ǌ�:n��z+��ͅ��#��]�;G�]���Q<�qɺ3㷘��a�쥕�=łt�2����?�mݝ�	y�QZ�oa�7��7!=SB�{Y�6�]��1�N��h��ӂ���dj�s�2�,F|f��ݐq��:.�~/��z�����VP�ʹ�:#�M�_�Iu�D3�4�����3�(��:D�n��f�n��)f��!��e
�����Qǯ�-���`���8jf�50����d��t�I8�b����(����ʥ9�P�)mݮ���o9��:25�P��xT����Lk�7�nÕ��`P����'�.MOs�
y���0���P���R_H1�HD������w��^�Bby�=C�����"偒���"Zշ-�����Hsu��I�@I�/$~�PV��sؠ��m ;�B�~N�W�s/^�I�����c܊���ͥT�%E�{�ݓ�	K������.m$����+�D�%ԝ�7p�(�����e*TAG�%T�B�,Q��K��ė*��>��R=��Mä�z��p}�Uw���pk��6oi!o6���t0*|�0����72�v˻P�豑��qd
)���:w�A6�Ie8
�	��d��W�?j�&DC��=���S�D	��(6��X�����̱D�,t^IM�@�&�sq�4m]vn�$q���3��>-����%��0ﺕ(<94X
Cqؚ�*^[4�1B��?_���(�,���{��Hɮ!�`�)N [�}:�o9(�~�丨�f���j���;l\sN��Ŝ�'wʍd]�utRG��W�@e�&jw��� �o�Ȓ�p�\E(��C$���X0�%���k�.(\-�°#�d�Z��W�D��L%���|p�rH�V�׺@z�9��IC=��q��R�9ւ'�w�gC� ˢ��kϱ#4��Ӏw���R	9 ���AsK��8��~��p"��^�r~��&�G�����J*�y����c�biِ�.��6.zՀl�9���L}S��zGvG��f���㨨Y=���)�=8P;Tҳi��������f��Hk�R�#<��.��8�~;+�ь{�XdC��E�bV�I��2���=���^~�E��[`�q�.�G{��Nr�>Ms7a�6�Y�=���4Ur�f�Qn<�h>��`�!������!#�92��VI�>��u�*'�_/D��m�����A`�f
����5a���힡4cƫ�0e��;-�y��{?�B�8�҉���x2��.@�\{�������~�g������>w���\�k�9\F~�E'B�:6����T�_&d*�sZ�p�t��C
����M��!?))�;���}M��	���/�Mw����ٗwiѼ��[�1Ka�6�C����{7��ן�ߧ����>ZIH[jp|�x����p�E����ҳ,�C0wh���'�c{>}Ȼ���������m����"�sE��&��R�q@�8� �gԖ]b��+����U�x�mu��K[G	0���1�A
G��"�dA)>м^��&��Rb��(�ҭ�#l�Ad8qe�j���c����='�%�h>
�y�J�5��@�f#��̡��/m��WΏ5��ug�.�o�UC��Bԉp������Yz�Y��c�/JU�����r�u�Z�����>���x7���X��ŏ��qW��P��3��E#�4���0^g8Ҏ��Ҽct��Ls�E�)�h,��j���ewe�'>�=���?���w%�*�C�'�x%ځ{�ۛ�b̧?�b��X�DV(,����<S��zW�i�46�0�M\��o��D�>�e��33�����o�y��e2�f�W�����R���q�鐎!���M�^e:wWV,�l}{�w&������գc�{�aJ�{���VH� �)0�繯�`O��_4zNZI�?N'иi ��� Z�����!>�ɰ���:L�M������ûs�x���2�����<�1��"?�C_+�"�2\���Ow�-ǹ�0��̡���0E�V[@��ǘ��ߓ5�)�|!��У���&YT�@�X�%�-��-��d/o�*lx϶p@k�l*�e��/o �Xo���B|0w&>X�Ğ��y�b�0�#	X�����v���G�NM k�i@Й�QI֘�X�O����
��4�Qݍ�\����S�x%~"2 �C��U/�<b�Rǥ-�/�7����_%{ջjX~��3'މ��*>���/���%��mg���k'|3�k��d��(qs�H��T��縨d�e��&���T S*�����6E����j�/�� ]���������?��N-���Ŏ����-&n@�U.)4ShI�w���Q�D�+O@��
���6lQk�;y?�r�QCn�ܾ�*�����ȶE*��=�߹d�t�m������$�Ћ�G��+��x��(M��8���]�Ǯ�)E����Q�Gح��#@��_2����yY�}�RL�7x��,��q��I�yH^_z�iA�eJ�e��L���D�������>��oK^�X�Y�"\x�I�5�glEwe�ͅ��)B�]U3g�%�B:s#���|���e %,����vձ�p;�0 �T�y��@EU?������3)v��V��4�C�V�@�L�	��7�I~����奬އV��ND���fe�$
��Id��M6��[v{�2]�eH=����e�L�:a"�e��qQ)p�7
卫�>����/1��1V�Ά�Z���)�ÿ?N���k�ȶ�.$S���+�i�=|�rʜ�N��ܑ�X���f��%�O�'�y���D��e�
�c�2A�E�Ih���Rs��lM�"�����RsE�!*`Lվُ"+�����c"���aA2��==�q/����U��2n�\�{U��9?�q;�����V��������ʊ���9w�_v������ʒ�~
���{�oi�?�F�z88�E҆�	� ��q�4n�36�q�h�`�10�.?��L+����~/7M����@DD��A�����Cs�KY/����2u��@��V��'����8��J����l��"=��h,��JG��#�hȂ��/�ؖAM4�a�#�#��j�(��D9RM ��1I��$�.���1�Q?M؟^$�����o"#p~���p����u��!i$K�X�O!�RX*�=�'.�)�R��#��;84�L��`�۷x��^XaSH�Ta���DT7٭Ӧ� ItD[�~�fagط�����K+5P�e��R�-�=a<���Q�D�$��	��
kl��v?y�����y�SZ�ea�;���-�ha�v��.�x����G�#�-�4�`��y��J�n0�o�H�Ⱥ+jD���[��5��(����cc�A={A���:���HKD<N8�IͿ�,�c
�L��|!;9�����C2_i3k׵u�L�B�ք�NIe]۝�2�KYk�K!�+���7��^߆b'Y����tCfdA�!9����� C��=�	i����joGp{n���<�#��솣(Z��w�a|:`���k�~�5���%���j�Q�hn�b�mD���d����DF�f�bD���>�>����`��6�2�>��!) �Aݏ�����~J�zV37>0�4�DnyOV��<�6q0��观^l=�3��v�Md�����(�f��D��<^��pi9��Lj�w�	O_��?�}��y-�^%p�ڋT���H�G�������}�q��a7���`�NH���_��
f M��Հ&|����b�p����+}6���]Z�m�,3t�{���9��&�0��ɂ1��D.� �H���`<'�N������U�Xd����s~Ặ�2�C�� egJ/),EI��.�l.4���"9��FH	����Q�=�<�
qY��H�ߩ��<���[ۭ�kW�R�o�I�r���E�������F��k���=�q���t���0��	��7��#�#�f��x`���_
��([M��ss 0�=3����q/�;;Z��~.�� XU�|Ax�?]�G�塹��f�w2�0��ć ���A�(�&h�9�H>�x�>m�JMT1���޸vM�gH�`�J����?���BY<K�ё���ĴIÜ�m��;z���泏}L\��SI�]�Ď��FD�����o?���Ə!H^i��'�^#��=�\�����V���t��V��t���*ZH���*����*e7���e0���˴�r�?z�]��!��D��Mz��V�*��<N�^�4�9Tƥ�O.aR
��*�A�hI� �=,
#� �r������m�h�n����6Hi�����w�7��|��Ț�oonn�<�E�������z�^x��-Ýek{3��޽령Rn)K��(C�Z3��N}�u���q���_ļ���2˅�L*���b�x?�̬��#�1x�z
ű�F���b��g^}ɈZ���Q�{1��Q�ⳮ�9����N؊����Q�	GG������#���%ƿ��~���[��$��p����
�09��l���A�1m�y�o@�Y��������"����;_�-e�KL���1>��ړ� `���Z�v';F������7�����kV�A��9��PdR���`�Am��ɲNN6�Nn�����Ci�L�k�a�=t�Ui����w��=�����T�֖�-lQ %���L���A��|��Kq%r	�g�sr�NB>����K�I�DSɠ'A2��/l�w���v�6�8}�y�Fy4//O�Vw}pp��Gy�k��i	EWG�����`�F۟c_�`V�54p���`8�����8����J�'V	�E�������{��@��`䜩>�=��>�Op�\WEY��qሻ�cV�z��a��~Ŭ�2��"~[p����J]�"����x�dZ�<~��Q�o!��#��f/�,�R�҉DU�,�9*)+k�s��l�p8�>���p<�������:�杔ɗB�L%���/���!-�x-����R	."9��}}?w�NK�Q.\�����䇬���j���\�����
|�E�F����脪f��2�/��W�X����5��.=_F���c� i�=���64��٩/0ht�1�������8Y�w�ߧ����
7��z��}[F�z:�C�Ο9Ӌ\"�]~��-n��,q��fgeg���<��ݚ�X��ny��gч��蟞�=qB/vGttt�c?��0�A8q�SN^�W�}��+�KVVV~o����g��}|����zj09�Y͈L ��T��<)n���׼�u��C�>��yk������uf�`j i|a��tt?��`煍����+++�h D
_���s���G�LM�������*'2MQ�����Q���&D�=��J�9���'�Ffgee�w�V�9X���>��h����4m("藰+J^�|G�L�e�P�'�_����eP�[�U5ǚh�O���W�ÿ�,����u䘋�t���&k�ȃ�� ʖ��j��/~a8~�/V�����?HJ����M3:�|�� �����lL�Dΐ��s�?i����B�����_�ߢR�`a��2�A�v¤�b�U��V]��zig�qI�n��u]
GU���s��j�ɑ���8e��3m��u��*`�Ƕ*}f�ۛ���ɕn:d�|����9��Cr���1Z�ϟ�9��9�&d��2��7W�k�����Nt@�*��Q"���p``�/t����RcS��&��C��`�B2�d����G/.my^P�����`©����쯥�p�Z�
�R�=&zIkruPgO��֦c��H�B�����d��lȉZ+����П5�	E��rY �>��/w&B��
��� Ͻ��a1�l��S�r����	��g��W=KK^�t�DC'�����/_�{�^�Vk�J9��zȌ[�⒙P�D���v��W���x�Ģv2�k����R��;�!% �nX�Ӥ�/��_�τM��M~���mt�T]<^swy$���p�e���>�2h�.�?��j�����._:���L���^��
��bu�;lY~�������*lpM�>����\���+SI.��72{&���r��4U��+l���>�M!��.���w~m�VU�H���HHpb�e�?3�溇�,n<H�Z�����L$+��q��_����Ҳ ^a}o���H}�.�+E�_C�oY
�B���P�BavC��Wk���s���UNٯ��I����_`(�h�i z������7&:��V`w@���do�H�����慨¯�3�x�#�J�v-\��4�M��oi�Ǯ0������t�[ղ����Ė9�*Şw�{%����u����gWݩ{����Y�|BR�b����"�._I������gϞ�6\UVV�績�����[�B���������`a�Zn~�Ⱥ�a1Jf?VՍ$�]�� ����nXM��tｻ�>}b���7�H�0�k��H7i[�� o��7�2�OJ�-M���O"��o6�JO�l���S��B��TH:>KM�e��z˰�"��'0+��g�u�㷡P1`��m����k�[���B|Ѕ4��O�n�"��j� � v�����.@��7e⽓�Zi� �J���jwru΀��=���aȍ?I�\kn^�g�X���g�ee�K�w�hW=Jg菒B�Q��ل����M̉��&��{�_�����{_�*�:��TU�G��:}�g�I�n;�ߴ?W@����n�YC
&~z�a�^��:g�#�[r�/@���q^{k?E�͊�M��|��n'��^�%rU^]ũ(��t���`w�z�����n>�O�5(��@�����5�:��w�#�"5��C����L��la���-j�&3�[ FA��X+U�)�s=�*6��`�%8И��U����7�J�VΨ�}K�L��;��4s`S��@�T��y���j�@κ���yU��8qv��
�S,`��+�)�J���>�t�k�+�9����v!��SRRR���x�ۧm�s��g��6r�k���h�`��[[[S�q���N���S������}O�Be#HZ1ۜ����@ྡྷ��e{;���C��1���/�����G~��|�?�\�����8�c�̳� ���747;�S(Y$8W}\�1򐼱M���Tf�MM�н���?#3�y�4-��ׯ__P��*��s������r(���������@�Bc䪩�*����� o���9��@���5b��.��1I�Z1-Wr��'��-��Ϡ������s���QC�*�Y��UG�&�a�	N����N�y��U�Ï�{��Y<ӒY�?xz��7��S����p�Tt�����@:�k�`7+Jn`�J�a�W7W�c=�U9iͣ9́Y������{�p�C>�7���`�B!����6���X��̮��!�_���I��1���������8�8;k`���a ����m���Z*�GG��b[[�m��������|��w��SO���� �9"�FLG����s*�o�����k���GH�S�sw�x<���&3:��SY��zj���@
R�b��4ȧ�-�[��bT�Y	*����o1t���@X���=UH~�k5G��^��m��� �Z��s��\s��"q�Q
/��݁����;M��bʁ$��;�KG��|����&l)��啕������;��w���c4��nQ�r=�� �a�w����TǴ��A�"fe-��Ao�������oA���<��T|j^��W����D�x�7)��i�Z�2�>i�%?㪾�~���bm2�H'-w���V�(_wj�9���]�ozNk�~���u'\6�-1p)>�K�`b-P�j�P6$=F�=�V�/��}��ԞZ���ϟ�h�S|�~��3�:�����rR�6
8��;rqs�����{gX���G9* hm�����v��BP@Ab���ޱ���f���L!�tf�	��s#�P�x^]4�n�����+gd��g�Z_��v�K�Ә@�k�;��C�ڣ�㴳�3��tO%r6�P���xk���qq"|�1N��|����/���Z)��+ŕ_�Q�Im3bK���\Yed��L6�y�!������|�7�\)�(����nG�L�}XS!�EDFTX��R����)v;gd�_�<�������nzv6e�,�@r{d>�譓g�^] �l��(.��SI`j�����e���4���7>�8O�x�?[W��g�猩�.�h�dw���O9�ŋ�<�ܡu����x^oՌ�^��[,�e�����0#�:)imu�Hў��tB�����8�Wq�JN=:%���x��K3&��r5�6�N�R��:�s�Sp���Q��L\΅����5������wl���w3rG��6(c��W�Ő��Ҡ��*�f��6w��u�b�٠KQs�:t��.m�&�Z.+N���t"�n7��ߏ=���e���L���?���1?KI�~��O /T(���qž���ԻSR��-��7����u�=>��ΈP��G�ֹ ��L����M��S�Ug������G�&�s�,��p�x��^k�@ħe3��9�yy�#��T�4�R@Eg ݞ�ǳ��P���.��i	���$��$dFH~����s�Ң�������O����ƾ��:��0����,ZY�N��ܝ�f�p,v��]Z_�rT���
�~���?̤��F~�٣�H �����2g��bc������5���c�E�g#fL�3��6���PE->�r� �*0��3b��]����J.�����-���<-9��C�ogtg�C!1����+uoQ[̐&#�f·�B�0��j��� %�6��PǈcJS�t�ڇ.��g���U�Ote�/_0[L�YY���ba���λ����U^�_�Z=�w�!P�vB��GϨ�N�=�� h�k����퇀���,$��ܤ$p ������9b�5��k��i�a�ȑ��ܝg<!�;W�X�\P�࠸����K:a�`j���Dd�B�d�G�w@�ƶ	݈��f�����3���Q���Կ�˽��6:��V��@P�O��O�&%<��g��?{�����'�o͍�+u��}���S6e��
����n>EN]&���QŠL�9�I�YaU��75Ey��ϗ�����{�7��2��㓔��%���O��$���Г��	k&f�ӵ���Q��H��;u0�*/[���Zx�5"�J�G�\
��;lr��@����8u R�TR؀Ϛa ���Ѭl#��Ġ+�A�����8�8���1]:�CRb'^;%�$�W=?��mPJ!9MM;\\R"�m��x�tS�Ё���=��;���{Bq���M��!%�1*�n%b끹zyL�k�kr2�?"�����.��d�U���$��`�q��I�+a�w���.{Ѱc~�M���b�?5̧#Q��̾G�oke�C-:�X� 2Uo <�$��$z\�C�����D9C�J���X�AR92{�R����ѡ�9"�7	�H�'�8���T���I,�r�������:w�"���L/��q��s~�� �sv���D//���Ass����5g��JY�AZ���QU�/.yo�Z�w���&o}�.H��W�	��(�`��:j�84��
zh�������~�v���ڒk�kd¸!!R�n�|�����HVeb��6����᤯41���9Z�n��hzbj����ֵ��=�B��˓P�E�~wK2Hv�;K�2�Ν;����Y�L�*hp̺6�!�3��?����w6X	I:::�[.�R�rJ����[U�`�F(G�l�P)��p�v�zn��	�z0d�g[V���>hf���چ�;`����D�}����|�,���?L��y ���	�=� w���P#O��yQl!��Ri4���f3�n0���7�RZ����x׭j�$FVǖ�"���Ƹ.�%L�>@�_j���L�m���޸���<���_�b<�����m�������~�CW���o�o̴�x/ڒ8t�ژ��y�ڿ�YRR��^)���t�͑B2��z~S$d�ſ�IheL<��͗N��;G[|6��Y�8`~�E)Dxccc��`�����W� �aP����<u][s��%7 ��IW�k��t�� ʷˣ+mX�@)�X2����}�G
tX�����B�(@R,!N��7��9
�Sx),��
��
�����G���p\�re�-����ij )���^�w���3%$���� �{m��~∣��_e��Z�ּ��t����_�#u+(3Oz�6���r��M@RC�t��}�3 �k׀��}�o�)%�`7�{�f2�@B|Lb�N����+���d@L��u�J Z�����H8ܭ�}L@}��`y{��]ףj�u�Ha��w�����B�	�j���ڵ�Z�;�c��٦`��O���R.Z��D�E&ޖ�6�:�%��͜��1�_6)�n[�7�A��Q����t���I�.���?�}c�.����%'�^�-U`L�.���2\ ���um�m�][��j���|I<���)����У��v�u�F>�W�){A�{�X	 M���f4	bȹ�����v�'>���؍�� >k6�w>d�H5ǚ���z`̪�LR�[�uSyyy{�x>t6� ��4��tE����[u��х�,uEbm���D���а���.�I�y��iruz\*t���[gee]3<�����fg�X�����Ii�ZqS�P���O<���A䵁]F���lN���dm�V��1�����AT(� �W?���=V�̗���Lr���Y��&�3���~߫�R���]�֐'�i�f_. �L��9�1%k�����WE�)���umdWN|�!wz�C�B<F�f�4��y�ھ�~S�l9L2�J�&���Wa�RT�X+�Q2p�T��q�o<@;f�X��+�cR�C��C��" [ؗ�VF�@�)���.�h��$I�r0�*Ր�#ץ��m�I����]?�#]F���:e�2�>�G�,a������w*.�,�lVY?�yXl��I��A�r���*7��L�%����<�*JJ��:*-�2�5&��jdzU���jO����33����gö�$[i\@@DԪ�����a�zVo2�~C$P'yxhBڥ�|�e�$���g��K�z�g�xi���_ _�3�T����rg�jE�WPaT�N��%$%!G���O���J��贿�"�wK��nH$,j�W4-i�Xʋao7tS�ww����O��_n�\�~��R�=�������[~e:�Z� 
�	u�����?L<f��V�I� ��y�V�ؐl�ȥ�:r�z�J]Ʋ�?�V|h#.X�L�����*cf�@Ĝ5���z@@`��������$a�=�K��O����^d]еY%�,�!Ց��`��?�-���k�cÞ]�H�p��4Q�MM�6W����a5=Ыe���ސl&�lhmݔ��w�%[�p��u�)Ӣ��2V�H�c&�v����u��06p�����um���!���@�&�|�y�bZ���x����s�+�җ��
זoh�{��f����^�аu�n݃@�\p�/��%n�>z4}�n~h[��Ͼ�j��a'[���\�%75�Ng��юYO$�`ۏ�	��$��2�)�F� �����\Ⱥ6o���l�����Z���*Q�zSӪfn^> gt�j��5mh+�t�e��hր�rؗTu!ҳ�VX�ݺ����H�v_�C<(d����-I�z������Pb1�i�wD�w���k{���)
�HLJ�oooO�ص('p�����5������݇$CK�v���܀�`$���SO���zx�f�i��\G��Kg��*�e2���4_]�B�ބ��V �߉�xJr�Xj���1G¡��� �_ޟ6k-e�iw�?0A�1������V�<� X�27�.��,��5���^��i��{�R
�-ҳ�]��}�H\	�E���!�g$�����;R���)��E_�迄5��oJc�ϖ� gJjA6T4e�����wU��n�Og��ʾ��8
H.�k�%�Tx���������{i�_}\[PSG.8�ibe"1�2�f�L%��A����`)H��%T1H�S�1�!� �(�$r��J����#��B`����n��I���y�Ӟ������'��u/X�k�jbgQHA�/{�;�����?k��·kt��GQte��b�o�j��u���m���h��p�J�.ݰF7�n�=�+Dt-,z�����Գ�Q��ϋ��<B�M�'��0��t�9Y�[�' �F���r�ɿ=��V�����~¥B�r��"u��6����%�p���x�4[�0Mۄ����F�7����B�_��G�dx!���īZG&l�A>(�5�DB��� 0t?�\�ݬ�e�_c�' "�� ��f�B�;]L���ڜ!gr���9�]{j�R_8qHHHD&L�!��FV0lf��G��ܸ+P�)E������nvE/�w�v�f+?Y�9�Qs�$O�|8�i�Qx�m,�U�����ϗ%�;�������@����N'�Sͪ��&㈮z��7�	�?�S/��1��_L�4�|�L�:%���'�ʇ�m����������$�l�\��D���.)|Mܠ��C���َw �{�y���h@��'�ۯ,KV�W�ZW�������xR��~�1���� ��2`Z%@�kX��Sخ	�V�P	���:�޾�}w��9�ьA���Bp��	Ϧ ���Qg	�KsZ��T�\�V$�-����nQ�~,&wF�rJӻ�p�䋐ƐK��Xn�k>=k���7�UGWvT��{�3��BT�*'��}�؅�Sw�߽$>_�o7����������8b%ؽ��>�][]�z���2� Tu(
\ݖb�tZ�ݾx}Y���x�T��K��V'Gmu�@ݥ�{�Auʹ�_�<�3�9�!��p�a�t�V�)v~��W�������[u�C���[�T���j���!��NA��կ�>�w��Ĳe2{���Fظ���c���PP�����k�+�܃m����C_�7�a��v�Zss�;U[��N��S�)����`���HR#0S��;Qv��U��of��C�f�jS��q[o�3W�Z�O�A{��y0lPA�q���j�����9��ּ����Tl�`�GMx3)�"�	�L���DՆ�3�7��^�n	<�CUF��Ff����G��-�w�`A�Y� ���*�D�y6d�N?й6O�T�g���\�o?�QbS����.V@����Z�o>�����<z�ǣ��fs�Q�e��lAϗyr�F"-p�qUTA�T�;z6��!+��^E�٥"�U�x�	mIq� i��Is����.~��Ħ��`)��u���'d�d�H�|�git�Fbh���"��t�?���b`�	�A!��5�~Ĩx��|���f�L�Υ@%���P�aq�D�0�=eB���2���8������QSc����d��b'W=d�Z��x"#�y5���PK   t~�X�|�	  	  /   images/e1d4e862-170d-4bac-8b1a-e4319ef50e6b.png	���PNG

   IHDR   d   "   ��|%   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��h���O���&���1�T��]W6�GeJS
ҹtD���m�f���]�1��R�,�9FAA+���֊�2��DI)�6m�1�5���������\�{����������s��<��y�s��4�ڵ��X,�V�X�***����U�7ܗ���<===}�֭[���4�IN�:��;IH:333.�T��l��EȬ�W�7ܗ��Yk��ּ����_Zh��Ζ��.L�B��fw#&d�t��������ķ��������q]����^8::Z%O�r��/��Ύ�q�[!��l{Y���Oݽ{w������nrr҉��۷o�&b��P.�xo�	"#<55���R/�}D$<'w�f/���)���/w����ϋ�Ú�#"�$�|�r�E�{��D��i�ؗ PT=��g��Od�ח-[�B
��v��QWW�m�"����P�c bD�a��Aqq"�/_!Me���DU������92)�E �b���3c{�{M���������P@�I�ɧ��J�$�Ab8�%]џ����ا��ғb&�u`��[��=I��E�2��8���6����K�%��=)9)�O�(s�\���>3y�Br�����2dr�w%�}mOH�,i�8���6����ԥ���\�'#������v#����F����3A���Tz��;���w�� ΃�876;�ֆm��I#\�4AEZ���<#�Νs;v�0�ޕ����ܽ-�Smȥ�J)��댓LkF�|`|�{[������\��d�o�T�CaD��{��}�H5[&���l�g�u���C�n��k�p�Q[5 �H��Q�w6v5<<�A�3*޳r�JW[[�jjj����s�@w�`�8��N��  �W�Z�}'#�?���\��ې	�T� �!9m$m�,���\�~}�ڵ�7Ƴ����_�gƓ8Dp������,��񻾾�555y�GX�����իW��h�����h�s�6x�ӏq�TV�\�J��!Ni�>�㥀+��%���U/�Ѐ��xU�'oi�9�g���LoF9�}}}��͛nӦMn۶m��ٳnpp�ف��Q����x)��[��ׯ{Ě���]��l�3�ׯ����d�|Υ���2C����;/ٲI����N@�.9"�$g�ʋ�R�]F�\
�h�L��JXB/����������$���XhCCCNi�^���$�Hd�
��� ��9ق6R���2'��e��t�Nc�#B� [NI�@�E���O��P#�-Ƽ��,�e�w���$�����®?�;4��f�o=���b�A����	[�a>[��E�2~I��YW P��Y_X��I�a�n�rq���
^^u��8k�2�S���+W�T'�6\1�
SdX9�n�800���9� ����*^:���B��7%�K�%i�fF�b����AW"Fe��G��n���8��&�@��:�gN���%���IK.��8�l߾���	wX��o���I�����EI�ZEI�J���^�ڭ]��[L1]�׳7��u��Ϊ(�@�ӭ_�>���@�=��/h����)df$�.~��?��p�����k�yCA��@������7^�q=B02��#��Bi�B�a#d\�l�<�3��Ȕ�T��C�R@?�q�C��8x��L��aez�:;;�� �&7�� ��ԟws��u��ǣ�����?n,Bh�9h��Pz���*�;v�X�z�\��b�V���#D�3�Ȑ�>r?7!��u�t�hkD������	9z����ݻw��+"8�<��8#p�ԕ��4�`6���A6j�:�Y�~j�$�{E���]!(��}��yJɰ�sV�d#[�bD��#s���W��K�X��f5��� _��hߺu�wV
"�r�Ν;��w�?�x[��UL?�Lo�SO�e�h���/o�Mm�DyUu��>��[ѨwvR�p��?~���xe4�>t��ok'&�1�g��~�Ns��5SS�YoSM�W"�*x���C����EÞ=��{���������������������������n��K}6�xT����?�&'?z���3��ӧO�{����>�ש�=)+�\����W{{�'��{V����}_R�X�YB�X"�ȰDH�a��"�!E�%B������#�    IEND�B`�PK   qyX5��<O  g  /   images/e63eccd2-2ed2-47c9-a1d8-30adbe2258b3.png�x	8�m��P!B�a�0ƾck�l��Nf�1ƈ��O����:�}�,3���'"#K��NQ�o=�|��������������w�׹]�u�w2�ڌ�[��D�-��8��ᄧxh�0��	��H�ۙ�Q�do���Lup�9� �������S�@)5���MwT�]�(vdD�?�\�	��]��u��K[���mT�
+G�yK}��*��~,�[��>�_�5��R��-]�[�Gգ�/Q�y���_��{>6�;g^bɾU�J���P���H��d+��Vfɮi�JÌ�x�>�?�UPUo*!>'�Y;]ʓt�m�ġ3�-b㺔�Ur��c���sX���^ς�cR	�'�&�q��M����_M�m�<`�S�|g�?N���	�V�{l�Z}.,���t�*�O��8���!;����EyZ��w�	")�~x|83纀ǵw����摧+�9˛
�h)Gbf4�'�I�Z3�����/r[C��k�.-��~�����2p�d��43����G~�x~r-:�@�󧨏�	�P��EY7⅟�'��65Z��ت~wj��C�bS�Jiw�0�I7R��n�}�Z}R"��Q������pT�^N�aBX��l_t�FD]Ь�#���v�c7�����w	`�r������q�
U	Jq��-*>�Do	^w�uk��[�^��{�U'�M�?/R#��J��[�bŅ�^�1�Z�G��w�Q5_�~N���g��~�F;�1x��䌞����jv�9&#:u�Գ�j��*���;�o�qk���^}����-}�P�#��o��f���)|�-���X������gs~�A�b$�I���[/�_H,�[���o��~k�����Y�ϴ2kφ�7�C֩�ʕ���:�&��c?ښ^GwD���nuc��ۙ7��^)@*Ƚm�wY�u,R$�`=�S&���i?aI�����m=T���qy���Y5�)R �GH�yIM�l�nVrdKެf_��rp@
�q\l��l$xY���M��C��ې�);�~{]{���>#����*�}�D����k4���-����p�Eo���}M��l�Ǥ҃_Y^�Od�\��̏�\]�Qm��(��n�{�l�8��4q��y8���;8G�h/'0k�[%�����[�[k�P��������hMK7�el���7ܮ �Sc٨Q=��.ubo�I� �Gp�fe������g+K����%{��H��K� ,�Ë���=qx�?2��������U�	��dD �>��A���B��zap@ 	G� ������a�O�p�}���B(D�h�v�B�O�q`-%����2XKG�S�[����VUVU����T4��*pU������z�퐦�fz�� ��BCC�BՔȁx����LY��
Рp�G�?H��$.�+�@!���;}Or0��K!x��\��_�|���T��a���0�����¿G�y���7. 8��IX/�G��S� ���� 2��C�oD���WM����.$��� �I�?����8�.��3	Ԕ��w�?A&₂ W# *������ 6/s
.@P<(?!�� 6�@�/��q;3����	���7�Q�0��3� �築T������,m���'q��2�+�jPU5��\C�����WV�jE����-T���OP������z��Ɂ$������!�8ΏLHQ�G�9�����# �� �S++�����g�D@ ������izzji�@�pZZPuu�T�ӄj�p���**j��G���w���x��p<?��x��������N�(���_K�w�כ�35�^eI�G�E$����k|���?��/Xٛ��3�6�.q�����)���Yyx�w(��������
�� s`�e�_���K��M��O��t�.�8@t P���Z���̑F�0��<�$��C/e�I������q���H`J9]vYX�r�b'��{v�]A�F�$K���vr���1��<@��loM?��@�����������⑻�6_lq}#�>Z�9�ݴ��`�V	N�Ɉ�O��G5m~it��!�H���mL\

y�F�5bmE�~l�q*%m���ɤ���y��+�Z7�Lo��:�8X�5���E�rA_1��ML�[�u���9��o����¶�Qff�);���=�F�u����t��.��2L9�����G��=>}}+B�aqt�}	�6���7�b����g����Gغ�O3���7C�嶷���WҮnWK�Q�a�_�EO��.�o�i�&V�b���617�=}�������fi��u�{��o�,���0�{������(?	_}��ڻ��E6��v`�����������?�WV�����l�i�؆�>���+�-���{u�%�)���PuJ�$w;"�#�2�S8��������(�Z�@L�.8o�����o�*����ϯ�'�\@����{=Ș8ܷ��7��-�%��+����e8N�=rfZm���X9�uƥd*	��5���g���r��A�?��~l��$x�w��}&�����6��>W�zw��C,W�-TTWy��v92cw��;d����h����`�l����.x�J�)�ą���{e��(�H�MO����[��� �����99:�[���Gx�x,�y������ثu<2u#ꢧ�ԏu �I�\���|�&6&�&����ۧϿ{ZY��.�װ2��#�ĩ�Ds[y�6#�UO�G�v�t����{�y�h�BM*[W/�R(�x �p��K�w�
�h��Qh{{M��ZX6���]W+>W�s�[Y��5�	F�Nf?֜!���vk��F�_�̬��j��gU����
�Ǉ%+<<��EQ�i�M��b6>�L���zf�J-�����.#�j�_�ē��j�H��cIl´��d��Ne�H
��0�n-�������p��8Ց�!�E�WK��Ns�Wg�X�����DҔPHh���Ř7�l�2��`�L�K�L֍�2ѝ"�5t��6�X��(w��c��{���]B:$sY,OU�j�]^���3y��8��:Qa�&f��7�3ya��
ZV��t��I�aw�,������C/"Jrh$O��i-�M�[ �sZ����;�%rt^ߢ/g�hȯ��P����1h�#*RI���h��n�Eq�mE�]���q� �p�-:���i��ET�5�}��2��r�:��COm"���v����'-��4���yQ1���JR�a�!�L.�sֽ�/Q�%:�6����X���5�|M�J�c��8����J�W�+9�^ɹ�B�-���h�H���HΥ�����y�K4�)SR����OR2�G�:�H��W��)�={֓v�2y!.���b�s�Z���������jz�BVإi_�)"�`h[�^�]�ɮG��Lh���4nꚞ@�'I�Y���Ǵ�w���<���r�#���󹤆&�(�L.�vE ��1�H�k��#04��_���z�dJv?B��j��%�{�����8��v78���⨮fm2m5����<����s<;��l!so�`�\`���K�Nz�q�f<I��	���[Q�c�F�m��@�GoY��'k��R'�u�h	�i�(]|?[Yux��M�SE��]��3�\	����d�Cb`�(�G�����yRv�|��|���X��0@i��o]0V� �=�hw:�E�B�C ���V�Ёt�p.˰�� _�e�i1�_-k�S2q&�o�1��tD�r�9����1`�H�/��_0Yc�ka������M�Gm!�ed���tZ'����`�DQq�����n�L�+U ��)d3Ʈ����B Q�5ya�!�F������v��Bg0$C��/�0�r�C�)Oi���`t��bݫCϞ������<I=(C�NUb�9|%�T��
f��9��MZ>���[�"�4��"{��/�b >ጅjGL�һ�,�Y�$D��[�z���|�B�x�,O$F�UӏE��A�"3�+��Lӯ9:E�V*����Є6ߛ4��.�ٌ�rE�C�yz�М��!�ʁ��Y��D�T,&ϸe�q�׿���
H�����@~5ٕ����T֮�G�lU�`�<C�W��tm����V��ɪ}�#�3�hҺ*&T�m��e�V�1
S -T9�ϗa�;M���W5x%�@uFʬ�K5};���~�N�(M�ƥ[�>ټ]w��Zʗ�0�gw��sq`n�t2Ӥ��Ͼ�,#��ԓ���nQ�С��{���
��(u�@�d�!Q��ߦܙ��=gS���z@R�޲�����KjM8�0X@?�<	��;��)�r����j.k���y�Ȳz�/���?^�&U�Z���e|��/�7���0Ԁ-2m���}��*�XS��Ih9s��<H�F��'y�E��ߦI�p�P�CA�l����q�Iwq�^Mʙ ��a�+���5�"�KI�����ѻK5��br��M���&U��y�����Pp�F��|��ٟ�qɐ���q�C�I���D�� �a�ާ���TdD�˩�om:�I���s5f�u�����S�{��I�G�œU�D��b6�#}�Vv(���R˄G�b�#���O&''��L]�||��}'�8&�d�����r���I('��mkÑ���O7�\�-l߅�_��j,�?�1<�FI�o:h�>z��b	5_7Tihd$���3��ɰWv�%̮̭{WK�2Tf�!}���]"9��98�Ԙ�ö��o���ų�۲	��� ��/�y"��f�狥�?����p#Ѷ��.y�>>����?���ߵf+�1��)mؿ0�б'0�z���O��M�R��D�ǥ�hE��G��i�"6�Vk��RRInr��,є5-8�[3����;'�2��M☐�p�F���^�A>q�J�a̙K��U��\(̣�?�>�}~��0�����{}D�xaěw�'��s�P?�|k��h�K��&��B�]�d�ƈ<d����,�`Ij�xe;5e�����w �$.��?�'�}��:�]#a������P�Fq��Pn��6	�%���fw)�<4GM�Pl��а��q����P��Ư��/�� ����b�}�B4-o�@����M��N�G	�[+C�W�'���w�Z�,ߒ�O ��_�}>(����¤�;�sGlOo�Ŏ��,-�Y4�/�"�3fa��b����%���,�՚�!㦓��b��c,o��۩��f�.�+9B���H��J����b!�מx﯎N��[��ix���r��y_����Sk����GIm�[wt܍���`o���L&9�yґ��*����n��'$�?�I�i`�T�#��j�j�5)o*)/�h.h�H|�?����}%��qd{ f�,����E����f����om6��ρh����>�G��v-܊hc��8L�&_�2~��-���u�5Ht�LZ�
x&��L:(�}r�HXJ��>�*�ez��ο�"�������wl�7���$��e�]��bb��bF��uG,|&�ag�X��C�5����wH��vH�,�;�w���ZCy̨����|�㓎U����%r�j��T]_�J�U�|s&r����	ZJ����[��7F�a�jw��W��1�����8׻�~V��GO��Xs�Yǌ�}�V�ߒe����� .�~��dm�q��j���C�CufM�<C���s��}��j9������u{����E6�3�G��m�w�BTz��6>�_޽6�c��P�Hw�.�9#kR��/���9�B�2C�_��R�|6b��j������x�8�Ն��B;���)�}�o;/ږ��zA�4r�e�c�zA��=^���H�c�z���K�@�.��Vy�5�`���F(��Ċ�d��/m,����=f��_`�6��z������ҍE�ݬNf"�������b��ɘn��w�����:c�i}�4�\h��h��vp�qf��V��X�������]�G@����q)�������e��9&�Z-�rLxC�����k�&Ә�5x�t�~�'>���j���-ᯉg�bI���}'��K4�r
��˦�$�������Ys]�m����0�y��%o�h��LMMM�-��=�R��k�}(���Sf�R�JϳU�4-Ϝi"�t�7D�Ϗ�O^}'UG���F��\?��%��?\3������h-}t0�dʈb{�j��tpuCC�jfwy���י����1�*q�ej�2K-#�Z���x����8;�ݰ��q��fＢl�L/�P	�j����l*�Gf�`t#������qp<� ����E�<�zg�Bk��[܃�?��&��{�g��?PK   yXO4��~� � /   images/ece94f61-988d-4529-a2db-f0bc9c1368d4.png��[\����;���@qw��b�݂;w+Np���&h�h�w-��-��w_{����Z׬�����]m| ����>ʻ�㿗�m��.d}y��ړ�49-��P�5�9���������'�k����!����!�a�o+�h�w&��c�v6X5��U8����>���A&�l�p�a9�3��U|-�g2��>!�#���*�G$���ާEկ[��닃k�'�s
�w%VF[�g���N�\�s㨣�����1t/�Z���g��[�sT���GN�[���:����E����P{��cY$�@�N��=ݯ�^rw���K���MG�.iHš���e{��� ������ױ��J��$�tt|�%p#����8�m���Obɰ^�8��Y���<st����r�����8����_*��up9���wi��@�Ui��a� ���AT�Z���x�Pj��D#L���J́ܣ�������п�}���nrf�)�W�%wV��Ftp�u:�������O��-qM���9Ŀ���������M/QT�!#
�A�>t+�IN"R��o�9��v��S5b�����p���A<���W唕?��m���3��S���N�p��@	�W��?�Lc�jjn�6dv���p������/.��N�.�-G�O:��M������UH���-׷R<�ѝ�A�k�M��-�r�	��գ��Ф���y���\�Y����s&�e����[C1v�Jܷ	�����ĲO�.̤0ᴾ|�C���]����ҋ]~y-pz&QugU�)�YB���\�$pkK�~�g�h!J���'w,�F�`�$�)oʩ9 ���ngOV�A��ʉ0����h�?N��o����� PI��DۧdJ���F���Icn��A�=�׬�D�]���n�\ݩX�YIX���AdZ����,��+���H;7���]�A���&*j���y��H�������]�J�z�(9���W�|{�YRĺ7v�M�y�	�FkղV��HuSrv��W�znci,��N@&�N�+hՁb�p��z�v��u�G�Ǉ��O|"Q�rnR��8�ip��NWC,E	�◦�mj�R���EltQ��7M�&���Xk2�y˵��[�W�Jg�]��}���ǹ��k��D�����L�w.��aܫ	G�����3�2#w��M:z~gj�����,O����S W�Zi�ǘuU�w �3߽-��h�>}qʋǈ/k�$gX6O �C�����Y�[�/(.�v^2д~@�>��������m��-..:+RjuB&���%g�m1/}�(|�X��Z3X9��_��%;2�>�;p�7��9Ys
��sq �G\HU��6��7I�et��rr��>�>���ů��!�����o��ݤ~��ڊ�´۹�)��SP� 6nS@>��,��/z6�?��ӱ���~�H��N��E6=�����;/ �(���_a}ee�!Ue�� 1�ly<Hu�V�|�!'a5svr"��-����8N���E_�q]V#)����r�م�zz�cC��f�v&(ó�"4Ar;���˚q�l�FKs�4��M����OJp��1�@5f΂Kύ@�8/:z�����[��ʁg�.�VE���hyҵ�3'���U��������5�0�+Ƀ@��4�2"�u�6-�?�r�Q�IګDˋ�M�� �,��O���n>u��iD��r<�y�	rd�dHqTo�Н�ϓ�:2�=&��9�B�S3��� �p^x̂��#E��7�!���X@��C�4eU.�8U2�BH�P��|�� ��	�9�����DG�i���1����ã9���jY��r��=fw��4DߛQ�;��sHT�Cd�X�{��?da�KR���3]��k}�,H� .��q��g8H�T� No.D��7�A\N��2e~��[�٣���|�����c&`\ZdH(�B��]ǣR���q)t����*CE����W��#��%���Irvz�k�߲}:]Ę`k���|�XZ=�-(h�ןӽ��❠�m���_�uM
 ��)�UPpo�'��:�҂�_��p��8 c(mH��<��?
�V	#��J�Ǽ�/�"������tT@k��J��>ol��>\�B��(p�Q+}����;;�%驩��{0䩑����n���y���G�E̓/���~j����s(���	�hNAB'�R�λ��E� ���+g��<z�����
3.ơ����AOE&�x�>=`���r���{��+&ylԗ��7����GPo��e��X
)x�Q�UD4��[�@AN��t�A��ıy8�`���7k�k�g����uo��;�i�������+�z�$`��D>iK���A�������5]a�ߜ���3�3�gC�D��̏MS�d_9$����*����d�t���D�/���ѢW�_T���'~�Y��5�C����C�&�B�	��C̹ !Bח���o� W���c��JY,%*�L���X*�U��a7q�}f�=;�p&x��'�Gf�,��Hr��W%�t�3
 ��Б�r,���D�ե�Y�*2LR3/�<ݵ�n��iOX���cx�W�_`��Ey��A瑻n�ލ�|j!BW�qsU�_p���1��>a�����[4��0IXǶ���@_���0G�>������67�
f�.��:�\����ƈ�����:�dΩÈ
�OI�Z&$/cX���n�vn��Je������k.���S_%剑Pݰ��
ǫ�<��k�j���<���b�Ť�%L&i픝��	u �?�� �0x&�����1�uv��bgߌ�kJ^U��0j,���8_�4��s}(g
S����H��F�76��D��'�7%}���W���v���������z�����cJ�}��".�K��I�'g��}�c��s,�_2�}О v0�^�ߋ-�Zvy���q��!�X��q���{���&3X�V!l���朣JDZ��&�R���P��[=�C�[~�tFL���^6.:�t�ϟ}ݜ��N@�_X2gf�!?�pwAv���Z��΋�+�������N-�i���q6���"�d"��
GOՔ˷y�,�u2<��7�-�D=A�bI^��9��X���g��T:�wn�fS%���H����lOT�Y��j*�L����rn{s�0�G\j�Ze\ƚ"��a�!�cY�4��'_NH-�h����D�퍾��E*�O1\7�TT�ٱ�[�hͼ���Z����	��`�6�)=�u$�wH�%��ʐ9���"a����c�x��<�;�����A�X��e�l�e�Hz8X�j�pv��ǫ0�\#����d� Q�o�i����Y�A ��E����1�+�;V�]�=9�&h7�e��u�CN#l[WQ/0[��K)��i�'*�p��}��b�4{�驱����@��7��� �T��ؕ:q�5�?��U ����wL����S��%(7,O�B�c$�d/o!y�>%b��ROY�S�,���bJ�~BW�>��W�IdP�(�J��-sG�	[iɍ�BS��>Z���^�xn�4>$*M�gWy ���p�Z�e&<'��N7�2v�Y���������E�l���aZ{bX�iOW<!>�8.dnͨ9�������� �1���K:���>X�[��Э�E�XQ��������_ ]�oF�������KBAE��B��Bw�����s��Go�~�5���b!މZd�y2�9<�c��эzZ
��=�Kr�_���X�E�U��^>#�|O� ����؛<�2�Qbʽg�W�0Y(�����YpQ��YJ�\�d#Dr���[(�n%�VQ��Ċ9ͬ���� ��86d����絒���S� � /�?
-�T���a�w�?��'!*r���=�tF�������J>>�ce���Z��1�����	&��Z���`�"���ߘ��sq�S���1-�fy^����.nQ�G��m�`��dc�,�q�-���P}�04�8��|�;ӡ���?��a��S���ψN$a9�̄��[9��j7b�9�'�J�x����t��[�B�,xtK����A��=�!>�Dd�=����a�}��c��7	M0�@CZ� 5o&� Å��JR	��i\�pR����Z�e��$=TҶ\b4$�J�`���3
J��m�m��참(��a�r	�$��_S��W��e����H��emE��i�-��*�r�@zz��m�ʹ��h��II�g춠m���ź�D�K!m�XD����<�n��(�'O��m���^~G8�;��k�%JE������ooc��£$u���z�F�ʪ^��ޱ5�o%�q�������)��|��3$e$ۈ��h�#f��œ�0޷ Q���t"���b˩w�����7�q	��9u���+����|Q��O-čN��G�۲;���g�}��t�04��r�B%,W�6�]i�/�4[B���a�.s�Gw�q�-�m��r��;�\Y�JF~���A�S|��b�X(�%Ȃ��*�^~��Zr1�pM��>�2���~./`�z"���O�+�ԭ��5M�֠��J�����JA Q4\���2)��S����<e*FS�� DR���).ȶ���	akr�& :LxA%e'�_1׷��T;D�c��1�%�S����~�I���u,!JBg��ʢ��ib���+��ʐ�|�������<V�K�E!UeJ���)gW.�z
�po�'��Y<v���i�,E0��SY�N���'�Ɏ��=*�\k�Q �z
\}��a=�Zo�Z���_d��7����f����XdA�f'��^�8���Ӝ�g |N#�<q˳?�����h�9Z�b�	Q����V� s2��a�3)����)� �����~�7HE$=���_J�t{ -v�^[:zߟ{��+�0��)%|�:����ˇ��p�����w��[Ux���ˀ��W֕<A'W-6�&�ѷ?���]0���H�W�e��e|��o��W�cF�Y�fk�2~l�(�\@1m���_3�:o�8ƨm�)6o��"W���^
�B�t���h�db|L���}�E���(�A�̪
u��uH��fDf3b�3���#$�|�8,�竍��
f`�r��Bk��� 	�ʐ��* \#� ����I�2��%��,mḱ)H*|ԛ�dNRȕ�8��o�L��lZ�:*�n�n9�<_*h���Fȑ;��Sl�K�FA���ɰ�qH�H&Nc���M��m/�;)��+V���+��8���E�	KTjG�5zH��H.6�rBr��mc
��A!�9`�}�,�#D�/7���a��'7��>�*��S��+!Z&�җ���W|H��Ʈb���0g'��%.��H�0Խn�!@r"�����Ij{c������2���4!*S9�**1��`"-��NE��V)�8�X۠���1赤��|�8	�@�\\�IoOb��YE�S��K�ho��u�<}�(���`cJo%��C���=%�^#y���(-q!k�z䅴��Y���~Ｌ��Q��J$I�yL�O���U���� Y�t��q1�����we:1�A~ � �&������z�����D�ءHQ���O��Z&}7��X�8xK��1�S�d��I��t��т���a���J{W�#�!;�4w���'Ϩ���}��p�D�"�%@rxX�MC��
T��<�Iz���|�}��ODNy�K��J�-!�G��R��P�@����ؕmK..嬄U���h�S��E�\7����F5�7�Ȩ,�������/m��@E�i�=�ެHmh�������6�лF�
"�g�b�.K�#N��%�i�+�k�&�f�l=4���@,G&�Id�3�k"RS�_b�Wi����p���$˪�R��õ`�Ñ��3�5��AO[�L�)��Y�(�3eЊqd�ʩ�	{�2����aZ�g���i�(���!���Zj� m�K`��JCJ��s9
�Tb�H��H1	�]�8}�|Bڍ�,��`"x���Ĳ�nGP\L�Ҙ���ʒ���Ԇx�����#�H��}$�B ��tT˧VX��`�B��?/1 ��R��qѼ�^��T���ԾHB�z����L�9x�b��<ߪ�R�^�3�m�]�O�YPR�=N�#�+��(��9U�C���N�[P�3"}�0�����~JXGN�m���Ǯyo�n_i�2�gy�EdV�g`<�k�a�(���+/�J&��fj	��s�Ag����\W�,ָ�"8���N2��xj5���*СXE���Z�����U@��i��A�O�\��Ѳ�e��"t��Ce��>�M�/�#��$˥��\t�|?��}�Q���Q:y�"�}�L�k��BΔ���-bִ��i	<��Y�8�I�]O��"V�.#�IE�hNF��_���˛�M��y:�z��"�m��?��<ļ�Ė�QN�.���Pl�Xw����Vu�E�#_���Sc�
E<�-�������8\�M�iԨ~���Q.���W��c���l�̘<a��3c�)L�}�豱���vj:�]���m��9��g�^�C��Ba�;��� Ʌ����a�4a7�۟�Fl��R3�?�}`�YlS	�l9�_w�5T�8*&��{O`"\(양|c�k��S2b*��M��Xy Y���+ϛ�T�<Sl��#����&5E�:�"�x����j�#Ɍ���������,�9 �n�.�]�Y�8����6�O�ٔ
��`o͋�jd)fN@'�2KdV2  ��{Z�`�t�s]������4t���K�sX�vlhNE�7v٘�83�x4��,�����-�,c!��Q=�a���L"F�_���">�[/zcȽI3?�ᱦ,��ɮF�*3;~�jA���IP9�!�ԃ���v����A����.��9VW���uT�����o&�|f�=�r��{˪lO�+��J(�w�8P��~Y�v����3�d��6�#ޚ�U��Bt�ax"��_�K��CǄN�]+ˑ[t˲�$ˋt��E��x�zO�ld�.��Fp<�4�l��J7�ԠF�D[��1�]�3h�%�#"���Q��$�uD��y�䵳p�a��"�e
���1�:V<Msk*�/}D�Ȇ�W��.!�=m����$�C�0ؗ�G��P1�y�$�����\�-2F�z`�Ͳ5���j����!��p!�`�Ut]��O�Di���#t��1���/�#�!$v=S�3��ޜ�-L���_"���\���b'�)=#����J������9��@:�R8�{�CEW\�U<Zasʕ
|�r4[��X�d������'#N��)j�I��_.������n��O�� \�v��*�5/��lО?�
0��
�TY:�|wxN V]����}2�A8'�5��K����]>!l��i�i�� �q�$P�쁤LDC���^�r�A�#Yaj�����
'�PV8�7��3|�1v_"��O���K��5yVa�Eҡ�� +�?yJl��0d|A˩p�c1���8�9�49�p��oϩ;,�-kp�PQ�sOG�)i�b���>]����Y����'��&~E��en����a^�y�ǲ��s*j1/Dה����	�T�;�霿(t�eS�U��:�c������$]���s͞��%�ɷ9R�ynk� ���Y�S���c;��!&p���4O?�&��Μ�fW��-�+mF�l�Q`�`�����qވ�����3��,:���orKu��k�Z l7�E��Vy̟�|�ޭ����6���7c3Q۴gUc�]���)��C���w�q��۩��͖X4��1�j7�2�
EPY~D�1�W���T�+�B�4�07�e�+&��D r�#�$ �C=�g����ThE�ՉXe�9d~m̶���\��ӭ�a�e$�g���r�̲}�A�r�?�r`(<��7�9�Bʎ����8�
�~~j��'��D�)��#Q��4���M���ey��s���7��U�"�é��i��8:�`���>��Q�t,��{�6)���A=:bW�z�뇠�v��;����tօ�h�	R�0dx��U��`#�i'{����R^&��-�����H�8+]�Yo<r�j&�V��RE�b=I��Mg��5�?���
ĸ轗���x�H�Z]��B�pS�&�+A ~b.(�g���*���ej��������L�)P�pz��>�R�=�S�T�a�|����9P1N��1(<��ҕ��ی I�,2�YeT�ݶ;%gX���A� �ʪƤT P����!F��b	�z�����9W��P�u�����u?ښ��*P�{Nf�]�� %oj��8�B��XI�b���7z�A;�U��Ҕ�"���,���TWmg�u��݉ѝ��{���ն�)ܳN�EMh�y����'�2h�
p7p�(�IJ.F��	{���S#�v;����ߘ+�?宽P�R��*�s�bP�$��W���q�7FS���f��ps˭�Y�q�t�������D�!�ӽ�N�_f�kf0�6cQn8����L��xm/��[\m��ňՂX���2m	;�nF����.���*'\��V1��͑�jr�Z��P�6"*�l�aߌ@����O�L��p�o�J�,^��b	~�����a<�	0p7g��$��j6���5[�G���D���q1{���zhޑ�KQQ�ZK��?�{�{L���c���uxO��nI�����:�~-�=�"S��@��]p��J- �?�P�i��H�ˋ�n�E�O���C"Ö#y��HR��{e���) ͋�]=���'�N�/+� �;�&Q�1v,�S�v���G*|9���#��r+��g�Pve�&�.z�6]S*�����>C�t�V��i����P��M�x��P?�h-��_�i�3k��w��	5�x��n=	��Ui��L7�-@}jx�D/fD�U׼���4o�D�+k��!�����*�����	K)~��6)�SB�i�3=v�k'�#[��TH1(h�sr���2K��1̯Z@e��T7��d[�t���S��&�=0�ډ�,�5S���v,84�~Z�bA~`��Ix�6�=r;C�sR�/����-��o0��a���ҕ�Un���>B1��E��Ӣ�.��W�(�EȫX��g��a�A���*�K|�v�S�>�� 
s�:�k!����Z��F��O�� u�#��#/se��Gj��J�kN���ᬏ\'
�5�{�o��0	�&\��O��Y�\ı�÷pL�4�tj��+\� *l,0ؙ�a�*�|-�g���t���"�1?�U*!{ꦢԭ�S�'I-�B��oa�����u�ڿÂv�%n쮝i3IY�o|*��(��x�x�s���L��o��='��
�%R��	�1_��ð[0�?�Y/�_���+0}����8�-�Fߡ��1�P	������o�#`=Lgu`/�����.���䦅��L1d�������ny�{���z߭������A�<[O���9Ζ��A��?Е���o��U|T#T��nڻk�
�Ӗ�;�ܫAQ�k���L|)�����9���ຂ��e+����^���,h$V����������Eý쮖�V9�%J*X(y����'�5x��^*�×���o��y�9�==�����
4�{�xd�V�\�K�}���Ax�\WXD�Rm�d�NU�r���	
�ގ�b�u�L�9t�IT_�E�-�E�7Q-J/f�Qi��ڪPp�A�Z�1�G5�5�*�ҡ#Q}i"��~9qc�۶*��5"T.L��l*Nw���NQ�?���UX �bn��D�S��|�����\�����@���j�G������I��R�U�9��%E�� Ē�
|?�yU;�K�������AQ�L�=�C�@��g��ѧy�H �R�Б��|@�<�B��5ߏH���������)�V\V�ꡟ�$��Dr��.�FX*c���)ÌG~��U��Ė'�\�!	lި6W����A����f�n��'�ϣ5�	ۭ~��V��!��䗱O�'�:�i X>��q274���A�
��C��`����� aG�"�z}�F
��(zkm���1�Z��{#�����u�I�yR�doW�۷W'�0xt⽼q?U��}s��c���{�/�Oę�����N�����I�`9�Yv�X#�����ګ�U�$��$�K�2�>�1��r^�Xs,�k�nT�Nm]�V��2TX.�2��f�:G�E�ih齷6��eV�u�3M�Ū�e����Hd&�;Yp@d�_#)6K̔�_�����LC�|[ �D���$�9�(����u�h�M-&�O��I�&_�E�-d�O��6�K��;;``��n�����sJ	�5�޳F����?y����k,u���e���2iLݫ�����XRT���������Y�J&QA�tl�"W-�S�]���eTօ��'V:d��\HVI�
#.J3�L.�h#������祐BF5%��t����	ci6���^?Ie�4��؆f�ߋ�� �A��oR����qG#����d�iP�lAuV<F�ا�	G�M��wƍ�W7=ɀ����c�d֥���=�7W��ې�3��[M����ky�"�\9d�ۅ�����:ח�HO�Dq�7h7:�ux$�GmOdR����Q�Y�]�⠫>��i̮�+�1�֭��}Y�
��l�웹�Bj>0й4�z�����#��ks����BJ�b���0���`�)ϊw\�6Db�(�����&�d�d<J��0���؜�a�J�LP�̍�;��V\�Iq�golUL�������q�%oOśZBw����et�����$�t��}&����5������+&�hO,�~t]���O.��G�N���'>���y-�������O��:U�`/ьn�f����������ɬ�Ґ�7��_9U(4����3
;����ٜ�Ă�!�ƌ#@��`��݀p<��ѻh�I�9�V���L���~	���(��q�l��f���������K�S'h!*d� �ǰ�N3��I��z+ �O�)�Wɘ:�96�����,�)4QVR��o�����d֑K'�k��K�֙Ӵ�Q7��2NY��?�|p����Bui���鈜_#�N��x���5����xZ)|�s���؅޼T�F=^Ylϴ�0h���r���ChZ4��@w�o��q��^\�#3��<@�5ڠ�kybA7�7՚-�b�Br�0ڪ���+���nۏ��Z`��6�-���Ȁ�x��,��\����6Ѧ�ǞmO|���)V���O�j&�-��>ǆ�#a#�\m��lc3��@T�ư�QV����x�bQ/H?�.����i,4:-֏��i=���a�W4�����>=5��ť���s����W �۴���pߧw�zR��R=�I8H��#��#�Pw��5u�J\���C�l�Dz�^1G͐�������ZY�teÓHb4 !4{M9U�?%2�����v(�� 譒��h�ŔFp�SYi�?�� ?L1=�
sk��-���{���@/|�Ƥ��{1�J(�Ӵogr��&�U�W�~�¼����]kN�Af��V���\7�Ҷ*�]�R-���Z4N�n�7zr�/{%�P6�/r����֌;r���'���H=����'l���!��+#�&��mB*h�C*C�h��g��SMac�G_[2���]n���C	'�@�%K�]�n���og���J�����%g��5*�3�2�dBxv��Q�@�z�w$��'�O���J��2ax~�g?���X��/	�Kw��I�+��)�Ô�������g���"d��������di���bO�,j-k��`N��uە�˕rY���HyϿ��r_�Qzf!?�N[ɖ	���uxҸ��T")]j�	2�h�W.�su�?|��:��FΕ�ݷU$��eSbz�t
�.�7z�u��P8%۽:�lVa�]�Z^�#���-�#P܊�y���*-?���;�R�s:f��[�D�AAKHS�ε/&a�y�0ǘV�2z��hN��zД=��������4��9�N���t��`�ͮ�������h�T��/�tCFG˦]�䮥���P���k�c��.ߔf��O�%�c٪�ߙ�?X4�}�ð�Qq@��Yg�x 4������bv��#�Ko#B\9l��8�gT�i3h�Z�8�����^�p����s����}��W�Pt�T���dF��qD
�B䤋�?]wK;���6ap�b.�'Ɏ����rYͥ�ſ-��x�2=��O���z�.>߼��s��w�c�x�{�v�zp cY��wpL�-��mx��,Q�O�K��d�2n"�8�󻶼&����w>���%πMG�7vz7����k>|�%+�˶8qDFV�ȃ��8|j��Ԡ쒬;MNk)`�fx�	N�)�ܤMe厣evT	9���,�2.�ɿ���"��&��	�ޡ1��6��k�3L�Dp�eE�h{0�y�|��5:�j�&�Mm�~��;��hZ��}�׈�Ԝ���0}��"K
�����g�{?g��j�m���~mB<�K��zd��)LalB��4���!�}|V�G��O�
c.i�?��ѹv�xx����_�o�AկH�+�G��?��D�5�@��e�Z��f��:������<.�4�ǳI%������$.��$��/�T>����Ն!��JKɍG�毒Gk��E��`Z6_L�5s��R�r��7bS���?:����������w+�-�@c6{6�.� �v��ޗ���<��>a�ѯ��/��iY�D󾇄�˗�Y�msl���]��_�q�E����NHrٝ�x_B�O�\Z}��u��iQ�~��?�F�\���{ka�A!��������J��d��C	��5e������^yk/�ѷ(�Pl��;Ȝ�Q+����7u�U��� Pإg��Q��ϋ�N`ѕ������wC��<�gX�����<ہ����d�q\UZS�!�Q��_!9�jF���i&�����C������=3�c"���s#�%�Ħ���3����j����cB,���S/#�Jh�S�x�n���?�Ldq 銏��x�'I��4�
-~��nr��s ���F�;��?���VӍK�(�𵏄�_=O��p߄gR���3��Wzʥ
�.���nSc�����`�L>#�e�Ω�����=��we-:�pۦ��u�M�a=!��ặ/<�fwu"�e�!!}�Z�ť܂>�@�|����G���G#?Oo�A	���{M/����j�j�q�����Zq�`�fhp��y�<��i4�6��P�l�YA�Nۈ�ED?�k�b��x7�E�Uܨ}a֟�_�"^�	��~Ө-�<����R��7��J�[���{4��X�vg�
]��N�G�I�6j#�ĢP�؟�^�j�VС�tR�TW��Q��T��7�n���Y�{KٕS�CPu,�
��%��ۈ"�[yTn���Ɯ\�����oK� �g����f$E�H����:uU/*�,�<Xlb$/�d�N=�X�x�z8Q&`e�6��o����!��y.C_�a���3���Z��D�X��C5��D�?��&i*���p�&�LΉڀ��Ř(��+�ҝd�R�id}�l-K���֯���[����b�
r����˒�H,�<���З'�eݭP�Kg1�*�w��~~��\F]��
5)�Ѡ���;tY�wm�{�C¿9�i�~�����s�&�X�`J?#"	�:���/w�7������x�q���km�
�'��Џ��=�������<=-�	SuB�������i1��~�W������n\=ӳH#2�u�L��(;{oԬ�!�L�'s�#�CB?`� 9�9w~t8@� 탎��XUn��:R�Ëg��{K���q!�6=�#��@��n���?j�nE�gh`����!��?߀�,Z^����Il�G��\�M���@�_�Q6�6�!x�(���N���Jā���-D�"�`�u@�N�A"[�&��d��󏸂�����`�3����`\��t�Hv=f�X����N�3���)��F��`���9O�fx�����"�FY.�T�o��KUtdؚ��M�_0��۱X 5��lqޕ���]A�(��f����*��M� �;���9��3�-4���C��ݸo��4�򁪿 _q2�_�V�eO���v������W��x��珒�&��d��m�
H�?[3���]b��?@�#jR]X�6�kzm������֔Z���{�"�U�pGt��?���C����OӳOi'5��k3��ؔ��'���&p�����C+K����y��
rȭ��;�o}m�lp�"ビ���#���j�)E�\�xu��Y�A+�Y�V���9\\�-)�O�U�ht$ֱn��P��8S��#x�i��%NV���G��m�	�[��c��m����#�Ri�%A&(����{o�~��|�[����$�|�����9y�Mk�e��SE
 ����vI��U�xB��C�;�H�zտ;�ޠg��n{�*G�}O�������'ł�p��E�	���WR���#��]��{s�g��0�����kA�����}� �p����W�Ub��:,l6x��K��%l/m�e�|�-}i��8S�m��>x(���L�4t?���߲z�>t��/������"��O%X�`��s������S�U�ܬ��\�Ԓt�)�<÷/�V[iT$�_*��~��NE���?G���@}��y�j�$ޠ±�,oA��(��2��P4����r� 1p���0?���h�9��O^�S+�-�[�Z����j���^�.	�0��{�����%�w/
pHn������waw�g���r�pa|�p�����oq�B����V�g����N�bK[�_���9�J�d��Q��ݭ�Ds!A�C��A���
0��aX�Q�������[�p7���5.���O���-�[U��ݚT��ͱ��`%ȢJ�mt�c�@i����Ύ���_�I�f��^=Tk���O��?���C���z.��(�,���C�U����!�-� a����DKm��;�2xA�8Ei	ZA��w���meXR*iƋ�$���ձ���T�/�Q���t5��j�2�E�"��SaW5�8�+�^ۇ�
//���g������}�����H�Ȣ�iHP	���qjE�C�K�}k� ��SU�*���ug
�F�e�L����nx����6;�0�"[O���[Ρ|7���O�ޕW7M�e�Y,�Y�;��(x�íw7%�S������#�v�"�<z�%d�;�I�o�_U�Gj:g!9Ģu�� ���5|6y�:{h&����D}gD����r��Y�[�_9�ҹ������{�,���Ռ��i���}|�(L��#�8�,�;{_R��t��UKg=�=�'?�$���O�X�=�&cy���L`��:��X�ڍ3yPx1	��;\7O��Ƌ�)��b,[D.~��x�|�;�A��=�g^��D�O����ՅLgm�=��«�:D"�?;@��z�j)�x�_�%^O��FOH�:&kW�S�Ŝ7t
�/��#/�f��󼎚���n$l*�.!WD(X�dSh�K�hꏝBw�F>�`h�6w<���m�H�bm<��JnO&`ې����x:W G��#�^�q��d�"����\�����zh�QZ"�G���*quA5�uBd�G�ie�e�sLw�SXv>v/R�եX�v��/ط^3s/__�X�ym�5�����6y����4Ǧ+U���oO���3�9��K��m#;���?��(<a�n�u8���x�&$~c�4�l)ǳ71�;������)Ղl3�`>�xKq��"�m������Or����8�-�d_��n�e �-�����G\�	-�Ks�6:�I�'[;�tzbr6w"z$ZW��1ZJ�K�F��|��o��a��"Ԍ�C�v�������.K7�N@�!�6 �o�. ;��`���i��/c��u}<� ��p`+�p�1N���&eQ�~NW�T]'y�������7Y;����7����yJ��uV��t

O�����*��l�R��k}�O�}�'�%�;+� RP,�W�=�n����1@ο�.(�j��k�;``���� ?5��(=s�ܙ29;]�m�Z��������/o}�[�����/x�&>�^R�~q����+9`�rmw	�~uyo����yd�6�cQЫ���"��L iK�n�*|z�r�N7�=��H��%���?�j�����b��"Vh2��Y�r7�=4z���M��#.��S���/�%�(��i:�3:�t+c��ؚL�0��g�Ex�o�p�F�.�C~���}>{a�=Z �Z�*HA���bz*^�c��+��#xqb�I�J���Ǉ�}�C�'���w�N�c[�`�'��3"s�,�d�����Ԝz�5qȖ�{FH�.�/�ce��`d^�=�'6N��6�Ș;IL)�r�a�3gN����K���߻��ȇT���N�ıS�����ܩ�⢼7(�Bǂ�s�ϔ�������Q~��>Vn��WrFs-����ó+��׀Sw@��դ�P�ϵ.��2l��C��J.��s%�u�FC;�I���vW�����YV������@�g��+�������w������m۶�~���P���;���������V����hV���a��=�sUѪ@�s���fʩ�ԫc�x������75&e�?�N\�-���/��*��(/<U^y�L9{z\F�A���ٶ��i��dШ��C"Zfd��M��%]�G����{���c?�c�G���)���u������;���|��Ry�];�G�:��2Wt�<���=�����5u�1��I�޶�7��^��0�����=����H�Co2/L�1h��[�0��e���O?�l>Y C�&14>���{��vb�0�kj.���j�r�	��c����Rݵk��1G��|"ͨL����Ϣ3��h�,��Z�+��J��{��w�x8�M� ���_
P;$N���J�����z
���#��~��=�������"����13��x�xq�L��àS��-ӓ�nfrJ=��)MB7=�<)�-�(Pk�|.�h!e��_�m�*-�+}x�4!���S��g$'�c�0�:>�.���.���(p��58w�u�OB~��������<�)�/;Gy��W�a%��`�2�C�y%��8�[f�V~+��8�ì%/���Ds�!���R�uX�o+A�_-�k��Zt^�&��Zt�+[�� x~����}w�ٟ�)���1���z�-�tT/Tטj��Y��P�Y�+��s���L\�,gNł��'O�Y�d���L�ƹ31��H.S�gΞ�d�N�,g�rbx�r�ƟQ!3�#/�xKN�sT�9�����K_�+{��-�=����A<�Q$:|�5����Õd"�,h!��6&��h���{��ޣ�j�hG�۶m��"3���k���s�m�� d� -��1�g�n��*/�tУ�Q?�l�2Z����eۖ�}�.ѷE�i?	;���u5j`��m�0���5X������ܹ��P/���{�l�5*����'F�@nV�e�i`�d�`(=�����G-<�@y����3�Gz���B �1�L�C% j���(|f���2�V$h&'lf�OZW�f����&��՜���Ey���7>��]�z���m,���N��C���s=۳�&"����C��ǔ|�o*��#o9E�G��#N:��������c�j�jI�#�ge<�C��E�Rn0��rw�}��?~�{�X��a>���:�V��
~o��7������.;���k�a����J��{�t'�+A=�+�ϰ\����Zh^�Ϋ�_��+��A�%ױ������P���X���^��T�g�t�k�,|�؈>e�h�C?�D��u�����3c��g��c'd̜*s�S����������uw���u��\*#��a�[,,B^�a�ǋ=]!�ia!\>���	݋�%��Ve0�v=s�M7�-�7�^�v9y�^��Q�0�(��G��$�Ǽ��C���w<��#:q�7o.�<���Ў�vҖ�gљt���7{��Bc�R���I��lՏt���I#y�lh�9��53�;����껻6���6��n���ܱc�:�[E��P��
��l1�/}�K��DcƔ�I�!{饗ܛ�q7-�KkE*�����*��w��#���r�m��w��򶷽�x��Q(l'���>�+���~�i�f�@�.��[&�a�˅^*P@Ѥ p5�"H��p1��;��]뒗4hpk���a)��.�_A�DY�5烬���w����=^ 8Ǚ3��(���B9�^'�n۲]=�����%��!���zk6ggh�R`�p%/8��/�᜞W��+�(\@�G���8����	o���d�ћ��ӳb32��(��Qx����]v����֜:����@.�0i+�q�� �Vr���K8\_B�r�w�զ�^�N�Z|X)l=|>��_\)�J�K��;pԟ����]�E�Z���gȨ�C�9�彪����{�Suf\u�d��I�8oF�GWU	9t��b��:"�ōenf��_��1s�;r��?{�gT���ݾu�:;��0�)���)���3fճ��i�w��V���#�f���)Fl9�J:�c�G�{T��zXk������i�Sw�n�+Fm��M9s�_N&G��ct��]W��l��?��A�Q���A7�eWkD��ݻ�<�� ��If,���е��t�	O;Gpf�@�:$���n:��a���m[��]hl���A�y�P� �gپsWa�p?�P!����Ũ��0GO����Ҩ����t
Bv�4j��0>��<���m(ػ�SǂŰA 0�0��������Y_B8h�  襑�5?�,b"�]ZQ��W�G��v2z�q+��C=�@����g������|G���>��q��GA�[�S�ϙٱ}Wٳw�pm,_|��� ��e�2�~rT��O8φ2N���3���8����PР�|Xl̷i8��%��^=W�.]����Hٲu���tP�S�D3
���,��� Mu���V�[	����W�q5i��εƻ����JP�#	</�M��*@�|�����>�_+\oވt�u�u�����P�ŗ�B�fZࡇ(?��?Qx�>Xt�g�#C�Wq҈���`�}�,֥u���S�������'|�v�f��w��*��U�uNwGS����~��]��,����	�0!}�W�[un�T_���49�:Bf0V��¦^�W�5Fmп<�fph�m���Y�1SM7-/�e��ԛ�������-bT�z�Jon�T���r�}��-C���ю�~�����Mc�8_��LMqt
:6G��� ��n��n�Y�ܨ������T�J��a���k%Y��o�.�J{���T��ZX��'�(�0�g>���	�0xh��h�7����_c0+��>��)���O�`��R6��\: �q�a� ��AH�������������Z)��� GC�r��O�JX�����F dy�|��r�����������m��g�t_��F�6{�$۫_����o���I�A�-���Z�&�8�����Q�	�\�a#n3i���i᧐UZ��P���<�l%'���I�0rp��0:�=ɱ������S*�1�@A��t��a[�u�vX�����X+���}-p%|���!��)���\g���2��%�����yH�@��z@������ҭ�';����W����� 7�����w��)��;�19_�.qR/#!*+Oǲ�M��!���޺tI�pn���l9y�l9|�U��s�S��P��tŀtg��/��.�ғ�2Z8�dQ���'��ȏ�c���:������#u~\��7��HQ�@��k�0N�W=N=r�&���g�nwVY���C�G4ƌ�]���sk����j�u-8h�͡��`0��{:�=����~a�<���n�0f��c��)*�M�?�4��!����6���:�s�?�b�_��Z)[��:e�y���BAcWgGP�x������{#50&`\0���0����l�����A#J8�RN��f�����v��5*��?���������Z����w���j������)XC�>ƕC�!�}�ɡ=���I�s�-�e�k�����|��j�	��:Xy���(����G�����T�����-�9)��2N�<U�;�O<�*/�p�|�ٯK��.�O3+72J%��K������3�@�y&7�[
?�d�"H���*G>�O8�½ �����0�L|�1͐�`��1Kb'N�45�gÎ��EMMwnP�n�&��S�N�P�
��G&�`޵4�QP�w�je	�n��Wk�G��}��Z�RfI[�M���yO�f�yNE	XYz1ik:6���~�i�py��������Z��H���+��i��p�wumP=�*7�zS���{_���?��~�֛�����U�L:GMLU�8�c�h<�~Y\�X&�ʙS��c�� �w��U�S��~��K�{�St����g���g|?>>YfgX?7'�f�kffgY�H��������U^9���%G���n�o���9�Y�{��{냥�$�cl��(��X�]|RA���^�q#��� ʬ���1_^7������#��7Io������ACGۄ.�SΚ��z�m�3�(���{���{�YG�6�a����D����Oħ �S稛� �#���N{�%��z��6���+���(�wl����<Q��7��W�u3j�bb�P����g(0��Q0��a|�Xp�Npy�L�.����߷�r��A�{���o�˕B�ȡ��i<�.Fq\����{�8h�2S���yb�Ck*] z�u��WK����W����c^�Ű-� S7H��Ƈ��?���e�&)�������s�գ'���lٹ}w�4����¡��o}[=;>=�P�0.U���(�^a���r�C��|pO�	�׬� ~ɟz�)�t�G,���ivy�e�h�>� �����K�C'.�=�GH��7�T#{c����OU�_Ѐ�P\4m��w���;��}o�������L����w���Ȧ�I8��5�K<�	���V*M:�B� �@f([d |�7�7�iȺ�@�2�@^��D}��/��Ce�M{�[����:�ݳS�����1��EP}stp|z�P�*D������v��3���3��I\����g�}�ùs��)u�Ν��3^���=��ґ=��t?#D�г�㯜P�h\:FzTx��W�jb�ǜ�7��:�":vR�Sb:
:�o�v5�JG�3�����X����vNi3x�(�5 _�\v���I�;_{�Y�`�':�e�7�'�x2�L�����3 ����R�s���3i�^z6�r��c���ܽ�tʈ~�������b�f��-���Ѵe���f�d%��ؒ2�rb��رcf"�f�s�LaH$3� x�KE(y.�	��>��yz��:��{ｶbQ�Y� �(Y��GQ�"�r﷾�-�C' =(tb��Y�2J�|�%��|���4"��>]��V����ʋ\4�%<���;�O��O�}�wK�0��^4$����྾!�:s�|9x�e����� v0���I#�ּh���U���澹��7���\&�z������p����g�;�gU"�Tq�^¼z��}�
/<�ɰ��J��ݠ�2[�p%f����Ufcqw��^v�+�e�鸚�u�R����J��u���~���o����;��/��{�[���w���z���9��6%tl(z�tH�����#��!�[��������	�YX��	�˗����#���~�7�طOy��c�=��e�/�� a�ևn*���p�N��¶�y:�����q��	v|���a��P�1>�],�H��U�;zԉ����.��<T��]�ih����\���q�#r�U�9���aU��2���O�pR���Ӻ�g�!Fl���,J_��͛���'ϔ㯞(ӓ�
�Ε_c`�D�%@=�>���vbG��{�9��)Fd��pO8ʄ|0E�#�Si��	��F^R��L���̶C��Og�v�p�7tp����,zy��]
�Y^z�^�D���[��H/�.��dn߱����
���}�@�e�ax|�_(��q�Foߺ��TA��`���%ɫ���">�a��촧~�G���u�r��M6^��Ð"���*Zl�E�G���@8 Z���|�Fm��"���Α'����Y������B�Q�s=�jPYX=��|زek���|���mo����	��y1��������q)����Ǯ�W˩��c^|%@��(\��# �4j�*�FA����N/rST���,ǔ��A��g+#��k��*�~���=��AáЁ���lX)<��c�!�����˄���9B�5<�?����X+�k�-��X-�v�p�k:��1���|���}�s=�����m���Ŋ�`�6}Ӊ@60�O�h��G-���p��X�u�w#�� u�x(]�:����F�:����e��ٺuS����dx��;���.��g*�&��$�@�Pyƃ�4b�����f�����A�z�K6(0D1*X�̚B�tIvv�H�W����15%cf��-e@��F\����M�]Ӭtf9�j|��͜���;qؑU��P#�I�����󎪏>��C?�'���cph��ɖ�^|��={�!t�;.�� F��뮻
_%���.<��;��o�a�RW��e��v��x��,�6�Pwh��PC���U�LF����ŗ��;�u�Yp���%N�z]���|5,�fG���������~�Q3:�>kX�u�{��0$����G�pE9�f��xOO����5�Q 68�òDr�w�z��}. 
����m���8|��7`>�2\)4���^ǹ�;Փ�K�L��"mݺYa�<���I�4�]9�y]��K�[��  �p���Vt�o�_����No�f:E��:y��*|�g �����s2�X��^�%/�J�ouCDD��$��*x��L�����yc�/�A����9<ԯr�-��LI)-�@ӱ�T
��y�1���鞝�NY��0}�榷�O�P<�0>-j��2�J���J�@�_�9�^��}���t�2�3�����y|���gp�ߣ.��b$g`�������>f���8� ?�sp3zC8�z�;›�Z@�tW��W�Jp��R/�ځ�������z��H_���e���e�C�����W,]��a���zIuh^u����dp0��Pe��Y�Q��R�`��m*�����;��m���]�w�}7�-���,#[�K� �T5z����햡ӧ{�d��XFX�:.��3L�E�9F��;���@b����F�4y"��?�!~*o��	�Y���=��Un���28:��B�=b8��2Y�\Vz���k�ja��Q^ԛo|�2h^�2����3"r��q��}�����r$.Fi�sىG�3O]۲Em���.��_<+�t�6��:.�v�#c�̪N3z�Cm��y�<�Y�p9��
�f�d��3�s�� ӟ�X�����vʋ��X�Ӊ?22��oZƖr��wG�+vr�,[���.��y3à�&.�h���R�4�,�7oR���Z�*��F,i��i�0��)P�!�����|��o%��oG|�#`��̫q�/<t�?�03;.7i^�����r��[#bV�3��N����`��"R(�C9T4�.�	��Qq�0�e��k]0`��4h8:�<$#���������ĸ����*�Bݱe���>\6����'��|V�����z�S�H��h^�iN���۷K�u�#G������2:<�rPX)��w@��W�E��]��Zo{؄,�k������,�#�j@����8 �x��C���+_��W�W��%)��m0x��'/�T���������g:!(�|�+R��i��a�p.���+Ft9�V}� ˦)+���sE}رmkٺiS���Pܺ��r���?�[f�g}H��*���U�'W��a�O�O�\geXx�G�]�TtKW������;��Ŷ��m�pٺg��ܷ��e[�wێ���Medgo�8 �zJg��n��}�:D��!70�YF���-;G˦�Cehx@�Έ:Ò;�IbK��3#ZU������b���l!����V3��Y兏*.Ȩ��4S6��Tx���WFW�>U�E�:��t�o��{=�V���T��O��u���7�_��_���_UL|V'����];���j��v�����s��t$YS�og���M�F���x9w������)���U�}�Y� �o�����h0�%��e���3�-�w`P�X��s�:y�Za]�t�p4�4�_��:t�E#������r��i�[Vʊϴ��O���{�{��O3*C�ABc�W�c���51�GA^�X����S/~��<u��S��b�j�j
��uH��~��?�8�W��h$�.��p-]����)U�����e�ezF�������䫧e���{�Ϣ�/����q���i�����s���S9�!��0j��i-�&,�I��`��p��4vz���y�$��q��I�7���0NQ�觗�1���z!�S�6�lDU�B/�c���_:X���s�3�<�Z#z,*�ʲI����z���J��î'���j��\uE~�B���ND��o��o�_���\~��~�|�O>Y��ڳV��(`�2:�g����c�ɠy�C���O����˯�ʯ�pL��r�|�΍S��+�z%���Z��%�j ���(W�<N��L���O�+7���'��ʾ�v�G{P��~�a���������x1�
�j�o�c��z������p�FZT�����{<����]z�T�{��N���/����I��BtՒ����)��.:�ʛ����N��%��m��"�.S7Yè���q6��J�j�F������燯'O�,��r�L���(]>�@�I��s�j�����n1$��F<��ؽy�wxf��������q4��_�j���]Dײ��C
�|��_w'���֑>��9�9E�����uy��Q�LV��vI&˞�۽Ac��=et�v��W�k��v�zC2!�QA~� ����!Jy.)/ē㙰|��i"�+�@4�(
�![�\���	Q�-�}� V�#X�j�9��߾u���P�ı��_����=��y]�8����
���!L��f�a�����ƈ����9���쓇�#����\� ��3���I�p�G�x�(eB��Cܼ�GY�,c�����{vy�#~�}F|��o?$�_����Q(�P.ճ����S/U=�)#�.�����0���}��S}�1�1���Y��|�<��\��=_�7�Yg�7������� ���|�e�8?����JO���Βںu��k0*��da"����/��(��iI�K���w3�֊����PL�Qo�@~��%���D8�o��_UW�ڹ��[�p�Gu�3�0h"��I�
���GY���eL'�p5�:#½itXu|HT_R���?8��_5iT(���j庻��H�� >����!����*C�=e���޼p��{e��,��Ge$�ZJ�4dC
~�Y�'Wt��@&t���� #�
-}���y�]��[o��2�wL����e�x����6[@C>1ܸg�Fi��<X�&���J4ԁw�rքBk{d@2;��7�����>�rV�>�F�b��B��zf�=K��)�`�z��~hդu�:�iآ�΂�h�q0,�kp0�V@�MF1]00 �^={*9��s�V/��Z!��G�B+�19i� �3r�b����K����kY�U8�����`*&��V��0k����n�EF��eD�����Fbh8 >!�b:�H%�H���B~i�ȳ�<�����W�a���0������&.zʐr����vx<u�\�xQe�n�zf���xY_n�hO���,��;?���H�<qH"r��%�^aL���0e�[��
���7�)��Yɽ�^�J�?��5 �1��{)��_(����|�q,������C��Q��R?�#?R>��{W��R�.I����7�zA�3���&�7u&�{tW=_�W��w㭆��
�?p�)����mۢz8��JG�!����N5����W�Q�2)ʒ��dԈ>:=t0zuսz��7�z�a�8|�X�K�!FM��0l�Șa�ow����g�/�ܳA�{��#e��meێ�N�Sa�z1v�����ya���kf�Z��1J�8��ha4���B�[e��nd�V�^����*����,�t+�C���bqt�'L�\Pbt��(ЃtLUz��8+�YB�����G^9��c:��^w��(l�.��a`��27����it�kY����nFM2�cP\
U�Y0���Ռ��L���Ƃ 4��.f4�4���"�� = ����X�/�I�4����jr��Dڙ�:@y��=�Ƃkޯ���T]�|�oEw�}w{;[���7,��d]�rc�3�2�,��yL^��%<@3��3�M�'B���{����ÿ�����i�b`�:9��z�_�fN�i�|ס�=���IoA<���r��i�*�\O:6��.5��铲d���[�鍊�
�I�V��tc�1�C��c�yӖMʳdfY	��5�w����H�K��Sq����bt�`d�	�p�a�*kR֐v=}�c-���P~�g~�kne�4��)��4%6�w�n����G���("rδ<u#�!�|�{��w�ڲ)fOH��Éu�FU/U��pJ��qbm�wU�x�U/m�T�Y+�e]Ũ,��:tFЩ�7����e�':<3��{��tvʩ_)UP�wc7~�C>��6�ƻx��֭�.��2bd4�n+9��̦ �9�%����X����_?h#Lώ[e$��-2�K^#�#+�W�X�m=��c䛎|g�&2s�������׫=r�:+h������w��]g���7=2�h�c�>�[�)S�t�W�
�� �1�������ϝ��,�>���|�<�VhQ�N ��<��f��p�G7*f�un�T��� ��8z�(I��qO�ʓQ��=���pԥ���*A���:����믌��رM�,�c���!����`�H���k��2jR�d�"�m�\�2N=n� �9��y�h���V#�q�ⵌ4zu�ƠT�n�fa�� n�O�Z�8���."Gl���8�[���T��t��1R�Ϻ@��1 P���;���B΢����+�^-|�	e��N?>z��r��2�r�W֥� ���z8�lFa�?�Xc��w���^����o��l�4j�xJ|��w�1=�ߕ�$�p�|5�R���SwuhWwW��S>��/��Y|͉����?R>��#�Y�F\���~�w˧>���Ǐr�(���1~��|$Ɛ�R(N�u٬���
��\Q��LȘf�}��G~�7��:��-�8��Ϝ�(�¥�2�������1���՜�h�=:T�C�a�����.���]c� ]#05
�{�]�Ҫu'A��g��b�p�XL��t��%��Fּ�8��BY��Ú�c�f��M����Ѐ����L�0����+1}���8�9�A�h͋����g��rϽ��]��`�GÞ�^��j`��k a��J ->g�������[�F�^�uF�'L�c�|�[ߒ>=�����׀Uҩh@�r���cG-��^̙7����2=�>��D�3!d%F���3&�e����U*��	�:�1���adN}�$
�g�q!�SAa�`�,*:����(�����h@驰��J��� 7�HY���ث��:l$1����_��_�����w�#l�u�/�S<T2v�`$0
�2GHH�|@���%^*��L�������k�Xx���o.�|�;e�l)�Sⷢp�y^�O�u=߿�&�B�8��-~IOt���e��V8�&�'mi�0҅aB��3p��� _�xL�z�����%C����bS�ʤO�l9s��*լ���#=u��9U��20�lKw��������cѤ�B��O���ϔsRLq���d�|�Yy�|K^����x����qV��P��Z ӯ�7 �P��5É��92���4o������&2C'��������W*����� �b��tX���%vf�$=���Z�v�a��,�G<:D�i�[/���k�xF���3�����R����-#���1Y Lo��`5�
��� J��(���I��Ƈ�I�Q��T�����ǈA��P���x����,�\/�-�Y�X�~�p���E\���4u��cH1�N�~��5AW� ?J�F��svN����C���D��c���9��sv�p}����I�g yNx�_+w��஗i{��M��닒�q�֧�[n.|��uh��~��I���o��(���z+:_�ʗ���{Ͻj�����O�Gv�^��q��ԛ	�����I$}�_QR:h@�0��]v���ͬ_�R6tF[|=�jZ��4�8*3�(�Ka���* ��u���4:��`{5+��
7�eGX
�����N��a�\�P�Q9 �&%P.�!_4�|��|cڡ�{
��p�+yW�rp���{�ua�C��sҌ�g.{ӛ�H��Z��K��k��PU�͜9��8��vҡL�9�V?S&��P�0��Hㆸ1��h��yZ�@��~*
�ͤ~�e��La�P��h�8����l����12��?[9^���o�#����&d����Q|^�v�)��<��y�H{��]^E�3�EY�MYF�	 �q������n5 �tY��|�n�o����n������駟.O>���S��:2����kү{�����z������O�i�g�쟕���y�W��_��o���a  �����OuH^�W�f�p@;M\�� u��S��;p��ƣ<�~��t]�:�-�e�:/۷m.,|�O�'Ӯ�G�������`�&��d��``d&��Ƈ�J:LӰ9�?.�j���?�Y7!����ݘ!�Qb'�(��ɂb����jr���X���F�|^�Ϧ��r`���(���(�� ]�{7J����N��n�Gэ��,_�_/�$+���F�/KxGެ�Twn��6�ҋj����/z@�Ξ�)�H3� 8�rW���>���t4m@*=��/��|�G�Jg�{ �h-O 06��]J���^*��S��~� ��:C�1 
�;��@�����s*�D8FJ�`/^p���)q)������&
(]A�NC��Y܈�	��`�9�J������w���G|�#��8�?i�����y����DGh�{@�޾�>�ӊ@����YiIa��ƔW���Q��VQN�a� ��?�L�)|Ɓ�(pq1�C�'���'(�_�c�xOU�Q)���ɂoG������H��(ιS��+�T!��b�L
_7LQ�����S��Z9x�l��N�]�:�#�W�����	 ����Ӏ,g�e~F��M����A7�L/S70h���@��g��`4s��}���;�S~�7�#8��˿\~�~��M�Y���;��:��A �u�:���˔���|�u��f��lFT�c�F��RW�c��Pq
�ɑ�F]�qt���SE=9u=�V������¸�Yam�
�R��ȢIYw6��,"��Ug��UG���mlB�xR�Fi+x� ��Ӄ��77;�6�jD3��'ߌuxT�##��Y�_�je�z`�r\"U��#ll�>s��X9x���)�"ԧ���ڬ�e�3�$o�s�t0�� �]�-{����6���%ڼ�~�k>F�)+�'!�,\�SS@�#��w�R�*s��ͨ��Yd2�KF% �TH�^问r��
����g����So@��5�1����b�
�C�+Ct�q��Q	��<\NCsi�Po,��Gq!�(q�CJ�JE��C��$��������� ��C��z������a'����a�(,v������:=�Y�(N�1�-�
�O�)҄��xG���_��;��1O�6�V.�а��s�K���fk8��ʠ���o�k����6*�2�/	OȐ䜝yO9�g�zw;E��&Vs�|딲dN�u В�gÆa݌w���^x_+pXf"�nHE�^;v�#��wA;C�Ⱥ(֥}�_Px��V�������;?W~��~�S���hv/·�U�5�b=��z!�*�z�Й:A��z�z?��K����469��:� Ì�Р�NcA<FK�t
�Ϯ��)�A~6lɆ��S���ClȠ�� ��X�I�T׍�x0��¨�QǏi��ʊEő���aeh��F��o��c��u6|w
�
ݱ�S*��<
��a#�ȷ4�	)q!�p"Ч�Ê�+�dԠ�(x=�H�2�_�(`=
 ��G�d�p�#�?����3�|�|�k�xwK&e����E�1���կ~U:��y�~F^V����#_G���#�!�%�_d�N��S9/���x� Cȧ��F�)���
�
0GC�[�������̐8�ai�Μ9[>��OZ	2r��~N�e����W�TK|��i+��� �P��*p&�~���A_���9���x�F2��e��Q�0�iQf�x)�@
�Z@>�/�~�i�C�^��Ba��/^/c�Q�����<�v��Rbq34qM��Hy������yɯ���V?#3,n㣚�EĢ�N(�}
��l�IX)��.�*�wl+;d��&	�Ya�2�=?�b��������6Xg������gPʯw�FO_?2u�h�1s"�\�P��#�m��QoW��rh�2~��y�{����s-�P�� Y������_�җ������|�3�M",h����hd� �G?���я~���G���
�G���X,����� ���|.�y�a��+�MQ�,�fT���-�Z�o¤K\ �	#W�'�',�Ĉ�N����٠�o�E8k���H6:�����#}��)#BZ�w��t�Y�&4�����a[x�:/tJYQ\�u:��.�:9|`�_)2r�B>��82�X���;@r�������5>��8�nC���	�Χ"�$��,d��ĳ4ˁ���Z y�Ļ+ ��C;�t�g=�"#��}���ϩ=�ڳ_��Q�}_��^��8��9uX{�3_����>�Y>_uX򊑄�}FF���E��r9���CN�J���	Y��2ŀ �N����
�̯7�}�0�`��!����I�&!l�U�:���k*!�Q�Pܟ9{�co��6o�XDF�Fo�ѓ4`0|N�b��-�g+�b����rd����ʫǏ[!�a��f�rO7_e�w>�U�`�@�'ŀ� ���0'�2���.`X����h�v��7��o�����Ji1�t����7]�Ռ���S,ޝw2V�G�	�၍	e��k���F˦Q�c�# y�0(�6ﾊʟ��|@�̎]����[�L6�ѭ�2r���3�4Xv��Yv*�V��F6�w��T~R\�F�I���<�,�"��#�(9z�U�ӳӢ��m���rr��8�x���(e��!�,8�r�뀲�rY�e��)W+eͻ����<�s;�����{�#�>Z���둄����,���w�� \.�������t�r�]wx�S'�2�r��6��T�>�H����
�ͪߋ����~����}�iK�Yg�+�y���J��0�D)��ϐ�xz�Tr������+n5Ȳ ��i*�@�͒�={�����[[˾��9|B���tRa�F��4lT�,���S _���Fu6��z�0�m��FFJe8(���[XT���^�<�$�L(u��&�{ա�T]e��P��˕˩��/Sϝݥs�Cݢ!F�����ϛr:���SV]����*��h��Ǩ���Nh� ;@Ŀ򠜔_8�A'N�g)ANqR.�1�%���ja2�U��\�6:����/�1��g`8���Mʉ�|ʾ�:hX�{��C��p[���OI8��S�����W����퀘�OQP��� �h����[�i=t��d��d|��P�H��޽��a��薲�;�Px]�ҍC`�� �4��0Uñ�|!t�z64�X��|�0�"�Q�q��)Y�+�iX~_��	��0(B��0H�Gc��C��O��|��Ҥ�sT�� ������QZ��0X��ş���h$'%P�e�:� /�(�{p'nd����wX����+�#�B���M\�OY`����B4��o�����|`��JA� ��cD�#��t�X�Ϩ�4C�T�ۡ�����H�ta0�Gիtz���XN�%�����GG�4(ݘ�W���ޘ��p�w���'������E�ތ�x��^���o�JUWя�aK�8���C��US�S6L����?���d�������_��|�1����#�<������|ZF�s�Uw�ث���o�i����<u4>���y��d����ፎ����w�s��u�wI/����������Ӗ{ҧ�ڂN8ۍY�י7
���}r�� dZ8ї�B�8:Kt���g	IW��|���0�e���0p�҈��S�����C���A'�ZN9��͇��TU�H��uB���-ҕ!!#�u+���i`�1z���Q����Au�K�û���W�z�H��M�����(+�pH����0@���`I�db�;6e�m�n��xĺ���q�(r޺dԈ��o�P�.L�VɈ����	����z�YF��:d���Z!�G!�)��n�V]C��đ�ӷ�қ�?�86CP��c��%SY8�'�ӑCoƧ#B�K��{�oϞ]�W�p��ˢ����u�H���O{�qٽ{�*y��� &�#N��� �\�T�A5b=�cF!b�PQ(�d�[%���0L���L����j��,�s��/�O荰Aǟ��H��i�i�9���ӟ�S�����O�N��RXq�l,^�A�Q�z�1�J�C>X�F#9>6nC<	����?���޽Ǽ۵{g���;�ta�yu�"^̗��Y�=� 1*ZY� �O(�%W��ߎ0j�C��E�)����A�`p�=�'�`wJ����E���|�}A##i�>���}�+��oc�2}����>O�&Iɖ�݌�H��(��4n��Z��SQΊ2�q�ӱ��Ƙi��Ο;'y��kt¨��	R) r���[�p�#��p8�t>��~���-��ۿ��ZL�R��0u,�G�\י���g�Z=ɗ�߲5>�(�-#��� ���O�a�������g�K4]р o%�	�����F���#��C�F�/�#S��?�j�A���^�h�+xE]dښ�zY6�QbF��	�p����>���;�lQ��yJ��P��
r� �w��t�ꃍ�r/��b���ޮ��t2B�H��`D���@,$&>y!Ȋ:�^��j(�,<e������152f8wF�BM���t���[;��~ιY�3i�aθ��^�DGy��C��J����B:�Y�e�;��V��p�"~�*�,pb7_4��DS�a�+F_�]��q� #7��9���r��aOsJ1u��l/��i%�Ы{�p�WwyIx]��\P[��a��������0R�Q�����u3j`��,¥Ң� ֱ�E^*?F��
��^&� ⵌ�8Wt[�*@�鹡X�U����i<a	�{M�B�G��Gt1���?�T���?[��`�)�"�@h�B? .��f�y�Y+�9Ut�egJ�4�?yKÎ4�[�ė������[[�cZ��n�h�v�fff�L��f���7�	����[��=1�y�g����e������J���ú�)zg*!9/X����](�.)@�t�Cw����;���*a��Pr(�P����]u���uѨ����d�46�t����pA�B��gX):鲤��r.��F��WOx� ���2�Q�|Q(g�9���%%S�c��C�+��3��іx�'y���{�
�]~�w�<��g��A�/�S��.J:�����ė��2����o9p�;6�i���c奃/�?���/�~����Y��垺�1��a�:���:�.y=e�,���%�4ӹ�a*��	mk��<�
o�	��aD��`P˭��Z�����,����`Oٹk�{�a��,�GF�G��]��#�N�C=�蠎�I�)�>�n�E�1j�h,:λm���t�WsYa��d�8�*WO��ER��2j(/�a��A�A�_��{�����bc��L6"�i��0�r������a�=���#�Σ���(�� p�\�J�y%�Wp�e�� �)����x�S��!��W����^�H�:�:��_���Fھ	�E����m ��uH���Q��2jz�zTG_V�ƨ�J�����#5{ʞ�1��YM]^OX�&�ʍ��P���(��1���'��r����($�H�:x����1p�sX�]��y�Ϊ�r��r襃^,Ŗ5h�$I�&=��k�����.E��q��0�M)F#�b"�`�P&,LCy��A@e�dq��6֬��as+��.iҀ�0	)�u��a�&���g>l�"ErB��$@�8sA�z�<��3<���_Q�@\�4I+����R�Qy�bؘ�����Sx0#7+ł�#�te$�Ra7J��p�������n����ý0jt���[��%���ٹiT�{��O�LFm���H4�0y�z�x���!^ۨA���P������O���=S�'%��IDŧ��e�F��'�#��,�}��O��ﻯ�'�'8ݗ�E}���`<c���Mo�/yw�ͷX���0>����y��'�t�f;�_��_��}�k>_�§�)�Q5�������Bi?�NϑWKI�(O>��i�.�g�x��+�DbN2F���,U��H�\ԡ�
��j"�`+�^9�J9|�e��CZ���s^�1£�u��6��r���^c��2x��ǭ�f&��p��ӑO�sՎ�Uy�����3���G?*�8�K�����266vd��'�\���P}dk����1S�'=�����	��J>��A�1"��-��@xZ`��4u��4+��4�?yR}E�tz*OC)<���\��B���S�Tu��7�p���=vQ��q�����_�F����[��Z���3�+���U//����+�j{�?f�,#�aG!���������9u�0f�~�(N���󫖏v��B���'�ȓi�#�Uy�y�\�U����ãۤ�cv�zB�2��J`H�4�0T\wO*!�Ŀ�w���jh�9y�^!���Q
.H9
��D�x3Z�����r�<h R�b�<��;���[���!S^��s8��㗾�%[$�p�V(�H;����J9��J,G>m�=Fʕt��`�=�����L�<���?�aKb��l�X��<�η��)�y5�j8�����r�P�N<�(�/��bX�ݼy�S�o򇡄2eh��nj|cf�Aέa*���068ݔ��&ʂ�h��;����'�<�q1E��D��	���,}ݽ�'�U��g 2�ީ%崸�<;Wz�꩜�`F�\聱0v2L���{p�P��g�Ƹ��/}�˒��T��-j�>Z>��Ϲ�E��K�R�){ɟ�����!e��o{���i��<xԳ���Z`1�A�q�r�\;,��E�L�0,M���&�������ʯ�jyI
p��5 ��(�>��s?�?�.2 �d1nHr*�L��|z�E��S�[�u��>;Lm��������Řb�Z�h��YW�a�K�JǍQ�zݾ��t Ё�Ϩ6��E�Y�nA
2}�����?����ŉS2އdH�e=Fg�h�Yc���ػ�W=`�TlՕ�b��-����� ����6�z)~G��q:��,k������9�y���	_��Q'�m�;8��A�О���݉�2=��~ݸt���d���3/�T����ߗ�����G�*#*:0���-2u��ڎ�|]��^w�u�V�������:~� �D��,k\�#u�?�p�� qS�y�4!?hAVX������Η���g:'�����}�I���x�|��p�L�Dƈ�}������/JO��/���e˦�r����O=U�|�;˾w��>��|�^�n��
�>
@� 4Yp ̢Q��)<����-ͪ@��]����	 o�y�x��O�q����-�?��?*��X��/��ʈ9a�r��t���0�<�!�X�1�)����M:�c:>F�q�ҡ����=���pl<��3#��&'T�sA�~��������l�hl��һ8n�YdAp�Q�.NդlXI���\�(I��c�����߸�wJFˌ:U��
e��`�����
$� �X1�I�I_~�E�:�/O��Yc�?+�9/�97?���_S8�U�2�6N+_�����l�6Pv�����.9�6LI�M+l�ƥ`�흔�(W��h<���w��^��.�Ea�C���kw�퐲�qL�i���(�������f_iH�S���I+P��Ϝ>����7-�9v�!�L1�����I7�W�Ȥ�Q�:�=����'u=�N#f���S'�C��>�m���P��|N�a8��y&/t&��l`V�_ɭ����::1����}��.�=l����.��@{��d�za|�~s�z��DN��U���Uf,4�GUb�C�N��|��]�E�Ʌ�w��evq��,�ɐQ�~���DǸ"�AE�b���J'�6�H[�FZ�� �:���fM�;DJ}`M�+�C;�z�O��Ɩ����b��6(q>U��_1
��d��Ԫ���dʆQ�͒��{x
ϩ�t�#d,�
@g�������{�[�2S�eNf(��JPǿ���Zk�b� SI�=��:c��;����/���󮏌��)t�"���-���z�E�<��)/��6d��1�M�'r��ɕ�ZXב�4�4�0���gΖa�'�WX�W3��y&�����!�z7/�b�0�Z��KpDV9�؅1+��CH�xqp@��G������{���ţ0�ꏭ�(X��s��������O�",���
C�Cn`�\����/�Q�؁{ʻ���?���^�;��S��c���^[�T;�&'�Ga��Z����a��8�]��m�iv��'�rX��A�E�ҔrN�$�\0Vz+,^����)^�٢�n�<2UpA��ŢW-�E�<�K.���
��p�)�|"c�
�W��/N�g���wC`���@���{ʧ��������I׫��g`��v��H��������H�}��[^:xУ��ON��K�MC˔�eC��h"��艧Z�ea�9�$�]x~cc�` �p`̰��[n*��s�iA�kF�P�ߌVpR�ꔼ�����e%���NY����)����m6�~M=��o����Y�L���O���1�r�2�v���#4� �������p�4_����s�λ�.�N���z��0t����� 0�5r���)'�SC��R�C�:�|/�{`^�z~�#!�8�؈E���D/Ig]ʼ�>�(N��(MehX�x��SG�H�PGU�TO#�h�1������Ћ,J��Ay�%�Gj�^�4����//������+G���m۷zw��� ����+u!u6iS��/�~�a���x�=�<�aC'�S[/�Z2�^�Z �I��@ˋ6$FO�/���#����Vxnҁϗ
�gū�p�6���ч,2�>�g�)SӢC�f��dh���s�M�C�@y�ɷ��7�Y�zG��zº5 ��R��a
�O��6jPz�Tnڿ�a�ȡ���A�b�ZNb2�{��;� �1O�D%b�+�����/��G3$�4��Ź�U��W�%	��Qʂ�5st����a�z�X-.@8�	����'����zfA3��|����.U.�Pp��w�w<�I3T<G�mQF��������ʹ��/�~�wu3�+�CY��/���w;wo�l�i�� �%����T�E'��{g����2���/�1B<*6��X�K^+%������鲅׊���T(�e�X�J�F�&���h�κxn�|�+_+�%� ����*�������ŷU$��j�i�������������z��?���o���e#���x���A�F9aXp
�u���	� Y�.[q��X��N��
y�dS�l�1�(z�3s|6�X��WvB���}��z��^������g���x�/�H���	���n�����������w�0jh��ICP/�+�R�៞�3m�Y'��r6& ���X⻮���#@�|�u��D�5�3�[;vn/?�3?[~��r�<�-��FyPW���c<�l��;W�؈^#%�]፜�d��=*.t��	#EJ�5�u���w�_��Pu�|���lI9!O�g�<3��4�b݋t@z@~NA�i���?K�����H�@,�&?��� |� ���N��B9r��r���r��#�g��v��X����(%2��([��z�T-�F���?�e�3v�2j���H������A��z!䃜�l�˘2�Z�7�3r���?[��5�bUn	���٨�����)#C���NLŧo��L��(�ʨ����<��^��>5��\X���-��@i��9�e��K�
��D9���ʊP��io*_,�G�U@��	+i3�����`�D�v!���
]@�O�y��J�Sz;T�?Q��J�B`��#)���P���w���8v9p}�-o���G*s����ɘw�s�{4�:d�H	a�����Ȍ�*OOz��u�n:'��Ѥ=i����7��Jᨏ��Q(Ì�y���Fc�f�i���	#�NW(Y*L��Y���``�v���h*%���Ni�)�%�_���q(G�	���&�eb%�2f�̗����Z�Pl�?y���K��@K�ҍ�Y�	�4�+�\�җ�l��G>_=�i�G|vF��>��3g������9�vF�X4|��!O]�p޽Tέ��Ǐ�����'˩�'��쬌��gN�����c�62��[��4�E����~�犰�
#�#JċS�O�<�:���yė�4�F���+����A-�G���n�;�{9!��uI�|����3�<4��ϩ+p@c�# �P�M�'v�{�.��qU���k����
+Wج�Q� �I�О9v��.���y����s�ջ굀�WD�< ��ԓB⠍���Q�P�S0�s��|(�䇎��;�����P�T��~����37�P.^d��be3�#�y,u��Q��	eB#N��3#�8�w���?8�.��H ��	���k1j���*�g:�!Ӵg r=�y\o�}�J�|��T��H���|�M�%`M"���(-����{��r��w���n�����{)�
��`i�i��2\M�0��<�*o5F-�ϊ�9������B��V�v���_ �q*���B����@�I��ׁ|�)$3�Y���	O� ����'�����e�R�i�> �TYc���y�3�5�W�[����)���U�a�tW�L��G�ܽk��Fk�o����P.G�(=cKyzh�R�x�B���_(��[�z'��-r�
��ں�ψ�3Q(7�Q���g%�&cŠ	E�њ�em�7F��\>�S�o�2!�3g�Z)܈�<�\>#c��~{���}���O�D������S�(�������ِ�X@Y#����ԩ�>��1�O�w�Η�yv�Wa��(� �����jz�@o��k�ʝpL=!C��/�c`1���?����;�r8:�\Dg���ܵ`�S6�3���3��w�8cǊ]���W��e:��ҏ�ttع��NL;E���(t�����/��Qz+~�U��\�T�R��|��+Fz�1��p� 
�^�%����|�j��+qѓ8t��DTz�:SiR��!�AHROTSaU��cT�u4���_<�^���Q�x���8NI.����?:dA:ߍb$S�)� F2�K�= ��o������������g�2uȮ"Fvc="z��J����#�Y��
Q6���,�A7�zڑ���.�:����cI��G���8�{փz����u-��(@"�`z6�tb�V+�B�J��<�����!�j����ޅpl��&�et	6ֺ�8�X��s�
�BBZ�9�pipu��յ�C�0 ��Y6<G�k�T�� *�?��!����f��5�XYW��ʎ�T�s��/kq�L�����Y�L�@����lqd{/�ý���R��ٕ �;B�0�KO��ꩠ�aȻRVf��/�Q�- ��	K�����DxaWM��ؖ�*=�*����q]Co+}�nQ��cԲ&	|���g�P)�I���߹��.s�g�rM��ʥ�w+�@T=a1;���Xtz��M�C�Py��ߧ��βy�����;o�����o�m5O����1���'��lS�-������)�r����:��;�W�"2C�QF�69WN�8�ь�ՙ6�Xr�'���9H��h@ ��!�a�GG�!�r�D��V^�X��rY��"�;H�g�	�ӯ�Ƞ	�-fx������f,nݹs���{ֆ��ri��?� O��<��xS.�s�c��ϸ���7\E_�q�@:S^uepi�Ns%/�b݋V�"���FGU�0_+�=����J/�g�U�}
J9یzt��d�Jr6�F%��H�p3�Εv	�{ｻ���oUl�>@|�����y�����������Q��?���/����f�FC��{mM,��c�����>d����C#�S��_�_"rF�����G��|'o���Τ�E �<�����T"����; � �EC�ȴ^�=�C��Zv�e!qMg&V�����r(��W��{0��P�ka��HAU>���F �(3����޵�o�pe�m��'R>�O������B6*D	�s�Q��|�IS�<��dI�65��3T_C��de۶5H��O%�E�^ko������\��Po�褷4%|�y�Iz>�ʩlL�,��{���G�"���o�P�ḯ�G����uz���a@��3[WUl�N��*�(FW0FԻ��ʨ�z���L���I�i)���W��	����qCrK�Bu���0�LE,X�7�(�
E�0ЕuIK#�q�JtR"�؛�g�����c�	�&���7�p���|�^Gǂ{FqB)#A�(��QY�e�E�
ǁ_�b��:�yT|���3qpt��%�+�e":X�|.+;�U���.�gd��C��	�^yŇ�1ݎ>Lև�﬷�i{���4�\i�9�*o4�YX���0-��Ws5J�b�$�ɣ�QgymH�7����LIǗ�E��e��& �)F���������q~��,	��D�*�� D�9[���T��ho�����]ꑬ�!�g�G�
�����
-��'���)��������������xW�o��o�_���Z�����rI�Yd:�53�@E�Y�|\+,ɱ\�+����iA�_!3�݁�1��$1�<��i�"�S�ސ\^�(P���������p��c��J��P��y%Xbj�9�R����a� �������x��!*3�?�SZt�>�1��'���!/zf�O*^ ��9�����^d����a��,4�;Fw6e(�/��̀:�\f;�B
g�HmPovD��z�C}�ۭ�� ]��T��M�ޮ}�-�YCCނh�����&>��J�8���%$Z���:�ֆO>)������<�_�����)���25�0��(O��`J���vX*˫ ¦��C�,�p�3�Dj9�f����i���4�X�|+�5-���{p o�}� �����{�+<�� �i�����c�>�W�`�h�e�,�JAB֩KM,�G�PE�gʌ2=y���n��0-��kol4�:���2�;Ej�6�r���q���� �l�q��ġ�X߃����pЙ�ge�Ƣ�;v�G��?�����P&�I�R���8�>�!��#t��&֌r�A��p��{w������/0�LB��AGT�娋.~�����uhᒫxق�_�*3��?�Ī;�+��X��lɼ��8�G����p��K�(�!g����!e�h&��n��>�y��3��c}��o=_���/x�= ���e����ڄ�����vH O�<���e�怤��>�Q���q��~:�
��F�:U��s��@�������x'�5�2����K�_��Ǌy��W%�?9^�ܵ0ޕ�b[�n��K���7����r�!$�ʘ���ԧ<b�bjFi�c�����g1��^*'�ư �"��|�Ѽ�]�䠌�����={9�}S��^b���ӆϖ-2jz�$�i F���*'�K<$/*�Vτ˰q�w�?�C�����N�*��AC�6���u�UJ��.�`){ߋ�ܟ�p�y�Ù �!���s�\])d���\)��\{��8}�3����D|����0��y[�l.���Fw'�s�ϋ̫>�������3�3�x~��\>��ۘ�#0iX����~�����р���L�i�S�����0:��2r��wzĒu?��(�s�c�%4љq)�.O[���)c�]+,�a����t�r�y&�(L�¶������V1���XB|�UF��$\�Ea+]T�IzR���?����I�u��cQq1RXgI� ���|�� "��)a�M>����X"6|n�sޣ��rϻЉў�,�+:��pg�r�|�N�\�o���Jǃ���0(;��Ȑ��}=}N��m�d�ð�k� �z��o�G���Z�����v-ȸ�i�sN��������QC��TYq��������uxb&T��4�`>��@Y�����5Q�-�Y��뫁��"�S��:Q�䑼�`��rş���07��7Ȉ��Q��Q`���g�Rd�&����?��1���E�]Z��_�v3��oCپsSٽgkٶ}T=�^���@lc�~�*�@a�އ�u�S�rг7*�!�c���K���2���b�/ׁ�_"?���U�xV��$�aԐO%��Ə��r�Aô��!��qv,�h�i�QV��ѥ����ϴ^����lЋ?n'�b���+����@e�u)E��ݠ�r��o1`=�&��������ןG�����߲�ȉ��We?F���w��I�&J�F�ʖt�o�κ�;zڤC=`�
k��Q��#<���{hM	Y��{��@�2�?/I��n������O�4x�`�Ky��L?��Bʇ����9@nr|�ya�/"W�՟�Z庂�Vo�]d��g2��I��@<t��ڠ�� x�����J���uu��\�rx�����Ѹ��e��Av��Bb=���;\�ѳ4,2���]~�g������V��?�'����#����ej��JʔgʑC��^�bp�VGF���<�g�@+#F.A\��-h��khY/�S�Qޥ|!��!�K��z"v�.�V�' e�ES�i̠���Bd���Ņ��HH��B#��e#�����ݕ`���G\/�A)Rv3QiXP��n��*@�f�I����]N�Gz�C��*�� (�8�ɱN�kG���Dc��' q��=[��[�����V���5z���D�������Y��^��}�-���t�h!���]=Nˡ4�@5?�T���B]�W�
J��~��������= ���0����]�%�?_O�(��-à��S�/���
JYc�FB�2�\[ep�l�/lS�X��M��ber��G(S���������b��I�z�YGx�6ti��+���Ch�n��6�H(����e	,�}�R�ꐸ�_�G���Լ�@z�� ��������|��:��O����7"}⊬���a7��o�9�#�ژq�<3za�3i�G\�kɘ �>��s*r�Nǵ\��qIW��?똊/����V��R�~k��V~�2�X{��Fh$7tb8��E�m�������~���}�{o�����7��ʨyR����k͐����Љ�-u���T�(#��x��[I?���l�g�P�[�P���<�Ў��Hy��r��ދ���i�J��F���D�z�˅
���,L��hW

�d/!@	�{0�ՙ�_��;R\I �\&M�Gn�����kB$^
�N�I�8=預������C@���+�f��\����x��.*��ظ���g>0Fb��t02!~����������^�ASQ(T~("�1�;''���OP��&$��9�x&-+������Ϻѥ�@Uq[���#�{���9�����:/��C�o���p&�JP<_���q�)@ϐ/��qL��и�;|�۠q7�|�G\�m�GDQ����z^��G����*�����q��o=߄��ˏ���S%~�Ŗ��\������i4����	� �S�g�]v����]%,+������g]	�Hm�ZL�I��Kt��=��N��� �C�w*A_9�^qB�������z�%�ةkuu�7-2���E[��/��/��V:�'���P] ��/��?���5�#���=�G0�9�cF8�#��acDLo�{c}"��]M��ԭ[��}�n�c'(�&8E��#q�8���ѳ��'cꤟ:y��;��B؊p�%�� �"���������uX��j!�d��a�tNNj�?�H��|b�Q��V�q�!y�n #(Tμ�3̡�zZ,zEɆ��r	Y`�g#[���zn�r<�e��8r�� +�=,ͥ�W���¡!%O(3y���۸*<��e�fx*.h�����7�%ƔT���2�gT���l��P�h��E)�f*�3sT�A���/SX��ï�k���/!��y��ާ���R��̖R�X	K=��|;�7* ʆr��a���`a,C��1��c� ��?!�!�Z�v%���H�����W�@�ʴۇo��6/�ͩN��a�_i\A��񩾊�1���`(�ڹs�׊�C�FY00Y�C��n�Zb��aT�+�p�Q4B=��b�	|�D��m}��,+��Z1�p�e�p\��xQ�`'?В��2LB�hv/l�'/q���0���.��!�����1Ĩ��4�9��'�5>�Əz'������o9-- ��"T�W�%��U�5�B���xي�{4L�����y@"t�Oeͩ��y����T|�k��>G�� �!�Ƙ.	]�(���dy�_�����K(���t�1d��0�x�̹�����0�uF?�9*&�z�
� ��K��r0*�W���H��%��6P�SE&}�a#�҆�1����Q��[o����(�3��Us(�"*+;y.NE䫢��:3���E���]K- �JP�g*�4���
����e��Ǩ	���y�{T@�_�C��Q0��#{��wJCO!Y�>�P����؄�����`Uq<&-'�F�Z�T��T�YJ7*<�A�+%*����K~>�T�IG8�R�[�W�¨��]�����T��@�;���<tM�A#�Q��avz�5ip���~�s����8�h��kA=�w
\ƕ�r"��'�I���a���Η@9qt|�C�޶P��ް±�#�Y������G` �&���������џ���ۨ�Lz�4ʬ; ]�e@z8�]>R�t~Abj�w����)�:�y�� ���\���:�A��ү��2SwA�}�������z{�l۾Cev�W��%Ռ�Q@�7�ȲJ�u��G^�NN���M�:���|�%F.@/�K	�:�-e��g7-U>�������6W􌴘h�[mr��E��UΔoZ~�t���̱�#Fʢ����s)\����\����25=Q���o�������'����r�	ZX���E�ٳSx-�*�8��t�߅?�#�^+�\�@䎷-��@�S�[��+�+�j�L)#dF��N���c�+����'FuR:U+,�Va�0�F8�a �!�\�e�hE��q�4�G���ع�����UAհ�.���"��qy��_�1���?<4\z�!�]$(6��y�z��u�'?�0��hh�rhނ#�s�3�g[+=mv��&£��`T̰(�-䁇0nXk��)�ֲ����FY!��߃g	���r��4`��ܵ"��}�HkN�p��WH�2�w8�b��JV�cd�E�s�(>�O�G��m�v7�,$4O��r�<8O�[�z��G�_Q��+���䉪/|��8i�咲cw�:�%[��/�2J��,��W�Cq0lP���\��������Î���v�n��o��o��~�����
����4*a���F=D�}tC��i34���T�\��|\o+dI��\�&!sr@L���ZI����&�D�;:	ј �n�U�� yfʙ�a-�JCa\p�#8�'�JϤ�ᗉR�ȃ�KF��ВW�T~�?颧6���n�lӷ{�f�|�*���gw�̋_�\d��[b4�n�p�5$Sew�����/~�|���������?�184�#Br�%d�2 /�,G��1ؾ}�HE�y�y.&+�5B����rk�J2�\I�����]��Ͳ�N3<��P�>�m��ڨxc IXw��HE��shd>���Ҡ�9t��\䲑�zvY��{q��	��� d��w�юP�@�&�4�X�'TX�Je"\CMh��:nzČ�P;@~�8@>��k�gKoO���YUhvBy��*���]��o�Q�pYD���1�qM�����Ż��
��c#5i��2m3�V��`#��O˰1��s�%o�d~�ԉS��ݻ|X![bi�����'0F֢=�_����z�S�.Y�+���^
R~�5�o��Wo�V�>~���t]�xQ��4u��NȀ -�J �s�o�Ο�qv;}�3��ÈaG��;Q�a�1������H�ϨA�S'1b	}��F�?����@�C�?� ����t�8�������nLxJ��T�JЎ����q���n��#o}��^���'Fn08�]8W�� FV�z1b���?O��B\�bᮮIi�A���V9����P��/�>}�K~�)?��+]�·㭮�2��ep�IWͣ�������k�P9 p�*�onpR:1����x0/��"xB�������4=e��M7���y>��M�����y�;��\�,�7�ktDz��t
��={����/t8Yl�m��!z�@�\y_�&@.]K̏������W����up}�F�{{��;�T�Iv�{�u/�q\=o�\�^'�3���F8{50
k�,������
�~��ܕ �­�m	�e�Q×ty4C��Fǧ�95�<��'�	QJ�48�#�d��ޭ�t�Y��lP��Êt����c���s���O^�_�(�XMO������t�~���s�\r�k��/�W9�HON~f?
X�q�T"��!;�V�P`c�/��OxߦM�˶��|���$ϱ�	����W�k5�w�0��k�_7�P�`/�T������la8 ;䝞?F���x�
"�1Bȗ�1����b�.x��FCi0e��ؙ3gˉǫ3��c����@�QL�+�ܓʟ��4�4JtX��C�('��V:����>v��z�kj���I���㵔1ړj�c��K��u���*�G��!���m�U}��WܑaT��s�bFf���Tn��N���z�Q��C�-���ba�0h���wy� �9�u�����7W^��~qW�s���c
�3g�`JI��d ��)C�+GΗK�ЫL��_:/L�C�驘��8��7���\>��?-���>��G��F��- E@��[J��/�[1^{��s?�s����t���w��ϖ���������xy�{�S6�n�9OhУ�0�Ֆ��9O~�\f�w��P����:a�}�5��!�A��#(�8�,
�o,e����������5;Jňs��z���� ���]H��}-�R����P�4Wi�ĝal��g��}�o��ԡ �"C���hy�o�}~�fd$FjHW����7�����P��&�^����p��zpi�	SS��
,�Pf�*)�c�ǻ�YQ����u簁o�U�䅋o}�Y��q�� ��:9��Z���ɟg�snf��<�7�N��Jٱ}�elR�&��f�5Pd��g���r:�����|�?z�ʍ����2發cx��(֬�����y:*aGFe@�J��t=a_F��p�����}|)cWu
����D4!ìy�$n��w@�ì�q��1�;_�4�&g���R����~��s:��Pƫa���Ow���A�.�¨^P.4�L?��n.����鳒sv�����S����ev��WU ��5�7n����XS���J�n6���Z����s�<����-D���L�8�;CV�*t�G��s�t�,JF��t�^k��Ѷ��_�N�}y�̔�Yړi9N���L�0G>OJ�sӸcT�|����{����G�����ċ���/~�`y�˔��6��������=�'�o����*[�O�������O>��`r:��d^,��T+�ˠ�?e�����qwU�fzUY��o��;�d��s3��n9�.�
��U����{9������� �0�i�G�����u��w����N��u��Jy7~-�}��������ƵB�y@��r�)��4΀�a�z$4(��o�}ꩧ|(��o~\V���G?����'/�򊸠�	�VC��򟟣'���c�ޣaL��i�C��r^|'�d�� ǹ1�[)2��	��� 	+#��5�M�O� �������"�j1�¨r䩢��-��N1���!/f�#C�Gi{H]~c����G˅scetx��ٽW����qϞ��u�P3@Y�("#(�硢5�2٨��a�����F���i���`�M�������6|yxbṛ4|�C��՛��KTs�iz�3Lg1
��+�ciۖ�e���� ��ܱ�kn��v�>�S�r��)Ou��Fv����b���@S��vۭe��]����ÙӞ�r�"��)��r2ි�5��-뤫�F��b�Q��r���h�oHzic9v��?wQ|@�-a���v,���M�ДE�=*����Q��	p��㖺��5�к�pi���0RDW��]2jz�{�Cue���A�p٘�Yw���sH�"�92�3���ؤ����-�Ψ�_(�_}�:�e4B0~�P����_._��WK߀GtY��}��,����_~���a�w�|������#�=��R�rǮ>��/FD���9��0P��&�"k��:�Z
p	��$_U ��k�h�Hg%�O�8�pE��}�w�7���I٪��W��҇9��D�����]Pݯ0�Hc��A�A��9p��Q�,�c!!�����ѯ�Y�X���P',��i����[�6xT�)�Гǵs���W�eU�I ��z��*ߜZy��;<C�l��c��x�m�-O��s�{��vϓ^+%�-�4�C�4�����;��bQ%����U��}e`�����]�і����y���Ҍk*IEO-^܉n�l��>9K�����L�8�|�z[G�L�{��aυ�t�񯫜>}Ƽg}�/��ƒ�c'Z��Ze���\o��\��,f���{$#�>M���XLMÉq0��8s��d�����z��wzh��q���w�q�q>������c\.?����|����o.��=~�y�'�r<p���/�s�%z�i+t�g.^���w�,z}�:<��0T�3�fE�v`�-7;K%����-��5�uk�k��s�Ѹ���!g��}垻�-CCÖy���l�|ӹ���9��׋�F\��mu�J{ɏCv0Lώó�R9�0��/�>�-����D ��;~Gl��w<W4�U��F�Q��������;�v۲e[���OIN&ʨd�ȑ�edx���p�#7�m����������ү�H~��K�᜛]��H6�:� y��uCY��җ�T~�W�a�ÔI]0���]��9L��_�O����ma��{���*OA�=�O���7�S�(�T'92��S�7��2��{9�g�v�G�"�]Xw�f~~���ҁ���(�g�yƻ��Iћ�!���.�ɩIK�b��YP�Q[A�
�pU!r�B�l�CJ�}��C�����\i�e��%@��<�$��3}�Mo*��v���$���\rd=/�ȷ��m�#�
�˙�W�9(�m��*��`���^3�U^��,Ф��0`y
 nu�q� ��]���a�a�>���
̊�~-%x�g�ЕfdQ�=\.�v]�f�˙Sg�PI�M�g�O�-�?��Ν��s>|�|ww��ן�rCf����:�U�u��t��ƻZ��[�S��#d���0�708P��������=W v$=�̗eؽ(e�+����� ��aA�bVJ�K=Z��ߺus٬��N=d�����tP����,c�5"���(��d��C�Z�^#��˔�;A�`Z
왯I��z�w\9��E��!��0����vZ ����%5|����L�|=�ܳ������f�o�>,��n	G�-v<�tP�u���}VU����+4Y�}i������~q_!X
�G��F��2j"|8� ����x�	;>�_,�O������`���<���رW���΅��}���������/X��>�
�����qn^��c��S2�/�n(d��c�3�2�d4}�O>U~�W~Ÿ�#����d� ��Gi� Tƃ��g��r0�w-��:D�p$�Bۢ�{�,��
h��`$�!6ҡ�W7���Q��FMύh��x�� B�Q�R�ׅ�g���h'dU��@�(ȕ��}Z��/�\��Jq	��=����J�b� �7y1��Q�䇒�3�_�l���NJ��N(�P�4>�O�2b�|�3�.��ǫ��=n����Hٲ}�G��/4a�e�[qJWOW�ȰRP�L'B�i�	��Ư�������PB�u�'�a��,��}�Q=2M EL�/�:�3W���=6ڑï��]V{����k5�1�u"|̒vK�p��"dku <�J��Hh�q5H�B��S������I�O'����/�cQ��qǝw�>�)���I��i7��k��$����xG_y�9z��W��"�'�5�nxQח����1FS��K�G7`�~����261&ڋ{�:sʍ�L� �ԉ|��M�(P�)��{ɨ��؍'�D��'F�~��v��;/*������22<�Q��I�B��#itt���%YJ�2r�9���Fc�d��K.�Z����\�O}�)h���Q��_�|��0l\���~��G�?w�:�g��.���Awj����pF��'F��Q�^u�ۿ�[�UΨ�Fd�4��T�{�'Z��$���/�T>���Yg<���ݟ����s_�|��_,���O�/ɨ�T=B6��U���};s���j�8���ޭ>]��	9����-=2_R���VG��b�Ʋ�2jv�F�n�Qç"�����e�����z�ʊ��e���3Dp���.�4!�B7q]��L[
W�V��\_;��W��{�SI�L�3*¿.�|4���3�	��C/�\��쳪�������/������|����+TƗ����o:-F���K~�Йr�(b�&[���xMĸ����C6�ô�/��Q��0�*_t#מ7��pq��k*-UZ9�������UѶ,��{��4�a��ϡ�H�)�����Rύay��`РD���ڵ[r6e��㆑�o����Р3ʰZY�_k�KX-�k���尚;7�'hb;�;��Ԓ�8�iN�eJ�=��;|p�0"ضʚF��J��������^���z����0p�r��ѣ�(\C�˪kq�R������������� �W��")��%ٲdK��;�L&����̬����ǽ���f&���$��ĉ�ĎK�H�z��BQ�$�	�������Ã��| ���p�<�yN�g�}��g��}��E9�f�DK��9��!3n���<�����}o(j����.m�4QjN��Q��s&���T��g�2��*�0�����O��/���5����\>'y�w��v[��#$��8�>��)4��-L�#l�-�T��B�Fӏ(o��+���F|�3��￢�d�s�Q8m1�`���XT����ōvl�D;?bG�%v��{>�Ƚ[��;7h�`���)f��`����y�ڵyɤe��ԧ2u�T]+���3��wsm`�3ϦR��z��Gڃ�~�}��fz��n�N�d�1x��5���'~t7��ߢ�0�X�i�z8;�q�ud7��6%��K��b�<"@���,\8��[��]ʷ��+�ۥwᕚP����*YF��:��W~�W�o��o�i�@b'8��M�lܴ1��)>Ũ!�@A(��:dޣR�Fb 9J�ad.,´h�ׅ�E���o FC�i'LmT[By:�\����QFf��/3~���,��W`��G�Q�BbV�G~�Gڍ7ޘJ|���w���>�:�.ɩ�9��w`ot[B�9�1�,u�r��(�fDcDb��mwv���wR(q&��3̈r����̽I����p𻒑Ơ�:}_�IѨO+�Hyh(-b�;�Z�q����(u��l~6"\�B�=.Fl����ߐ᭣���'�J����/|�}>���+�T8x��п����t���~7ۂ*��6��M�AVJòe�������7 �A��"��fQ�m]&�y����Pb�6���xj�\wB�]!֓YWS���4�=婍�+
���TL	Eg�}U�I�R�l�����������N+p���!}�׷��z�#:M� n����L��(�����F�Yi��-����r�w�����6�%�"n���<_��fN��[BN��-����+B�nHY�x�ȔLC�P~=�T0F펜�9,�7_�EK\�C.�G�����(aT��p��Ka�.�|���!���%�p�N���٠ͻ�4�ͼ�▶�M�n��|�w�D��Pt}���B��f�2��+�	~:������q�m]����7�9��N�TY�{*a�W��8����ës��%�3�&��N���WC�W/�z.����yc[���O}�><}c�Z1 ��n�����w�����7����]�lMě)�Ϋ�SH�e1��o��i��!kp,�EI�gd�V�^yh��������ՕU�?��F��Ƞj��L�d|�0k��ϓ����h�C��s*��pR�����,���Y
�h �+%�T���|s�`Q�����*��(��q��1�!f�ը&��v�H��HǤLY	�n����(v����O(�O�wM&=2-��
R0I#p�>�S��Giy���3J�#'����p�=t�_�`Zd��[3�Θ"]
���5�w�%t��?t� Y�t�h��©u������:=�_���ޢ���#�2�߬*
�6H��S�/充�<�,�gI���o_<|U�ܮ\#cJ�o���F�7Ud0c���ť���-oɅŔ
SY��K^��B�O]�c�� �1�3(�N�����g�X���:�>����v&��\A�C�TbF�@�h�hFI1}b�c�k�W��5I�m��ޑp���S�T�B~������C���l_�0{y����fo_�&�[���V��.��?|��O�l���ÍdD�g�.q�� �ڙ�[(,�M���g�~X2͎��m����έ瘟�0����C��2r���_�R(��ؘBN��C���@�/��<�.�i`��a���}�����|�qj�L�՟�"�m�~�A屶p��v݊\#�i�m�ʿ�����RC�0M3�J�/��/��l��z��ޖ�o��o��KM�I��:tı�A�H/�H�@��,5�#�Q޽ȓ���װ��1���
�}qO� B� �/����t_�v}���
˯���Sl�p�N�ޞ�]s]�Ї?��y�=m�3����=A�}{�p����<t���ؿ3�~!��afN�du2z���3Ѩ��s��.(��v�ĝ*_xA�C�De���r�# �aN	�i,|Wj�������Nzf�s��G�:;���y&��#b媕�ꫮi��̩)������.ME���ɷ�zT�O�r�3�����Яx�B��S���}��X���<b�^3���.� ���#M���LB[�;��GS�ہ����Ve�1ڕ>�:t�P�A0-�֔Kc��SDX��(P����Y��^��3wNZ��b�-ȴ�r�/��H�S��XT�[���C�$-�`�ކ�x���;�����:7L�{�u�ϿR����έz�{�����ח���|E�o����|-�Ӿh�k�%�MDw xyq*�K�.�4�y��Ā'�w��@R���۱��F�lN8�[H���s�
L��~�x��N{�W��̷�lAXJ��*\��2���3ez��ʑߜ��#Q�Ϸ'2ya����+v��m�]wc[|��Ԙ�3�\�뢐;��]m���/��d�s�m}�꽣�Ϭ�(�d�,����,`�Of�$�N�I,:O�jp;�9�bO����{ڊh����O�����,�Hȋ���ۮi�x�;�]w�׮��N�o�9oJ����0Xjt0�_��_l���s�k�3~s�̌���1B$��Ⱥ ۛ�M��FYj�az���"�����b��?��4�n�Q'�ׅ��Eʌug	���I��8T���J�+��u�W7�DY�����������ڑuY7�i�i�}!����R��i%��=�SXwEG��[�ze4��9_/\D�q>F�˒���)JM6�(g�u�ߒؔ�)Z�����d*@�Ր����)/$9JH���D}8{"���Q����O>�t*4
�hx}1��v���{����cO��?�8��4�%���z����D���ԔBS� x�d���^O0%gø�`R���t�H��n�����܈�E��D_��Kt�ùF]�ϗbM���l��ݺ7�ޣV"���iۣ���y���;�謴���o���o��#�\6اf�����M�!�s�I�I����ˈ� ʹ�Ԍ�7=uF0Vo�z�6�0H3�G�Wͤ.�iUܮ�tk����-]��}�����r˭mͪ5m�ש�Lȝ�h�ȣ����6w��h+�ߗkAm���m��Gǿ�-��vQ8�t�V[<>�h��!-���j.�;g��N�l9��g�շʡ��b�����#YqR���!���U*��Pf�}V#�nQ^^xqK{��R�]~�ʔ{�qIf�����gv۽cW�uZ��~"ih�f�ާ?�����}<e���T_U����g!���<�B��U�Y���t�&`b��癠S��0Lq�w0��$�\��������;��O?������Ҷb��Pj�koy�[�ﺷ]}��Q7�#�t����sC&)�m�F+��T%i����@��i+�2N��I\r�2;��;Gًv�kvZ�N�:�n�e�r�$3�)'
k��ҩ��� +y�����r4Fp�ZN��Ӷ���~��\����-)�L92��a˖L������eGy[�'a����+���mʎ�n��l�p��1U��E]u�T�(�����2pu�Lw���{���^ƓqO��(,�E�Pd��g�Ť�{O�h��{�����fӥ9�5�s���6�ű@Pd:����ѽi���
���N���+��� ��w��D;n�zP�{}��MY䅉ѹ���-�A�����d�
GT�������_�'֠��K�>�3tƓAB�K|۽gO�ʨ�K���:/�8t �����][ܿ?��>��сiC�Q���B��r�z�f��p��w�������a�����`A4u�-x�\{���k���E�~)h���m(@;v�l[�no{v�z��bЅBKY�W.��4�C��"�U��j���w�OR�O����7�[q����m��햡��H��HnPbw�ړ���|*�07o�<����:.$��H�$����֏?�x��oT��ia�o��3��x�d8c�#x�����4N��+��M�<�<�͚Ƥ8NMWB"yH]��$z���yQj���,6�9ͥ{�@�NnԀ?N<aYm�a�^j�\4n��=�N�<=p߳��2��t�?f'H����d�L�F�.d� �I��8Ho�s�WP?�?̣2��w�?t�;�bA(�d�|�5M���̍v/^���tv�ܕʍ�޶�~j�K��]������x�hׅP�G�I%f�:���j�p����N!9�F�K���/���Y���"d�?���ڗJ�7����^�u��ԇ
�n�,�p��N[�F�z���)�;ˠ3�|�hN灪���z��r��2ɁIyNrӁO�6ZY�1æ�N �kGCu�=��H1�|d��˂C�A3��ڜYN�S�N���]�j�d�i�׈�AC�A��	νYʓ��}�)�m+�|Zhl�%�a�K��N,��]���u���%Sz��p9�����8��cq��g v��8��FC�#�{���B��c��9r(\��ږ�{�'�?�婧6��_|�-�Β��;�x�������εh�Dmd=uf�ڌ��;�q�KpM �����A�┓� �{��4r��� \$��D��{*2������o�(���ؾ+���x�������w:�I��[���Z�"yr��y����c���=�\���)�,?-$���?{<.Ika|	���\�v��d8��脉r�G���	2r.\���pJZgU��F9d=^�W0�3�L�[X��ώ@p�!�7��hΛR��E¥4b3�.Ⴉ	��qv]Ь)��0��O.�}'�G>���}���:L�V�{�S;]��dr��x�{Ô���L�<�����h�ի�w
��& v��w����R.�=����p(&��^��R���+��h��B�-�7?�����.o+W��Q��P�vm��r�Jt�ۣ��#����.��P����#���]	�@2���4�*��21���yU�y�hs�'�2oj�K�k�w��E����!؞n����ڃ�z(���t���n��[��)^ziK������ݙ�_��L�ر-�l����Sk���X'�����t N�=�?^He�����G�㡓��Ԝ���������	�H��LG�E̮x,^�4]M-��S��sW�PB�����Wy"7xuw*�����q�|��Y�Z����[~��zWw��K95r����=��l`���_z�΂��֠�+[���F.�50��ɴ�޽���4vȝhw��������������r�t���╫���v���91Ќl����v���ٯL�z�bF�\}2�x�=/������%�;�wt�C|����,������jߡ��N�Сp�����ȗ�pn�:1��:6��ٱ�=��3���^n+/^���^�vl�����ێ��i���lѲ��ط��}�\���#���2.����/��oV�>]����I�? �ˁ���|�yN���+�.�o�C�B�L���t
/t�S�_a^t��-�����+����K;Qܔ���ύr�-٘򘕶���p{-@ʜs��	����ب@O�55�}�)����}(���A0b.#���<����G2�Tz!CdB/��X�D;.����qtn�b�a)�A����$a	�M�6,�o�
��`���8�Y�$�����Zc�*���V�C�Cc�iA��L��
��w�S2����_�ë�R�)��}����|��ys�����C��������v��rC�+/�-��J��Qr�2D�u�Q�w���޾��o��=;��=�,��<��t	�ӑ��^zY���7G��5F��Y��6�d�j���#�w��Ic�C��8$΃����_(���T�O�W ��٤t���^�N���*0��3>��]��Py���ӥ�w���d�Tg���� � Ι�(<�k��J<>Z��Y�Lo�6�\{�	[��N�lbű(ڴ�{����v��m{���O?�6?�l������c��NɈ���+X�m��6W
(��S��8Y{r �-+]��I����u�S�QSL�܆�k����۔�m����7�����9���R���d�rEx�3j��sv��E� ]���V_R�pp�D��F������G* 1�:;p���ANɎ��>p��ѩ��&�_����_���^g'���:�{���E���S�i��:���/8��g�"��Z�d)aVa�(� G�N�ޡ�����+3GCt-�ù,�����]�7�_�J)W��<�1���6�5k2>��"cq�NN��4�<�߅9Pe�&��x�!�{=�Zy��`�gQ6g�N�WNNX�PYL�/��vb^

�2;L���4��m;��T�Ϲ�c��w�]��R�QpB������=��Xy��`�A�֙rL�=>^�Y��gz��'�C		��+��Bjk����b�\����qå���RG��3N9kM�m9g��s��GE����?6��t�� MN���x����7���琖�NCG_H��Ct�J���BB� ^C�=���o�ˁ\���G},��pJUX2������:Ϭ��,�߼��T��+���~�!K�!���.r���Pt"되����n(]FZNG�7���ӎӅ��{�JL��."�1|!�2�=��F�ݶuGZZ{{ߜ8��T�� ������n�YF� �D�s��䭍Sl(<�#.�OU'!ʧvG��g��{ʰx�g��)5��e�4���t�����,N��0ه��xҍ@ܡ;0U�LSی�����f݄}W��y���2_8�^;�J�pUѠ�]_�7+�AU��
�9鰍�M���q�E´�i�SI擣���|ႅm�fr'�m�ҳ�e��C>�D2X�1�U��@���p��%s��	�i�C}K���M�|�����]_��Nf�q?ߤ�w���=�+�	��s�닩��as���A�OCa����S�)�d�ŗbx�~J���E9��O}d�H�<���1r<p��
!�L���Ձo�u̿m��W;��D|{)��C�_yM[�hi
�-[^�t��ȏ҂�̭�BQ=�ޠaGYJ<GrX_���� �3u��8O�G�FO��2�x�_*|*�-;_��S�Ý�ezȰ��=��X(�e:����^hY�9��[3��%~x6�-�M$�(7�w[�mذ1�~V{����SO>��X�P�ȱT�,���~�ξ�do(;{���w�P_(�k�,�S���(7�k^��%��D;Nk%ƀ�{��V�H��� �H��.p˖m�И*߾}WNq��XL�aevo�s�L9;��8��&��44�/(%���.�\�A���d���~�T~��1wN[���ť¦�f�KC&��u��Em�n: �ԛkH��w���V��@}�8���=,�L`�&�eJ>��C��d��_����4N�LgQ����s�xF۬%�}��ԦS�x\�+��O�f�Eq�5Y
Q)=�s�D0��ओ��F�,4�ň��wn�WP��zV�a�z��Q0|�ʣ@C����k���[�k���5,���7kx�Gk��tN%aG�.�@�f!1f���SV�px=\�6r��"%<4�Q؈#�Y9�߯8 ��S7?�Jg��!n��r�X�ٲ%�b�i��˹��+�n��r[����W|�ܦMͩ3u�h����8a	�m۷��!8�n��]P�^/�9]�0��+N�����?5����� =���wt����.���x[�-֣�a�CZd���8�D������(�!�~TiyKc�IyL��[�8m� �+�
;�C;���h��s Klbt�m��u�lۺmk�=gn�ֵmA��CfЮ��"a���Q�R�ʑ]���V*�����t\��jCVXD��E�t�q8�K������{�A1%e����v�ύ�L�I�bp֙磍��W^qU�����4���W��s/n�A3Z�{��%d�>��ǉ���W��P��v��ypP/���8/��8rK���!wY��X
M�WOk<��]f�.��j+����o����7���$�G�\}�c�=
�Aߐ���u�״M�n�ӝW�^|�����9p^O.b�p%F�����O�)��"�)�&¨�ULU���a�סS��4�fF5R����'�& 8��9�t0]v���C������-fR����)7��P3*��(Fy���(�Q�m}%T�ӳ��p�T�}�/Fl��߷ߕ��C �h{vu��5k��+�ݠ��oz̜�gR��ys�*�d��������iǶ�����W���ܮk!7%ŉ�C�m��SO���@���]w�B�`��3F�R���a�G(�����^��K��ҙ�	�<p��S�T��7������J�K\���J��|��,�2Ȩ)J�\��� ⟒�(~�wZ|�p�ᇸ��&�����~J����7ov^��x��hޗ%A;��YS����S4%K�JC���=d��CGr}�zp��6�'��=gĳ�*���,^�,�o)�#�m��5����L(&���U�Oy�~��o���
���qE��&f��|w8��6?H��c�I�f-~�����n�)/K�3wns�-ڏG�J��!�=3�i�Cv��RlX��9h�t֭>j�6��O*�'�Ȇ��(͊�-�?�;�j0M�/~�;���j�oWa�y"��
��d����W�; �����e�_e��ӟ
b=v4���Y���7]r�R�Ѕ�CB�TO�%&g��=O)5Lv��<��#�7��E�r�:�q:i��t�\}��\�XO0��Oi�)�t0]>3I�⢕�mA��Nء���B���A���Q�*v�9��N�*�nAiiN����Sn���i��fj�\|�s,^����s���Ie��ڗ&��e�Ҳn�%.��-�pv	�Q�ӐMR��%�/�HӼ��7��^~iK3]FAr� !��j������{s4E�ShXh�1�{y�KSV��wR]�k�S9P�jU秃�a��Н^�3��xSV�n���;����:�W��e/KE2�㈎?_���I��]8�+��sg<\��0���`���u��:/�0�nBz�0L�޹!/�ߥ�H�?7�&K��[�]r�o�a��Ӣ�L�W4u�-�Plbp�j���ֱ�7l�׋B:��m՚5��̶�?ڭ)*������"VJe���97�����{sʉ�1FAZ�xi��YaM!SbXhM��]7^ڮ���H�Gc �.<i�YF��E���%�8�2<��q�&�F��{h��CZ�a�z'G���nPXy��
Z����k���6ID����v՝��P/@�.}G ��K�>�'�>���a�N�3��V0Fy�C�p�UW�r�}����O��]�֮[�W�l��o�_���E�#`zɩ��T�їIPCcV���i��i���#��o�\�-�a:��@�rg�l�N
��, ��ܨ���	��~�@�B�>ԋ�[��)���� �P,���E,.�_@Nwr��ʅ{Lȣ9q�`���Ͻٹ�e�;Ҵ�{����v�ֶmN�ޖ�ؙ9���I�!0���.���R�;�?���Tmܰ��x�-in޼�}EOgyjGA��(.:�7�pC{����K�9v+�H�z�a����aM�w�,'�u�/��­x3��p�Դ�SO?�#��g�����{�X=�L�yHg�{:��3��x:gH{ô�XeM���0�ש���վ�ۥ�oVS.x_��i�bՎYk�u�ڦtp��m�_0� h��HLb�r�@�騳~����:�G���i��&�ԩ��8J[�V�Phb���K��w��
�c����{�y)��ի׵�K��������Tl(Unܾ����5�r�j����Q>
�^,���ء���/t��-�u9�3�}�{:x��/�^�:�$����AהYsf.}���o)K��'���� �'75 s�;S<T��=~g���/�e=w<=���_��m��~�V�)ѳ���oW_se����1��OB�ELO�����_JM��!�0���F���JV@�����f3*]n�W��;8sU���a>����1r�|,4:t���e#��{v��p�K$�C�l����]fÌF�6���E9��,�#E|��j���z�7b#0��"C	�ʍ]��4)@,"vW%2�R��0ҿx��m�����<� N{B`����ږSc�ol7������j��/9(��s������H~r��!���,4�)�����A����tux!`�\rΰ<]yG�'O����o�q
��e��ʖU�%ОeP}�� ��ѽD��:&�DQ9��Ok��40��,�0ޤ4��Wn��aȋ޵E�)����Cy��V[��SjXmB�� OSzL�R4��ݓ���D��Ӣ��:6���Ӧ�B6o�z���h;���³a㆐-vY�vf��T�)߾�Og&<�/�eEtr������@碋���D�{)��y�+��ʴ9Poɒ�)'Xn�w�ץRs(�*瓙ަ<�Bw�����D_�O��s��M-é ]Ѵ�u�~њ��/�+ϹV����Nf���(<�+�r7�k).��0J�0��*�ݮ]��Z�Q�&oLpC����Ȅg�7���0�zG�xi�-9�x�ѣQ9l0���kV�7��b��v�%#K���׋�LἮ����P���󛄚��H�)�fͺ��Lv&(�'���O�~OG��^���y���<gJgð�Ci��m���U�(u��z2��A���M�_I�~;��u���t�~i��}m�!���B�F^pt:4���W=  ��IDAT�����+ڊ�F���Xx������5|-��nL ,����ʄ�XB,:<�<p���&�SX3I��,^�,��7n���+�r����ukC��`޵#���'�S�YX�N_��WR������Ba�-z�����uq��9�0WN�?'&��Qn۞
���Yѯh�/��7�
l(܀,�VþND�Jh�:,[�+�ITޑH
�
�r�_�7���}*͂ӥ=�S�� 2�xR�Ь��FY V�BAi�L��pz�\K��kwhLyAo��)�s��Nޙ5���.�hP|L^}�u9HbY75T�xu�N&_�zm[�tq�G1mKӢ�<;y�y�y�a����r]�˪]RN�6���W��:��(o�^jmG~����t�m�g��_P(��/B�+��,2�l�sE���6�4���i����N>(3��N��'"�8�ۛx�|�-��xg{�=o
��:i����7����Y��S���d>�b0t�P~���x�#_Oƭ�♳�!.�^}��k�5�ђ�1��3{V����~�)W׮s��%�_Xx.�h����P�蝅@�Q����TJM��M����o:��0*��b���kI�l��t��Ѝ�t�O��ӓ�fQ�\�o�FO9)��bC�ʂ0�ݸjd���L	\r��PRbdʊ��X7ܶ�k����=k\XU�����`hN4l�ʒ֝��w�\Za�ZJ�
����ވ�03o~����3��I�7^#�K�o�2\������l���C)�)f��̯3C���u�+i��%�"�J	<4���B�� ����W����XL����?s��N��>� ��0��R�ǻގ�:e~�}u����(:gt�:�	�O	���}6�3����(�S���-����O�������ue�ł�> �|��]wݵ�[��VZ"�B�ub݇�A�W\qe�y�ɧ'ӻ�-�|��X�|��eN&�S��4�y�f�iZyo(?ڑAAoK�E�ۖ�b��b!=`�)�4���}�}���h�>�X��U��[o�Y����5����� T@��}����7?5�?��\�m�10G�t�-�rw����J4����������e�o�� ��/�����~�B1w����{U���o���/�%)��⪫�I��/O�U'�}ʈ5Gp�w:�����0��Rh��9��g�O%-��eW\�;��z�p;�o�׮��v��7���^	>��V�Z��RS'}�;�pA
9 ��-.K�邍��t��x��!�=���#��\1Q�t�0oR��qW�`�s���N�q"��-����x' u.:~��V�\�L�mǘt���.j���в�.^�tK
�51"[B���q��{Xv�؝u�l}4Fz��3'�k'��p��p�ڂ|�[���y���c����;��m[��_x)���۶�۷]�i�ϼ�x�Ҝ�߽kW
�m!<)FnOWF#ʝ!���!�MsX�����2�ÙU���d�p:ڟ�^�p��U���w@�I�s�Þ���p~�~k9JWt�)��MoJ��Q6'/�j�/�C�Rj�M����~w*��Kz��iT߄;�9�Ҝ�QY)cU/UOSaG��5�������ȁWř�F�4�v����'��M�`�lݶmk*�S,u���-́����b�,�=�w��L-���)S�;�M���<RZο��nɢ%�ɓ���Y�6'۫��,���̙=?dK(��f�$�鿎^�'yO�"��[�M5 S8Sg�xp��ĕ�X�v���db*��_J9&=ʅ)e��e���v�1�GB9;:�h͡}1h;Ѯ���}�yw�?����}�WR٣4��O�Rf`廴ܯ�M 
�~�r�����7|�/�� *���xܙBů�����T�5��?�d�q�׹Q�!�C�/	9�(�Ή�V�Rs�4�����$���>8��Ɯ��J�Ί�p�.x=�Tn�����ӹI0��L�tq5fi�F:
�{uL�����rҨ:!��g5~ʐ� t���?7y3����7;��ӈ��1̅»w�i;��v�껍v�����4�ڶ���B��mK����^|%���8km즰^����+rW�2�z`ͪ�9�T6y���:A�/��?�r@'#KJ�wB�:�q�:]�V�ޤ|
������0L<9��;?t�9w$����B-L:��5[@��pu@�=@k�(����n]��t�y`�@��!}"l�9��y�;Í�O�>r5}5�xD�t�ơ��6�~�83��U��^mM�3��W	,�����e�e��6Y�K��6��KsУ혮��t�G9�8�zۍ,̵�Z��L�,Z���Z�5�6�eKW��m>�v��Yo�_m�"`
�-٦�Xt,,��=��	���������.mW^yE�,���KG{��)'4�	�t��"� �ٳ���c�6/d�5���zK�e��M1�Ж�§����3��I�--J��������k�h�i�O¿�,¯L��g&0)����U߼i��紧�x��
�tA�#��9��D���]q�5Fk�/I$�_(8/J͐��5(��h�����~b0OK���sjb:Bϴ��aXAg��-���q�_O���{Z}М��a�+�?�\
�&eGgd���+���bR�L0wwm��RnBa�Fo'C.6gד����m��P:���㐭}y���{�
��p�j0���Mp���av���k�h\�E��]�^�Oi(�VSx�u�:��G���L@��Mʇ>'�!���x����(�����������N���V��e��g����Z�>8����������'�O]eZ�'��9����/�O�Iu>�oR����7�	���No��?�C)�6ԁ6Tm�u�'�[�t��-[�Jq �=iZ�b��r�>��O ?m�oݖ�t�OZ����(G��J�>M��+� �C[��|/�
.i)'\?{�/���2�r�k>�6H_²g0�r��b�'��m����a�{�i؂n*~��m����d�͵57�v{���C�٘�<�J<�ԓS8����"�����r��=���8�f=���g:����)���ˣ�X�ݩ7+xΔ��@�8v0�pN��+C��3����F�W�}>Ἦ�)Й l��,f��K��A��G�x��?��t�0d���������Z����E��F�&ӎ?�O�~ ����:s� ��!8��P�p�t������8�@kw�Y����Q�S_ue[��!a��,�p��X�� .Z�,\B!�.[��2b���fh1�k��m���?���uA;��0%�Fa;�;��h��^a��u�L�o�Ȱ�Ur��^+M�?%�ѳj}X�އ���|N��0[ydر4�1Nbv�����b�s,]y�%�y��	U���/[�뚬�(��X�������Si��LKyR�x�'�w𥃰���O�,�L�(���.����i��0>E�) �䩶�7k%ڛ
|���R)�XR*N����`*�E�֮��v�6)�@���]�����,�O���Ć���/��9m׻�����BI�/������{��ŧ��7�c;i�޼����w:Qr��!���CS8r�]�xI��@�g�իV�̒��1����pxd;}{��?���� Q|����4�:�<�� �¼�+��~���3��I:�����	���x�Y��F�Ξ�C~?v8�)�U�K��K6\ږ�XJВ���s?�pޕ��hP�z�Rj0*�c?�R3ZS3Is,x�[�u�Pq^K����i^/H#G�4).�-}����De!	O! �%ۼ	G�ĔJ�-�����N{w;�9~�ړsȶu�../Ͼ�e]�1��y��޸O�� �h��n����R���e3�Yn���Pn�M�{'T��6G���K�)l�y�aR����~���N���Q���K��0o�;�"���_������
��1j���(�YkC���RJ񙭮=�H��<����N#������ѷ!�9^�Fq��J���u�i?�y�D�FgOߋ�:[���PZ�m�[�6�ZD��P(/��e��g��T���7�[n�%�Y�u��ń_����Bn���N��ঞ�k�A��8�xp'��<��^���Gy$wв���e[(A��o8��l� ޑ�gx��	�ևP�D9��ޙx�>���\k�y����O�����n��e�L���k,�Q���{���~/�M�ޥ}O�t�L��]~�kE]�ltpfp�m!B��nkC�tӆ~��u��,�HƟ>�sA�Qi�1H6���Q�*Y�����n��_��Tn�����H�?��?ȩ��a�@�I�`gXA�A��7�9S��>.������y�)�\_3B�	�%t�Fh��k��6��9�R����|�`o��AYS�Bŭ۷�Z�=Q�L΄	�S$�$�����ڴThtv;#]#1��Vӳ��̘f2��iS?��ɜp$�Ϟ=�R��ʣUa��#�k�X#Ft�u<���Za<�n@�U��u��0�S��0U�x�J�����p㐥goZ�$\�^�����fOPV� �#�v���r�p�a=��3uj`S��)}Qu*�	M���*�8��a:S���^�
�4�8M�F�s�^a��+�v�%���^X�Y=��+��`b��U�I�s�[(������YK�*�y՟o}�S?"���H]�ڟ'��S>\�ګt�)\@"��Z���ck����M&�[���ôk��w��W|P�I�0��S�T�B	!���v����vv�^nȈ�s���b��1�sƒ��T�#�֚�5�RV
�8/�t���xU�*�8���/�_�Q~s�Eᣜ'��6?;TW߈s�-_:��x�e�-o���������ޖ�Xx�6	���.���� �J����e�љj�:S
P1���C��z��L�v�p�.n�1���k�3���w�(������G�ӸJ8�C �r��bw�R(%�tZc���2{��r��΀����h=\��d�m�+2F{�3M�X�[�uxp���(+�B�\�����rjAG8��F����"U0�������LA�\�y���s�&�x���9��ş��(δnH�z�'��uev��rѸY��[�Wh��������H� �w�ę*c<��8���!����h4�S��gIG��3����VT�
?��t�ݠ+�{7����i��^�G�n��1�Pgv����Ah�Qʏ0,g]I�w��;Ń����7��c��i�d��W8j�� m� �G�5m�}�\���΃�H��C<�>4�9�Ů-��	��B�f`_���{rǓc,�UCٱ_�(�vb����Cτ�J3�~�R����?���/9<��_��sCi9q4��5��F�]�.����b%KM?Qxr����B�N���$`�g�R�!����I�f�ΝSJ�t�/�^������~:�I��>;�8C�z ������ids�w0��D|~��<��y:j�F���E��?�a$�{��ߗB*w<,3
���nk­\�"��~���b���8�6�e��#ջ����/�2����c� �G@�[�Z$��(8��;˟���,o�f=��^o}�J�Li�L
_~��V�m�0�?�FR�ߙ�ͦhO��#i�{)����#��0xƉ�R�9�I���Pt��U�i���Ql�3�Q����)��C*5�x��4��:�>T�
��(���_Nw`�d�6C�锶��p(}JD[[��[�tNvHj{�ֺ�A�S���ۥ�R0�l�@Ĕ���q�X�N~Plj�
^��S���f��J&h�e9����=�݉��>����9m��5���*���c麠��}��էZ����f�����g�_���+���l��T�8u@��o�!~�e��d�SaROI3އn:��}����W�3���속~���6/t�5����n��Y(�����#������e�i�������c�������'f8����oo7�tS���}�=��m)�(~��9��}R80v�p�~U�Ӂ��wp�x�
�kRYN2�IF�� Yb��"�48
�E���~[۰�"��z�zXgC����)�2��(Һ��[����eA(!�R�x`�n���Z ,/��d�(�M	<������n�`$���	��6[߶I�jL�޻R��� ��v��+ׅ�I(ZԳh�w��^8]:U/3�aZ�:�|�L7*[����i`$�ŭ��w:P<c�������{wߘѫo�E'����Sr�G1�W�Q�&����C���(�/�IP��>
S��)rd,_o��l��l@�ӥ����;��I��bpb���yy��k��:-�ھ6jP`����_�-,�j��6*}�E�"�n����ϻ�c}��wKQ��TG��j�ڷ0������Sx�M}	GvH[xm<�Ȼ�~�>��ߤ�C����<�\����(���ԃ9\5q0���w�+���w��p�U23�s:�;��~У��C����V�������@���'�)g��v�D��j�����%���\�~�G>}��m�ƫۂū#tOcf��~� J�) �����;��;�~�NQj,L��8R��4��qTO0#�nRe�L�����J��.޹�j��g�W���S�ܽ�ͽk��)�K/�Ю�抶aå�-LA�2J�߽���y�y�֡2:�eK��L�j�e�q'�C���\�G�G�2�Ǩ	ц����}qy]hi�c)3oqA�;\�2���1E+�s�K��)��i:��2ݨl�SbF4˘҈���=uf�.��'��+��O-�[a�2��X�Ѕ�w�����Eȴ��\��G��x�;ʝ�����6�So��a��CA��= ��o�;]�%�AN)�uN��`��<�Wk0��_�����θ,�l��<J��{��-���~FPdp�'=O����F�ڨ���aiڑU*a�˟|�ve�R�(1�_�Rf�'��!0���M�D?����"����۔��c!{�����wຣ=��cy��3�J��=gR��t8S��T��z��އ�֠Ҝi��=����Xeb � �ǣ]�<?vh_[����n����O�h�����uW��KVE"�3c~n༮�ALS�X��55|�4#.��F湙�L*��pUy�0�g5��o��t��5L��*�ʿ�z�8��`!�8����;b�a������/B�n�M�]�'zNFnV��Z���X��-�w����T�Z��<<�͛� O	�#��ݸic뮻����v��7�n+SZ������c$�9��i�:E�!@�Y�H�~ʥ��������Pw��ßO��o3uE74�����
���4�#�z`���syԥsK�M�~ݺ�f��=�T��Ϊ�D���?�IsO������;�v~÷އa�3~����Ё��@�1�I~x�~�w���#�aW��#.�d�����X�%�u�քP�L'�;Oa��%-&�t���P��V�~T���va��k/�Ԧ�3]� y�+�'D�ѾM���P���R~����]�)�a&m�`<\��i{X��ijƜ�n)�ԉ�hm��$e=�T��${��12�����A�`���i�3�i��_Ii�sBY��:��t��z=�֬���~��1 ]�-Y���_$vO#�?�p^��!aT��ai�~[�nMN)5L�,7��L��q�{7]�����}�o��s�0�����+Ӹ�������2������o���˝�u۶�}k(8����L;v�ܝ�ۏc��̌��o�m�{_�g_�h�V���S�h�����dN���/7l`��'���9F����Ņr����T�^K=���ƭ�W�L��q�y�5���o ��2�������ä�	3,s�n*��2��Dյze	����/OI)�wޥK����u4#�L�p�9�G}��4��I��~����*�I�M�s����`<���h��yt�iZPt�E�"c��
y��S�/^�;�6\�!���<��7;��滁�6����.���a�-N�`��Sd��4Qh�O�o2Gf���t��b}������с���g,!Y̩r���k�Lc��μ�
;�w�����r9wI\a�x���É?pgg\�a�f�k�W��o�.���g,�v���Pj.��l�����^��-]�2��PZ����y_(�Q)*�V煑��-5�3)5ETn�>;	*l=A��O�`&i�K��L |�q\������0)�:�Tj����L���l{v�m�C�!`��iO{�'C�x!��0���`��.
�Â�Q��p��{Otl&SX�M���}�J���@{�E7u?�����m��`=��S0,ㅆ��t9�	'�KcXӾ��ǂ��&�x��F���G�����'�~2Q�.��'P�"*��o�Bm�ܫ�Lbr������^����.�ZZaF!^��9�aZ���L�)`�g̏�m�5�`(4ꇂC�p����Š����b�.��,7��L9n���`���my(���ܮ��\o� �Ei��V����+,�׮s�:� �V�gU��9�~y9��}�o(1x��s����NS�!���}�N���(W��y���:}�������|_����<<*��w����o����z��?��������i����7u�9���]y��5c�z������q/��55���h���	ј15 ������z���Ϛ�Ü_c4G�-郪��aXag�;�>)��J���]��.ŔC�7)����QX��۹"���#0���C��S�ev��k����4�Z�Q
�<�G02m�Oi���k��&��4G�U)\-,E�sRyA�yN�~.a�~��P�¤z(8��pbW
���>���1�;ǴQ��o�"; Z{���ۜ��$���Z�(8-#��;O�Q>S����`�U�Cz��ĭ���t�y&w<�$�&���7WPE�ք��YS5p���u�]���}�O˚v�~"&�nۚ
�||˩�h��rʁJe2mS|�R[f!���:*fn�ti��j���r m��J� rŎ�w�qj^�N'��Q�E���w�`���ur.a<�*g�7,o���O8�@�rh��=��Z���=�\������"�#���5�^�����iw���v��7�2�~O����mMM1�ad�К+�i�:3�m
����Q�v:V��°��^K~3�ך�0�x�&��o�����I�.��X!�2��j�	�S��W}s�6&�8��6ZN�,5��FD�rh�9vkf��<=�=�%����ECa3]�N�����)��6�\P�?�[[���H�.��jwӌ`�~�o�4�ā�.���o�~��d�
{�Pmc<����ۤ<��^���Q��I�_k֬}��2�S�#��k��Qu�m�[J
�G��C.)A��\������ /յ�__��g�ӟ�t�aL7��Hǚ>��C����Ī���z=�Va����od�e>){ε�@�rg���9P��s�̅��;��o'*�6�A8��0�j�]~Y[���f�0P�4�o.��֬Y�.����]
��D�g����KM��1�h�F���~����/�nk(Xj,����ߧ���c�Ða�q�pJ�U���,��^�P�:�*g�{}1s	
�-���ɯ�p�4��C R^+�ʃr"�������:��r��,5v<IK:3-o�ͳ���/�k�E��`:\�rbW
Ð�T+�A^�6Y?�L��1��r�̨�}����d����P<�q�e����R�����&�#����Nc��������a[*��'�?��P���c�>eE^��.���v��dפ�)"�'�m���m�ON��p�����)�x������rcNZ���l,���t?e|n*�.�56�m�t)Cߴp4;Y�4��Ũ�Ym��~��~���O�$�����ـ�O��Tϯh>`�Ǚ�Xa�Wwh����,����!u��7�҄O}�3N�if�Y�t~���k�[���v��w�k��)xj}|얟�}K��@��)i$��+_�J�����;kH��zk��{�o��o��nT 7	�_��l`gX��0�p�
*���i(覣�8��Le�s���󽔘RL|�NHR`)�ar#+�h�4	>�޹�OzB�5ҭu6C��\�^��W0��|�0���S���p�:��r���Ki�� �sL��w<��B�Q��-�H���S���&�8
[i�C�3�f1,�ڹu
~��OW�g[�C�_ �rS�=z
[ߊ���0<𻃶pj��ɟ���loy�[��j���Kh{��j�G)5��eucA�u81 �������)ک�g��"4w���͙sQ�b�@�mo{{.Dv9@1R�9s�~=���r"p_�hA�ŲV}
%�t�f��c&�~��l}ϐ�C:�^(�aR��2�q(�E>���$�#{͘Pt��[����ћo�9�����?��6�Ĝ6wv�����tɼPx�k�z���mwܕ�O+W�~��J�y��0Ӥ'f�p����/�[e�0TG8�kg�!Ü.�L`�i�M^�agJ�IyT���п��)F'��m)%��5r#5�n��7	��T<�昅v��#��xO0{�c'Ȥ)��J������X�	�3�:�z�P��SSK��,�u�?����ߴ0�}�;�3p�J+�N�^fn��[����:���)T��/W����9�B|�W��<~�r�!�]Q�ю(3��[��?��i!߸�Ҷa���
���_�Sd�i_O�Tx'�D�g�qR�š+V�̭��gظaC[�vM��항��E�n�}���_x�=��s����γr\z�}oظ!	���vLZd��/��	��ۊx_���◥l���Yu��״k��.�����紗)2e(�'�oax����[~�+M�
_����T���l�+np��l�U��zWe���d[u9����Y+�3����pŕ���.k+W�m��/$��-�U���_��3�1>���M)5�}J�1u�1�*L�I6��<�cp6iA��m�ϻ`�m��t~�`��8T����T\��QO ���
��ݝSFh����z&bB�"EP�G�a�o�'PŧԈ�7�����`��L��4,���^K��IL
=���8�"l�)�Ù�LA��8I�>�g����Y�_ء�4���	�4�[�H�W�;�%��z�A�W�GP�*�����k������`�)��IF�� V�Ev��(�(%h���W�mࠐ��=ߓS7s��ʩVК^"�w�ܑm�o�k
J���8
�|GSԑ6�����R��s�����۳�=�g]�ٻ�>x$�90����	����v�3���V��?�����=��7R!�򗿜7_����o�?����?��\\l�W����ܑ�Nd��Uvؒ1SCZ���XC��M�z�ڑ��ίd�:)�=�ې���T�Iη�;�w���N5�1s0Xӂ���8HKY��C;ui��p�tL9�M�����s�K ��Y���y��"��]zن�i�e!�C���t!Ἧ�17g����VN�
�?�G�(��Bc������l�?�x[zq6F��$'�UL�6�21C1������|��V���/�L�<&1uA��L���x ?���a.������ڽ�Z%u�$���(qQn#W�:��n�g�E��w�}�/)%� ;)hO�(�I߆0�\C�Li��L��$�q��P�%������p����1��OⳊ�	�3�y�|0E�Q���x��0c��|��߃p���:�ն<�IA���w���9R����O����ò���>�+a�.��Qz@X��t�N�޴qC{��ߞS�K�������A^K�S��?������?Ec_�3�J��3��+SA!�].i �c3Pپ}[*aK��~�<���f�+�4Z
�8(�g��9�����f�~�������G�G<GF=�
��TnJ�'~�'ڇ>�������O����R)Cg �!T=�S8�)@������;W�j�(�{)E�o�����œ�
']�{*�s�N)\�oiT:����9B,d.^�����'2�����('��-����~���\(8��m�����k�l���M�{��n����c��D�����aW0��b,��F��@��dht[4x�B�A���s�����ϔ��r���>���^���3ř��z����w�7�g5|�54�R���\���lT�]C�A�jpi8q��!��$�Ko�q��tn���L`&q_K�b�ש����OrC����7�l!�"]�S�N�ۤ�������x^�9)����$�8�ĳ�|�{�����.wYsU�x�Wf�����>6at����H��V��#�q��j��G�]o��]�|Y*G[�lm��}ߛr�2A�~���Q�9�Ú�
B��3��k,<��+[_�x�o�`��Ge뛩x<���!�7G>/� ���o_�)	_��N2�e���-6�D�RV�7���,��7ޘ}�-�>s��n�:�|]Nu9-yϞ�m�ҥ�ꠑ{�ȍ��Q��Ԡ;���:}�?q�S��/eFZ,�\#��p��$������K��]�ҥ�\4'��<O�OU�&ůt��i3%�Fھ�p	W4�'�~��䭧7onsf��+�����nݚ��M�^�V�Z;uK����	nW�6��p̜�$(�Sk��eC��T�*�B�|{ޘ��0d�!^�d�S�&��{����8�3�?���f��O�N�0�x<�FǪ�*���5�p3d�6��[��Ix��a�H�J��J��R�za�3x��!���Lr��f�r��1���o������
*�pE�OrS0��~���ff�q��ɾ�~��i��֡�پ�i��#7��CM.K8���x0lk@�{�M7������g�Y�ly*;��y�g��~��r-������moK<�vy�5׶�n�=ژ�k҂$mꎝ�ۗ�����/}1�,��-��핶5߷�W���^zyK��-����¾�^�|.�/���֋Q��^~9�F���!i _�z��'ڱ#G�뮽���-oIK����t���B$�>�����p���E�!C����ַ������|�Uz�Ν�.�dC�������w�����oεI7����=f�fw��in��t�؎4�F�#GV	'�=�k��YJ׬��[2�+��{:�u)P&�B�\�rE�t�J
�g)d���˜i���:G��W��<��kۺ�k�>�5�Z.�_@8o*T/������ ~�*cX!�]A�w:�o���2t��IG@X$��=����0�I �0N�.�!�ô&�{����ÍC�3���~�F�5�	�:q���g������d��4"~�X�g8_y�`rK�*eP�����d�0��A�q.������x��~�B��x��`���g�o��eXuQ��w7�J��U���sr=����l�pM����6`7��?����P) ��/9�Fh֞~��~�B1�:�G�فz���!��*�dɲ�b�6�J%�{���v�}����ۢ-�Zot`��T`^~iK۾mG�.{�H_w`���o��������+_k���g�'>���������O���������������ݱy���p(�;(u�]�.-2w�yg����s�rZ�ȑ�zPt):��
��Khqq(1�x�;����ϴ��W�j{�����/�k<�����}����7���h����~�����O�D��������g�����������C��|;��Cw�;|S����S����>�B��p./�z^�D���F�;�W��er%ő�"
JWv|�<u�����L��x9w��n�&�Պ�%'�3$.0�7�f
�2UDi�&W��1iF�Vn�#+��PֿI�����
�U ��~�W����d�Q�b|t�9D�����c9P��+��d����0ޠ������C(�x/�����&�4�~�2�G^ꗠΑD�6�Z���{��t�	��2�u]y �~��|������8L�?�7E�@��Q�t����_|5���v�]�0���8�a0H�B�T�:����]�g�X�w�m'�����0������t�9	�w����'d{;~�k�ɤ'A��+�_����/|�}�c��e��~/����'?�kx��~���ӊ	���b]�+寴~��9�ca.�x���?�6���kӲ���(S��8�޽�=��#�djv%����E��=���m��}m������Łۂ6w��6���DY�9!Cŷ�E��Ӊž;��]����n[��Cu�ؑ��u��ӥ�,Z�(�f���t�=o��ѭ�Q���Rʤ�U�}���:��n��yW(4����Tlrg�;�XS�P��m��K�������?�#y��K^.Ӆ������Y�`��<;��\�pq�kw-����n^��J��\_4on�uQ��c�||n�@Bg$�Z�-����Ѽy�z�h{��	�8�yPl,�����G�軏��g��9]Pn����GR9]�9Y�	�e�GP�@Eak"R�Ie�$�>	T|1�ԙq���^\���&�0+pv4�Y�_�i�y���C��b0�탫W��0s	�
G�F�E�em��x��3/\���{�+eO��,�b�/���ʎJ�ba�uQ��@���nH;��`X�hUuwj^x����W)a={i�{�ܕW���^�~�'��c
�h��zx=��F��ʝ%��tlC=�?@$M�oIZ��~N���SG�c�����������m����?���a�����~�?��?J�Fx�X��Yb��o����>���������N�0�����"�HZ��LՐ�p|y��9%�SO�W�E���i�����L8�Lq�yi���պ��w�7���u��펴��Z����%�nd���|u�A��P<��sv.��C�Z SFγ�����2��w��]�am�i$V*�kVv��w������ǃ��f^�CkvXնlqۑ\S�w�+�O��:�8z�cJ��.���>��$�#k�����u�u�z��3?�p�®�/X�Mi����o�<
�z:��(�l�آPZ.j/��r۵�%���"�螏D}QTNׯ����q����TQ$)I�����.@}�ȫ��������K�<�3F_$Z���(աW{
z冰?�U�Ҭoe �ŭ�z�Y��V�K.��ojT)�x	k��B�8���'�j(+W�Hӧ�L=	��%4 �%JXI�g.�h�)�og���5"�ߜ��	Sʍ4������ӦC�2��U�ql���x��W��);����f� ��LV�=����˞���ך�q_kYF����[.��>�g:߁:�&��قN�Q������w���O��/�f#7�8kN�ϐti]��ɣ�H�)mA�Qޔu��t�9`ZGgY����<�`�+�x�)X�!�F|�h?�C?��n�ƈ^�9�(�˛\�T팟��ݮ��P����.���T}�wO(@��������������z����v�wf8�?�����ko{��R>s֡|��?�����j��c�,�t��O�����Iꔭ�!_���z(Q�F�!W��{\~Li[�� ��n�-�E�>�������k"�7dy��I��/�����?h��;�����G�=���F]�㟼����jS'Y��K�N
���;���RQl��2H��Q� Ws�.Ӑ~�m6�c�&.4/]�ʋ�$x�i�GE��c;��l�?�b{�����[PߡD5|��T���G~�મ��?�*��o�<�/��;�c��:d.̀�t�+�� ���T~�)<�W��NaP��(9�,h$n�]B�o+��{(*c=��]`23���탇�`�h_���ݻ�}m�h$��,�RgݩȪĎϬ�}�8f��3CZ���v�m�w�]w���[�=����ʤ<�(���/+tZtWP�Y_#~ �T��x��R��z����s�s
��A��)�;�EH� �0�\c��)�ٖ�����F�A<|2��s��$�9�ǁ�������?~4�!�BV	9���E�ےJec��d��l��p��M:)�)��)�Z����u��]r�U�B�}��}_���F��2t�C���ƻR��p}
\�%[��mg�W\��s��Q@R���|B#�7乲�I�W^ْxQdL��(PL�Y�s�ͷ���w�5�%.�2�����K����og��E�}���\�aJ[�D0Y��	ʑ4��m�	����Sq��ƛەW^��S6X�~��~���������y������ņ,�SՁ�����l"�o���v�e��./���������=�ioy�[r�=g�ڽ�ܛ����v߽������y��7ef���������������`���}�C?�>����{�{��?�����/�y{���7�w��������nz�ڍ�_���������ۇ?���zG����rv%��[~���r)�h��,[vqд�I����B�y�вF��Qb�b6��h��N��D�@<1)FPɜF�����K�T(���05 ɻ�#��\�[醶I�0��U4X���Nx�'&̟���su��"�.�N����Dz�H�EhhS]O�d���h�dfϙݮ����>�Ly�}��y<p�7�$�FCR������u�Aâ�$��t�fn�0]Z�D8fb�.Wǈ��#�'Z;���y�3�#��Q�mm��m��\��qg���{<-��M��};�6��5G�¬��|����6��xJ#��2�Y@��Z�q���t���=��������*�x��_���\�xٍzA�,�#�4���� ���E������NV�Wr�x�GIU4�=I�r��\�n}�N��h�3v'9�<��ˀJ�e��<� ��t��Ȭ� _���u�W���Dޚ~�嗷B��|-D� Y~�WW�oa��C&�&r���ݡ�Ρ9���ٵG�r,���]��:s�3��l�7d�JuH�I�����S��7�UƗ���y�
��H����_�~#��n��~_ܾ��w����S~h��v?��pE��K������������>�~�w7�{4�
����O�ٻgo����甡�z����&� S@��ଌ@� /���Ⱦ��o�A/�wF�)|}7Ս����h�ǀ��w�����o9����Pvn����j��n��K�7�+�r������n�5��.o.Y}��ƫەWl
%��v��W�;b��|C�������
ӽ�O�Ӯ�ꊶ/���6��>�Z|���g����c�`�F��"����؀6��_��/��酄�~M��i1�Jż��ձ[T�3����5\�CA����<H��������bq�Zm���*-��)��@t�k�����ʾ�h �C��.W���-���bi������{�-�ߜ��M�o���k�Ά}���#��m��ݩ�h�Ǐ����� �ͳ�T֮��}�>�+�o����Y�Ey=��z�-Yn-_���t��\��s;��f�POӅ�I��
)�Bh�6�`TcT�J�����^H��*c��T�6TB�R��ƕq��hS�Z�8o��ג�03���*Z|��4��iQ&�87�/����8��T83�}IN�s����װ�Fe�����%���G�5\�x:�S���8��`���7�0D*�n�-Y�.y�!����k��Y�:wNҟB����p�9��I�!���i��������Tm�!�(-dF)Z�꒝v9�+ �%�D�{���e� �|���϶>K���D�T�}#k�ӆu��-b�]��|硇_�+`��-7ߒ�N�GC��-�����d`e������Tn���>�ϴW�mɭ��g�'�ڻr����<<�4�>�#%ñ�����rQ
�L��C���Q�KY��]\���p&�X
��;wmσՓ����+B�ߖ+�J�<y�-�Ո��k�e�u�W$mfŃ���ꫯzo�ߦ��uW^qe�:���G�5k��W�_vYN;��d}[�zU[��|Ų�zm�/�����ٶ��|;�W��Y��-
�Z�.�bc�;:࢐�Kۆ��íi�6]JJ��(�g>��6g�����Q��۳�<�$�VRlքR�o]�tq[�nC��ڠ�[�&��s�]��<\�Q5L�S?�S�eN��喛C�)�_T"�1/�2퟿��;R����7e����=���d@��P|��P�>��뮿���m������l�����{�t{{���;FF�	%��v�=�ŷo?�S?Ҿ���i�����������F��m�ȇ��w�_�o����1�5R`�%�)�H��OCU�ʄ���؁a����� � Y'֯o?��?�g-[���ڹ+���3��ϸ;נ\A	O4A;#��x�xI%f
/�á�8���$(^+�����o<�˝�e�o��7n�)��0F���-���hނ\Ӱ*�;z0���n0�p�'���A���q&Pc��r����&Aś��2��8]�3� �m���RW>�n�������a�Lu�8x��;�����w�+��N�<[�Շ��}�g[�h�K-|N�V�Y�᩾(�kW[!���0>�	��ڇ~�S���K�vX �ΰ z9t�x�+8㥶;��Anu),���x7��S��g�r�����k%Yn"i��󏗴�P��N6+;�Y_X�>��?��й��LP�h�������D�<};��4�Cɗ!/�����|�0��Y�����P�w؟Cd�&����سgw��a�������M�?���\��>��x���s�o��:�zy���L[�l��Ѩ��K�GZK��@{e�m��W��Q_G��=�vD�GB�X��?�O����������b{�Gڳ����K�xı0شҬ�ڄ?��8����l}���L��%���R�`\��`���7}d��a^��Ix�9��3q�� Ki*汫 ���Y�!���.��ceA�#��E�6����/����h�ȶk���_�Bۼ��` s�vtSb�@�gvj�,L��Q�L��������ӚZ�o�B�X�O�Ј	����7B�<,acT���6��?ϢKA�w�}�)Lg���S�\�N�:<��CCv��÷쌪x� �	�=�7rG����CڕW=�ӛ΍�龏�Oz�M�JX��#�'b���'��P�뒶 ���N�6"�.�9$��W^���G�rF��A��ۍ1Pȋ�B M�gO90�]�L�J�|�ҟ��w�B���e�ciM����x����F��9�^�	�>s���V\��-���f����{�i��������v{��g������]{ڵW_�B�ݳ/���v"�G`�iΜ| �ՁQ^(�d�0M~Y��M3�:���%��T����o��o�/}�K�t��۶nK�K���n��Q:cW%�G��9�`=��an�ֶ\��GM�X(˒m�9��P�XW�M���ZdJY��#�n,V�O�ә'y&/���,ס�垢��e����.������?�qA�,pr����|�K_NEI\�b���!�+K��� x�v+ձ��o��F?����_{}�eeEg��zLiY@{�=oJG^9|�%�S�I�x����	��A�텓�:!������s��P��\[�mM�؉��jo8���n�o�w�h�w�����z�ub�>6��������O�g�{�=�'�x,wr%�U�n�W^��>��/Dٗ�"�.��=�W����p�A�w�a�%��W�5���R��������Ԩ��1��7�cDJ���KME���j͍w��b��.�#�%�I��
�=���i�4���o3��y��N�ǟ��i�{"��R8���o�}��`���|��\]�`�s�}������^���/������Ov
ʡ<FT���ߛ1f����0/m����/'��K(%��Plh������abith	� ���tP�n:�l���z�S�����>NN�&�2RP !�W;a�-���h��;��E8dx��B�=���'}���y- �j�#]��W]����=�Ӝ��.��[߮�vg��c�+���ڲ�Kە�_��ǈ:�\1��������n�G��ӔcX>o���Uj
�o"x{���F�o�)����$7i�'�_

�O>l�Nz���s�i��ui����>ݞ~vstDG�.^yek���k��5k�����v<;�ay����M�;�f����`�L=���"+�ac�ٴc�����<�H�ַ��
YA���d�W\�mȎ�/|��yϞ��3�凜юt����D����S��U��n=0�Cv��M�`i�Ԡ�-�v�'{�LG�g)>W]}U�5s�Sa���
|dx��/�ɾ��h`I1���SQ6��z���wޙ~d��,��Z ��޵AxS���i#t�L�4��6��#H[��:c7���b@�M>}ҟ|�O��ڥx������<૏�L=����Ii�ʑ�k_����Ϻ(���F8}��DX���կ�©��b���>}���ڟ�m�S����}���o}'��ۃ�~8���>�X{�.��.Y�!xbE�u|v۳�`(�_�4�-_�"x �Ы�TjN�)�yŲ��M�ϗG��Iom�λ���0|1��, ����1�Ƙr4�h�ջ�R�~k���D�8J����f�?�ր�������χ2��Ï��a��i�.��d:�����E�/c�`{�u�3J���b�v�5i�����D[�QG������l�0.��������(^̱5�M�בI�Ӏ84������ʬGI�o�k��?t��s���_=�A/�weR?ʮ�6�����O�����Ba�ך�����|:=�ya�7��ti��<=��lJ���J�\Y��>��λ���X(�[^~%�����{��[o�����oLMX��7F�.%45����ЍOW�Ie�����u*T賍7	�0�zH�1?�~|���s�N��k��Z8;Ś��!��b����i��_�\H�!��V��v��>�X��8_��l�2P�Ms�R#<�ǯ:Cq()�v��i*2�Φ(O=�T��������à�e�R��7�%��� �m��c:���O:�_l�˃�y0�Q:
G��\۶����c����0�����ze�+)�o��-7����r%]�BC��>��@�ZG������[ra��٦�%�P�<-����(R��w���������w�d��P��I� �M���#,�Ж1�w�����(���?��e��H�K��z�+��+ٗQ����C�y(�E�}u�-}��.�����������7�fۺek��Em�K�ڟ�ɟ�/�k�'�F��L��S!S�mO>a�����b,_�ֶ��3�˭7��KB��L�����B`��K�кTT?��9sg�ի�ҽ�m�xY(��~X�F���%�!��;�a��t�em��������|14L�)4U�:u��(0�L�vY�Rc��*�����/��/S�qT��`��B�y0���s���s���X����?Ӟ��B4����=������ǎɵ+��h+W�l��Í�+s�9u`�SG���|:˥�+��u���\�Ԉ�����F�	�i; �yy����p6N䵀��&�.���]>���'�O�{2��$��pa09�Ix��|u�k�1�FC2���rԡ}�7�$>�'�	ճ�O�p�:�/WP��À*��w��V�a�X$����+w�(�_~Y�$F��RW�Pݱmg(����8:"a�oﾠ��v��+5�-:�=��=Ί�YJwX�*�8���E��K�@䔺)�֘1��j�a�U^N��cڮv�o�]��������ۉ��S�-Ιێ�ã�Gx$�
�qt����P��kp�eEg���ȳz ���Yt�!?L���!W�w )�w�+<��@���7<f����`,]�I�4�a��y��b��k�4��܍Ƶq��7����i�?������ ����P^�[�Y�� ;�GγZ��.�c��"�|��OP.���N"ZGq�6ʡ[�L<��eAWʠ#?(��.�����o����}���7-Y��e�"�?��?I���M�{�����V��T�v�r+��E;���K��p?��}��Q_�)|����_��Q�E��7�/�����.�5�͝��~��%�����<
�'��{�-��,J�"�¨����K#��wm�pm�mk���v`o����Y�H��z^�~m[�ry[8n�wxu�����ൠk��Z���c5��	i�e�Q��Ԍ��JT)*?	6���[���������Q3�K���?*b�Rs�� �7{v���7��~���C۽so[�`iߚ��7��>��i�i����u�����^�zm*1��$��$F�����f��)q�i6V�g[s�x+��e����}?&�-�����m�x��&�$C�S�6�p��T��p%�4����-��K}�v���3|"ɄZ������.2+��9B@��H`J7��?��n�4?�U����s���Fp:�I��������ehK�Y\��O�,�|�U���t��d˶W��f?�.=~�>l��m^����e/mBٙm`G��'�z:�6G��y9��\��&�9L�efR�q8ӷrCA�~Q��׌�L��!���`Bt@۶ni7�x}�":��A��{w����֮YѮ�����x۹kG��УTOu����x��SO=�~����w���������i���>ײ�pn,s�w"�vU�)���ݚ�K�1�-˕�I��O�D��G>��?,(��qFt�sЅ��6\�i�gݍ�Ý�,�%G�l����},*���;�Wc������Y;(��G��������Ǐ�h��,Y|8F�y?\�O�pH�Ν�ҡnŊ�iA�v�ؖV3e#�)��E߂�o�D��PV
�yu���7��-��PV���_��W۟}�10vN��v�5׵����yʰ0�B��F�3�9'�-<��*ñ`i�x��G:W^�څ��F�����/u;;x�9:!O�^6;q���
�?�����s��j�b��>�p7S��"v�J�5;𚓽V�q��F3�ġ6��p�B��m��痯r��P����t(����Q��u�S���w��s�9��Ь�˯��@��;��/Nvf�yv+?�$��4�KOC�G��u<�.��L`N�� U���{���Y��?�S����n�����v�nJ͟002��4s���o��v���P��ȏp���ʠ\�������^�ێ��ŴE����f��]@�!ȳ�����C/#}#=�K��Սt�������(Wm8�۳�I#
^�� qY��_�;~�銫�V�.�V�HѴ��{��,֔�o��,�w������ݖ���^z٥y�-<��ue��YN]��{M���o�xx︟��z@UpPB/�;��۾��ꢵ�<���/����-^��B��{C0>��w���۳�tF)�B�ٳ��HK�A���͓x�L0,��ӹ!���=���龁��
sJc��ġPנ�[�f��W��G�n{���ۻ�������kWn������x*9}�[18{:�IP
����TUXg�2��aZ�7~�7���}4��xN���i3�R��Q@�>�O	�Ϟ�����b$y�H�d$]w�b�����u��c-�֭�:E|��9Ѷ��`���G�v��#�<Ma�:�Jα�H�S�yw���쇡����G����	�1��b`�N�?�^QZ�G��I8iL��F�R�N�ޞ�g��|� ���/�&?�K�E�D���{�'?���k��k�+����ֿE�~~փ������>�OE�hM�`��N��>��1h*��F��t�ڡ���7u�H��ٳ��.�����8��PC"���]�Y�ۢ݇��8�D���E��3ԡH+�E=�8O�}���9����P��67�U��nl�.Y2*p
��uE�.���E����S����t.��'�(�N̓�)���y��+Ta�`��� �-�(���[�.;V���T���&�=y�_�(+��l��@����m�|�����3��t�vg�97mL�߱#:�=R��M����/��'��L�Ԝ��-&6��T,��)K�xRj"8�}aQ��]s�:|��T�h�D:�s*��acư E����w�ޮ���v��Kڦ��� (�/o���%��{ސ�O������T������p��w�bqCҌ�ɩ�q�{4&;vlE�����:��.�~&�չXO��F9�2�n����X�;�ʈ���o�
~R��r��r�!�<6�_>�'��o�T�CWi�O��������ݶ��R��а�ɂuJ����ly���rjĨlk�?�e[��;O=�t������^K
�I.����9�>�^n�m|'��y�����{�wz��m��U���n��� );���H��Ĉ�Ѽ>��!���Rq�J�k��W\��)/��F�d˃�;_�~2�7e��{���7��;Sq�f?�)�N�pB1Yr�]o��n箝�4=��)�6nؘʍ�Y+L�A���<���\���Wfyv�lc��%�lHň�ŗ�˓�Cޓ��M�܇�).q9JCN���e2p�*�5�es��O=�w�y�2����3Oo��� e��d&�K&�\&~��ճ��]�Z*@��g}��k�,��o,���|�2-�������n�2�u-�܅C;�����=��eү8֚JZ�:aN��z;��NZp�ײ��N*���`�2��f];Pݗ��kz�hȌxS�C1A�|ɼ���%K]S1����-^��]��I���>rk���"y�=��4�پi�m��5m�sj�$.���.�\E��x�e�U���)-z��D��T��D|��y�tOP���0�ri�:}yf�c�C'K�/��ܾ=��ѡ^����*�_�lj�N`�dÆ蠣��w(���m˶�B����Ny |(3FOF=Ui�Y[��[X����k��cP�RpB(e���"+޽�@��Nq��˻zА4�R�����BB4�d��moK��0�!w�=w�)��;o�-���{O��B��.Ҹ7I�vz��7E�ZҾ��ŇOw+P��S�Z��G>��τ�:�g?`���P�(-�NI����Gx�_�4���>P^4Wft+��`��g(�E��(��c��uM�V�¿8%�QT�n��X�~1����H�v�h�%���A�F嗷l���/;ہ��tF|�wmO{aN~����ϑ�7	�߆���g
���L0_��,�S��E�I������F�Qcm�Ǟ|�=rmo(�Le'�ޓKRi�'r
�u�Z;��7�KFZ����R���O~*��Cx@�(�mܗ]�)�YH�$�lQ�m�X�e����yvs�X��|����/�0�@my��@L���%��?�+��YJ�����;Ύ%W584p�&~�����oMĳ.�"h���l�8E?������u���$��omW�\p�:����{�dJ,������hZ�II��/E-��E2p�x��ڟ��'F�l��V>�G�zOu�Fc�] c�Gq�X���9w����ߟ'�+ܔA�h���?�D�sC�0Eh���N<��d9y� =
�����8NV�
ӂ��-�f~(&'B�Y���vI(+�w�h�<�H{9Ti�j)���sښ����4�{S[�2��(G����q��[j4L����  �5��Z�����B[����dP�xfE�U+��t���xfUi�S��Z�_�M������ħ��Z�qSh<}��ܲ�a��\վk���j;r�hV$�	�;vEe�|5 L_�b7�^s͵)�X{0���|���ބ��)GK����o��d�/�Kɸ�ZZG1y=�Ç+�5���~���4KS:��wf8�Z��U��K�1c��W]*���7:.Z4�-��1���7�������=wߕ�&^s��m��[��I�G
����k��NX�cq]_���i ��	�0���"�k�Ki�x�hXt:<�|���9�h:���k�S:<����Y(]F儿�+�^��F�U��޻��	�/%rV��.h2;��m}ek(?Q��W*��	E�r�`�[����.�$8S����o,��d�pʑ�g���~���¾u�/��^�B?:��=�G�xOd�I�q�wu�Q��aħ>����
���g$�O���h)"�zX���ۦ|𔎌�$����O�w��]�O�q̧?����ɶ'�Ǉ`�~���]_���7b��� �$�BAY��*@������]�X
@	"o(A� e����e���`:yV|2����k�I%����V*ڎ]9�]~i{�o�zQx(6���eH�����oSmL��=E;�l(d���+[�J�ܳ�$�F$�=R�+]xq,W�|��.��G���M۾����O��O��C�x6h���E?Vd�):���L:7~�=Y�i":�*�L�,����Q v2>t�͝57�E((�ND�,m�.Y
�M	���ek�����<������B�
"�PD��vY��u��5�Rj��j��fa�k�$��h�*Ú5�Јi�����lh*ނ�������~4OVQ��I#ڶmk0��d��s2J)A�D�~FX�D:,� ��h0v��|0:��3������i�>�T����ͷ������lǏ�j�?�x{<:M��[���!�Q��+�?��0P�00�&���Hʉ1<�#�r�F���S����^��_���hQ8zO*5�3l�������7����#޿���>�i�hD������k��l����,�U~���K�VG�=	��{v��$��6%�b6��i�+Z�3;�h��p�1���~`�Q %������� �Pg�HW} � u�<�~��I;D�j���#�4R�*#?#Xu�^��`���|���׮��,0�>���x_�4�,�4�ѝf�_qY�tݿg_ޯE}u�9t�h��[&#ր�t��E�$��>3aOo�/7�⢳r>�_g�_)�������N~>2��9|D]R��{�_e�?��B?Z�u�v����(�]>ޗ�k��u���_J��;������|��a�#w��K+���_��W��L+���4�����Pb�U��"�6(Ͼ�@~��9g��E�.�JF�iy=M(.�Ծ��*�0���L@O���V��A9Z��Om�N303 ��_�������e{]�a�/��>�o�E;�1 �Z�Ģ�	Cf�|H�:�:���~&�=��w�d�G�����7^�����Ƀ�cǮcZ2FY\���B{}�Z�n��]��'�(�[2�����X�Cɂ���E���կ�=��S���m�E���H����}����/�:��m�
�������������߶�|�3��d�,�m����w�u���p=��mm���Q��Nmf�λR�))1��0����N�����_ڟ}���4ɋ���&@%Z0�A�v=�BT�·r��ўK��*N�/ͿFևh�̌̉�3�G��tɲ`��!,�m��mkW\�ҷ�v�_�׿ٶ����k׬
��\��̳�cN�c6�����9�X4(���V�%@�ա� 4t�����y���,s��=�^}�{�b�����M�K]�����SiM+N@��;�����`�ݒ��V��0ʵ$�9q7�N8N��IN
��nW�֬^��pZa�b�d�7����܅:�|�F,NZ�B�u�����`�������`�������JƦ.�����B�rGx�7]�p����Ҳe�A�'�'�ӿI�&X;��b���|��t����n�uA�Ƀ)�u:[c�����-SG#N��CG�ˮ�<pt����v�=��(p�S���m��,�[�Xd:��$��U��}R����*���?�{=0Le�ay ��� u��iӨ���m���u��x^�wG���hˑXZ�T��=�/�/�E��jG�2-�=�Y�3��0�w?�K�N�&^c!������9��p���?�����SO�̡�@�[�F�!��@RF����fmK��Tj�N�D�-�l������p��������ڜ�M�(S�e1���A�uL:h �a2�� ��`� %�e�87ӳ��7B�y�Rm��}����]��"��D4��Zv~��=�y�\���x�����ڵ�]����cs������˽>��K.�J���8ιa�w��~=��Xޮ�Ny3�#o�Rr�bi�=�R���ٟ$o���N�����]D>,=Q�T�k����kOY*p(��6�?|0�e�����pU۽�p{�����lm�\|�9y��_��g�%x֬#m���[�rO�xɺ������Qj.��{5���TC��Ѱ`%ch��
bk��&:1���r]D�}[��AL��7�j��uy��5+�@�|9'�/��(Eg�~��d��X4��+/n����ٷ?:�/c?�#�[*�A��*��D�-]fRe�����G#�(8j�]@X��)2���chr\�q����ʟّ�5Eg��Æ�9Q҈բ`��V�^���1?���<fl
��o���/<��ݯlٚ��y7�|&�O<�q�(�SO?��CY���!13K2��f�/^|��<5u�>���'��{K(Y*�9�Ȋ��#-�{:��2����# ���	�մ��o���V.R�0�ɓ2Lȗ0D�Iu����[�w<��.ă㋑>�0�<��\.��A�->v$���+��jφ�m*u��um���i�&#�t�<_T�ʕߤ2��!��U:�~��8�y��U�Յ�ՙ��?=|�%G�̽ؽ��'�$�����J�ʩ��M����Av���.-��~��^A��*��O"cY��� Sk,�V��6�>��_{�u������T�e9tuGvGf�+ָ�����{�v�7���7ޙ7Tk��g����;�m-�݌��GSU�|I�S���9`�>%ek(K� ׇ6Hq8���h:x ���@�B����S{��M���h�dj�@������p�*k�V�l�������G,W�Mvղ\Ę�7��B`�ҿ�K�#Y��,D�^_�tq�t��CkEY/^�4�5�:�|L:�,Q�X"��,��a0h'�\����nj�.��׶m��׾��>��@���=�ʬ�1�E��>~^NY�7DqIs�Epb�:b��D��I ^5BJ�Q��Ri4y�.!+0��.���h�����?��ڵ^&7��,�d�sK��݊�(�[�G� ���טK���q�_wI�Cm��i�]������8�n���wݺu$�a��`�,/�t|F5F.@��(=ۃq).�)�Q�O<Z����U@']t��]\�x��`�#ZWD��,U�A���b�П�}��U)��f�ܪ�@��_�җ���ܳm�K[�L�b!�Q�y�_��^z��\�WZ<�\{���Cٚ�+����RH��oN�b7i��+/���X ���ؐ��3z4�#4����[Jk�*Ŧ�Fo8S�ԇ�m����0�F������.�W]KC'�f궄�8��aXC���Җ���TՁ55��sϽ�G� ���:�Z�"��\��E1j{���/��#��Cn��2��x�*�L�m<L}����8��a��^�S��$赽���?��[�z�＄5ㅟ��C�)��������(�tu匒�H��9ĥ�d:���ɐ����G�dg�ys��A���+���~��xߖ����1(qx�v��3����|7}f #M��~���/i����Cr��Td�4�t��b��7�ឡ�/����%Da�`��!/�x�����G�G�O!�Li[�����4�k~��>� �(�,���Y���#��a�g��ŋ��.
2�J"��Ƀ��Sx�3��@��B�Ģ;��n�%e�ylz�,�����ׇ̾'*�S�ǂ�D�7���v�UW���>�U��?Z\�NV6�6d݄�~�H�R�"���n�:�d�Y�ϡ��υ���|E.h͟gJ�E*d؆K�]�֮^�.^aG�G� �]������1cjf:�s�jU��*9�D�F<}�)��5T��xM��*0§�NG��;s:z��L����kw���`�ۮ=;��E�C[_
������m��}���`n�˾(WgFV�4�bxyQ�4l�����Y��);%FGi^բ����Cίj��u��DQ��e�?.��}�7��7���4�n�����"���8�ܴ�+�/Y֞z⩼#d�6��B�7���6o͋�	&`u�Yb݁ka͛���~V�Q�9_W��c�@Y't�h�~]��UW�H���oh���'��g���)�$X���N���h������������6*��P�~��<������?�Va�:�n
���Wu���R�g(ϗŨX�pJ�3�oE(b�1�qn���T~uF�B�J�� x�P���l��.^�{���w:l�<I���dô�S�R"����Ge��H��_)��%�#LF8���OA�}:��m(ʍC���U��n��������E����~�}��_ȵ����O�?��?KYd �E�3���n=����p:rK�O~�������n��R���\cc��t)K�)g�|�k_���?��?k���\S�� ed�8��������s=���p���>�?
/oe�>N#�d5��RC6}��ᦜʠ]�JS���d�E�d�EIs��������*j!帾�R#E:d�0kN��ݒ���Di�+�6���ƾs���C�k��&��ї=��3���<9f�X�M�A�p>4��	+�Q��;�����!�V��j~(���W��`�s�5ZD��=`�r�f�	��5��K7�1 ]�f][���`�hct?�pz�| � J�
"�1e�7�*X��^9��;:�ڗ�&m��u@��dT����7ׯ�Nr^t|�Gf�eIp�h��cJ��2���]��I�HK6i
���R�R�-kv��ۈ�PƜ�@9(F/���^��_����}��~����o�Y+�K��K�F�c�X.p�Ǉw+ Fא4pr�ZL�<O%̀8pF�	�?%���Y0�2��J1��,]vq���Y�p0���A����;.�5�`S4YI�<(1����3�cJ.pr*%e3;�H�cJ
s�s{(�K#��WG.����]]{���٬��_��=���j�����-F�=<�?���5�@��/�O��»�?�o��PiI[}k���TN�/��ZHJ��T.C��/hj]�#�%���E}�9\_�m|��K���@y'ю���:�̡J�9�
����<�{��%d��I�=H�d�������9	��7����7�oc6%ѭ��R�X���c� y9-6/Ġ�m�:mS�d���P8#uJ7�H޲:��㕍<X�O�|�ĠЉ�{"�]��1��Zv�d?+�ۥ��V�Ky�ʖ~���1�,�6�Y��� �!�8t
�@���]�i�=Ki�4 ��_�� I�������p�O�`V����dȖ�$��K��S5����iW�G�`A���2`R7�bʙxߎZ��K���6x�0Sr��f�MN%fi� ����M�<_bGk(R*GLW��=?S�G�E�<8��(F��..��F����Ϗ2tk�� /TK����OiU�T>��b*C0ϸ��,: ��RV�Zs�]�uҢ�NĈ^���\^�u�%�<��n���f����yd�q�f�v<'�bX�50J�>��-F�WLc����T]��Rl�f�qS�#��Egv":���C�BH��j p)��)��O�t�E4�B̌�i�:,�������������1�K�W�x^��!~��հ�KxZeu�M�)�o��
��дƾE��;�lo�;S���7F]M��[�G>��=����o������L����h�WF�c��GP�;���9s�rrX������ 	L�s����,A�B0}R>�p���Gi��̢b��<�9u�r��VJ�0���X���h\���@���\�O)R��ßLr�����S#���iP��&�����?�: ��no�%�~� �6�ko��>�8��~w�-W0����^������:��'>�<{;�tF��K	��~V����7��q�?�0l��^���z'<U�^�&:(�����o�:�u������*��O��92�����'��ε�s/������k�P}"��'E��!}����c�Hִ	���겤��R8��Rf�睜�� V�HQ$|�ؠ����uTx�BU�o�A^V���E��5�{��"���3�J��5L}7*˭���"m�G6R,X�է�O����&ҽ8�\Ұ �E'�	
g�����=��d�;��D��G�`W{)��{ty���4���2�'W�M���W/&�ɵ� L��R;�ζ�F�8:v̦�ҁ^s�59E�h�����+��溡]�~U۴�vy(7�w��N@Ŋ�V��GCV��V�J��y?�� �ߋ�玗���G��<��w�־XN��gPDc�o�T�̫�h�l������@�YQ~�Q� ���~��2�_�+%�@��Pp~4ޯ��(Ko<�@��s��3����ј4�)3:n
T=�L%��Np[ �0�'�q焙严K7�����ʵ9#�t睷��9'b���+��Xcf�d�A�A�ڠ�B��V,w��Y��΋���v�����nM��W���E�i$]eS7��
LӞ�i�'���������o�V�^;n'�a�P�ާ��I0]����Y�aC��#�&~eڎ�v�f��'BI�0���_�;�o���85����gA�Q"ڠ;��CG���cqS�6.I�u.�pŧg�¼s�4 �q7�2tS~��;�nT�q:�k@����H��*Q���ǎ�h.��9ʂ�ᛴ��۳����9eS�^VOiUz~�D}����'9}��gW�:ﻣ��Γ"#�/��<?S���)���\t-����Oa8��N�T��%p�F�b���LN�5�dU��%h�~�Rj�tg�����.S�؄����)�kOea��l��oڍ��^_lݧ�9�ѕe�f
�9��t�'��Ż��o���P~��ݻ�?i,k.E���{��˅��8'�eم�hm��OY'�; ���9N�.e�yǼ%� H@��Au0@E�@\�UPqT6e��`��M7����<Bڔ���+���|
bΎ�w��:(�#n�ݢ_��tV���b��J��V�ʱ��n�������|):f�c�E�s.
�Ƃ�����,�ƥ��J�������VHʉ^�Fc1���֬X�K�����}'����r���ܲۅP_LZt�F�^㮾;?�����4�.}uA��(�UrV�k��Cs7Z(�g��5kbh����;�#~/N3.KAa��lLǟ�̧����~��s���g�R���1m*����b7�6���t���`!:k��+//P��3�A;V��}� �s�،�J0U��#�^����T� �����d���괯���B�խM: ItE��v�� ��=�
��p��(2�b��/�B���C���K&r��_�k-��Sf�
�8�K�F�]D������_z��e �Lrc�g�B��G�2���)7)�	~��f�>�ʱ���m�I��7�h���	7Lo��Rw�3��~'�U���΢ح��}�8�ig	��:Zm�)�=n|����IKH�����!���xN�_r�?A&�������~��NymB�)Gx�㕿�]Y K�)���T�E�V���D�����y�E���"B�0���^x1�8>����_�r���?Ӿ���)����:����c�c�i�u��@?Mw5�@��u=6&>������u|䈻��#6��A4�2Q�/Y�/��t_]�F����[&�a��	����."̊FR��Yģ�Цu�v$q̀��:��&���o��:x5��V�Z�6nؔ���H�%�p�T�X�k�/��e�b�n�y:�3p����)�S#�������9J�7�(Q�O�6���g�j����:X���I����
�p�B��������8tpA��t�@��Z�/�'�@���wu��|�IvIЙ�,�/@c�̇?��w���Y���7������8o���o	e�"6e�z7b���ͷk,�SJ��=�������I��.�E�����z�Q�/�*��X� �OY����/�I�K�gX�=F���0���~���Sڎo�f
NI#������*�)���S6�p�?:K��b˼� �dX���.5k�	�*�LVI�n5S�x�N�hxa���V�������g�*�S�8�;L��f�Яx��$z�
�,�@�-�A�:�oøC�$��@��&5��5|�7�׮��X����t \�!��Qnm��w�\��x�)�W�O.m�L��n��ȍ���F��Rbב���`�B�@SK��"10X s����Ҧl���[���F�m�p/�A���ձ�ͩ��;�R�پ#���p��sbpr6�K;v� 6�2��+�X��7��!�]T��t
��"r���fE֬Y��$���L�/,h���0Ɣ:3�(Ÿ)(��󂲨0�E?�vC*.�����i<�.q�#��De�h��t1e�n���ܹc{h��5��$�`^�*M�
����::a$�J³�̈́��-�Td4��
�#Q;{���<M�Z�~��+����a����_ٹk<: V�[x)�c��1��˥p ��5ǈ�;�ѳ�'_��7����� ,�ҡ�BS�(����47ך�(����������)ˊ�+Ra��X�(n,l�;M(���X���)&�n�є������=ܓ�%4���(�L��E����_�۝:逍�~�g6M�:SWQ�ݿ�w���{�����#����h���UBR9�哂�7ת'#$ _���XW>��.ލ��g<N�
�s	�A��#�"��)}p'x��7��4>�8�xIW[��O	�<E��?p��ސyn��A���I���1��i�7��9C�6Wt��OEK<4�f�W��,\���(��V�Z�����=,���\$GJ��W�/��%O�#]7곰�'�r�4d��S�qA(<�]�K]�m@l���D�pa�g�_����Z��m���O��'��=��-dF;�
(S��l���w2x��P�."/,f�>���@�-ņ|W.�+}�BU���e'r�o7���GGu��a.$��ik*[�`�B�36�򛦇��9��#�CьK�ai��W����ph�;w���p۱}W{.��^z9F��m�����5&��|�K�� C=>�	�;�Og"&�<`+X���8z9����,��(V���r�����L�:Z;k��������|;�옲�K	�a�l�X�Χs�S����0��pDk�לvR!#��Lo8��hDu��V<]�g^����I����K?[$�`��T᠁Q�s�B,��p'x+��:���͈��"���෢:3/�v��_�W�U.V���}g��]����߆����\S��6߿�K�~$���	���(?��=!��Q�Q*	2�p=K��)y�@}K��I�;�{�' ���� &t+��}��V���,C�oC7�I�g�^/�.��E[�I0Ĺ���`���:��н��QyT��=�{�����gp�jS�YA���)�w����h{��ޞ2�2΂���?%[�-!�:�n�����#Px���;��Y��}%@ގl@~�9
��Bmv`�w~���Յ�F?a1�+�(</��b��,�)�1�w	�	�֐�[�c7��T��{��iUZ�bU[�be�{������Q��r�H�+HNʬRdz��wa�T�q�@��B�����Ԙ�0�y8�!B�|+��{v<�[�_�Q��={��m;�C?2��RTB4�HS��	(���׼�Qz.���5��WX���?k�F��hR|��#/�cJiL���L��F`�0=�L۰�l�4*�+�u�V]tW'���=�;��9x�ӹ@x��<�M�D��R�q+o�3��0-N�>A5�O���;2t��̢:��'��HŴD��U�����&h��Kz�*�G�wŖ���FU݌�o���vO�E#�"(L�8x� ���`"<�I���g>�[���(O��{�6��
�z���a���~Uw��[e�9�_������F��|�m��t0雴�~����ѬpQǹ?x�|������pٮ��1y�p����Z񬺝�~�H���,�^�o^o�*�!���}<l�>�	*,WP� gL��U<%���Ȑ��������d��Ͷe�����0�����?��q�	؀�-��)E�����v"u�� -3d���h[��n(-�|�3�/	
&N�����eӬ�i���브\G����K�ZU�\�n�zG��gŠ���:)�bli���PV�{�i k�ৌ��X��j�4�Ppf�8GЙ�w�
�;���h�!B�D#zO�L��Lb��9
���sT���:���U%���y7F����J� �*.W��� pꝸ�Ʈ�i���oi�@
wڽy�`�+�:{&B��p�oe��)�]�0@��16\�)<}O�9eqکPa��積Y�:s��*,��M����O3q,Ohf޴���� ��(�tL3�/��r���(:5#��m���C���_10�Ą�3h,΅nQ8	�f=�w�ňF���:�뷆e��L	�Nx����o�vv����⿼D2����*7g<��ƿ�=�>�>!ܩ>�WyV�z���cia������0:�4�AQ&(�G��\?�ʰ ��o�f�ƌ^a�{ќ_�\y�����0��t���wa�^�������J����pB�ɿ����;C7�
'�&��������D^;��AA��d&ޭ�����¸u�t,�͛������(��&���b�o|����5�4ىI�"��c�Z�Ԫ���?���5O
���Eߎ4�^Ɲ^��w�����`V�\���Nf��Ѡ1��N�9+�}�𡃡𚢚=7�KS�}u��zC6��H�A��|A�+5�tI� B1o1�hu�%9(��É�;�~�Xn�U�-`���ˍĎLE��s��1:\�i��tƕ��k��|�V��:�:D9�f��v��6q�Qsb��t��X�P`"���G�݌���t���7k6�� a]8��՝�[x������D�]��*~�r`h�i�����N���x p0��/�B/��ɯ�����/9�6��]>7%�,P��(,#;vlo�/
e�����}��>�t6�%Q���=iG�k��,��5�D��P�K���į�盎�"gi�C	��/\�Yӧ'����߆��}���7S��ʭ�p� ��z�]C���T>��Tv���	�O��������^F�v��H��<��+N��s�w���k�u���0�=���k坳���1:����Z�=�#�8�����s��v#9��a�N��2�O��[��AD�DI'�)���������W��1=6u6Z��D�!�1�_Y�I%+-|�[��,��hc��ޔ��k{C~��B~�R��R���Rש�^e��������g���5�ۊ���g�>w�������y9-��\
���XG �7�g�p[�20\h8�93�L���J�*� �1��-J*(%���wk)\���|g,غ� �9s�6�sH� �M���և�	\$�FC{SyYt���s��X:��B��k@�QEsޫqU�:��h�+�wP�I�^�U��WZ����+(�����k���7���8��N�C���r��<��l=�ޙRX(55��O�qZ����F���8G��Q�8�Ps3��-�NF4��u�-� py[��²�9�hA4��"D��i@����MyQ�E#阖�p��KE*� /u �\�P�ov*T��?����a� nR��>��e��'�g:�u��s
�0�0,�:��!x�-��O9�����(G��"�xV�TY�c������pY�:��{��Ey�I�[��(pѳ��D�$�+,?O��/�>�����?�'9(3Ҟ�5yL���_������?k��;��K����*���8O��&��%�`�AV��ݔED�ַ�a���˒m�0�4����~m�fz?}g�:�s�����ϐI�$�ڰ���Kֻ-��?ܞy�����������F�o��X�%;��m1��CH�|�]~�e����F_0Վ�|V�	��@ӔQ��/$�������S`�����wv��y����l��VZ��J�w���n�[�:��e˖�ʺ���z@�JW�C��$~K#+!p�=�'���W���7���M�3�1�3y4�c�����g	k�/o`ј9W���n���ҙ+W��0hc������aapX�_��wL�����+Z����o���V�[[b?
�w����ɻ����#�l����&�ʝ�y�;e������P*re8�XZ}V�����5�VoK=!�~�c[��ҋ��c�u���MX��n�T#i�BqD
%�ԇņ@���2�s�=�px��]j��p���>�v��M�Dt)ڂ�;�����*���x�?��>�j�����+�����y-n�+ﴦ��R�Ϩr���݂85:�m�N�Un�]�ZW3�����lp��\N��N�^
���!_8������J�} ��$����ҭ�d �$ �Um�p���B�1@��������y���W�W�����3��>���	���X�M�а����yj��)�6��$ed��d�8�6W�F?G���Βq�F�6Ҵt��7}�<;����sl�p����h�;��Ny��:N^?���gB��7�=t��\GC�f��h�<F�$��f��^X8/JM1 P��i�3P�u�F�Q�Lzv�Pth��RB���y��\�m4o�6�G���%��,�3�����w��i��f���V���oo�x�;�=w��߳a�1�'M�٨�)V��D�Lqѡӌ��K�)d�i �6� �HVf�����?�� [�����4�Zc���S����tH0��h���g�����*~�8�>��3�[�m���Y'��̌Ɲ��[^Y��_���F�]��+��nun��yv���ߗ���=�no~�s��$LSR��H�w�޶/p1*Y�zU��ha4�h4(��4�\�=�w-�_��7��~��̽.�
���o{*�殁�s�E�e����vE>%+�rC���:�J���j�+W�5J��/� �=���"����']�$Q���h�tԓ�0����;�+[_	oK�)��+^���g�!Y�5�4�֭��W��?&�o��L�/S��4�u~ү�އ~g'��C��ڸ�x~���yXk��W�wơ����'>�/�&Sh�(3�/΀!M�h�ֿPrȑ����k_�җRV�9_[��������0Ee�e#��L�T��Pt�gEf��v"�(��(8��D*u�0���o?���۵D��nڸ)㱐�E��۽���\��~���e����_r��7-1�bQR��s�.�����g�?�p���u�|ɔ#���v�a���o�]�
�Q��Rl�ouU��m˖�m�N�e��Ԗܣ!�MU��:�c!8�/Bg��fm[�v]v��_w}{��}o�ȇ>��|������Q@�-�����`NB\�*0��Q�]�1�Q
���4�P��Fnُ�؏��U�scD+��&n�%�1�C�t�v�(&���ś���1W�X4������[?J[��i���.T��њ9��A�IZ�?}7�w��lw�yk���[�m��ﷷ[o�9:���C1|ӛ�i���v�=w����r�}o����]�~G�w�w����|[n�|������w��t_�����Eߏ<��a;y�����<��푇MK˖�����=��2(��8F�t���/��2efnm5x
L��b:�M����C[�C�q�?�XZ\A��tv���͸�E��5"K+T��P����|[{K�ٵ��T��1�v�>����P�A������} xh���)������}S��e��Is��9%��#=�ǩ�*{����)�\�����8�S�{��|=0N#�����x���Ii������^=�]���4��wr�xt\.��<�]���w�T����Fnx'�}����/
�{���nڡp���c�!#�T>ȥ�g[��y.�E�O�A� 7چ|�}�n���'9M�aay�G��?Ҟ��L*6֒:z�6�r�|榼~���7x�=��ږW�����7ܘ�x��+.�"���أ�F�/�6��-p�ޑ}mߡ}y��eW\ޮ���6kα���1��ɱ <�����ǉ�V,` |">�x�a��'`�~Π��3/�< C�D�
�DŇz8g=�W�;���+��N�4�Ve�T`A鶜sܕ�C��A۫�SQ���v�L'2�����6m���ŎF�̀,$�_�v��'1֖�_x�}�S�m�B;6M�dE��Tk��W��>�h$�
/+�v��8᳟�\Z,:C��,S@G�ٍ(5��\$�x�w�(A�>I���^�o�Ey�����Ĉ�-3�Y��0�YΖ-n��x��ٜ�p�ץe�`��.�4ܦ��u뭍Z�V�Y��N�Zv��T@�i�ՙqh��S���j��}軁��pQ ����{b����nO�I����7N׶��ٜ#*�fQP��|�}���9�T
�������� 8��7"�ì�:��>�b��Ȫs�曥%nѷ����ᷡ�S8|�'] 7'x��K����6?����������J�����"h
����O>�40:�
ydV������;�
�!��[�(?���Q�7�tc��إ�W�_��7�����]�w"����'�ǹK�!T�&��+h�x�!�Z�O�Z*�8�;���d9N���!L���t��`����a�E���N���z((����wq��8���	W�>�S��IAg5f���ɺ\tA�tLՐ;��ސ�W�F����?�{:��w�W�������䜼��5��~�?.�qm�vҽC�}�k9ā,φMs0g	 ˋ�B�Y0��|�?#��ky8�����k+�x�GPH��*#SR��_t��KO��_}����7�[b�y�%�H���h{�����O�Z�l*x_�����q_���7� eQ�������i۶�n�>+q<�ǴƐ���
9�uW��ե�V��ק^�Ϭ}�+8/J�8��r��JG�[@h�淾���J�G��*.��uLn��'��:w�Hˎ-�75@!��t��m�+R* ��a�
͗bS�wh�:[���i��Ď!L|��_�ug��^������a�g�:�Ky�)��A)�3~�_�9Y�ΚRV�U)>hdt��i����W#�8��{��Ҡ��]���Ԭi�:q�Ǔ�0��ra$~$�Ѡ�޽�ï/^��y
�yW���;ǀ[�OI�8=
�w�~�Q�\��@(�����7x=#�F
�s�=�q5^���u��fݱp���'�L��G8��>��̿k�Bo42"΂�O�����,
K*��XP&����s��m�Z�R4��l��$�:���a��L�&��R%iR�@*5#����_�����J��t�Ҝ���}���-	�$|GYM�/<�~���^	���r\�rU<�S�I�-��}B{W(������T�>������G�۰�j����2D���W�3�0�q�B9p���
�=���|�������2�������%ǋ_�*�Ug�+ݡ�i�ʣ�M~��o
���"r�c����9��� ����2�p�_���C�?�[o3'�9�gYs���qÑ#E#2�7a�?B��i�����h���wܞSݗnؘ
ޣ�>־e ��}�K���|�'41���#e�v�P��#�쵝;��w��۷�7(P�Y�=I�t��W�B�lْ����OF�
����G����i��rC�]�;�sW�Y_�>!�Đ�_�I�9�8��=����1�]�*�k(N��ɴ?_pޕ�MX�Y�AlZ(������¨��*�􈊿��[��(��Nw��ܙ&?V������Q�{C�ؑ�m߾��
v�
%��̘N�y`R���P6�'&�فG�ڵ4���od9�q�Ղ�)5QW����іMװ$��S��j�Oc��-S���1���	�b��5Tی�MY��h �F���0��s����� Ĕ���mw�����є��-L-]��BQ[��M���R6(ꐕPȔOcDJ�_�gaq�xO>ٕ(4��w<aI�:kuEy���$�A����I���X�M!�$i��֨F��yv���$�z�Eɨ	m�.�Wiچ�s�(jr�Zi�)��:�����z�<�!w8�	m�q�I)���>�Saڋ0F�h���Kk�#I/��^X�����l�V8k^;�:���H�q��TWo��YO,���p��׾?������[o�=+�.^�w�H��������ѱ`R���m1�f�\�8~�3�ʫܐ�~��#��0�π��Qm���V��\r����+�x�"��qy�����*7�xc��B���xDx�sZ#BƲ�k.k$�u�d�4���f�A�
�������ƶ�,W|����C'M�E�]����w	o���i�uI2��ڼv-}e%k������ՖqJT?��y7��)��/���%��:~­����؈�#����������ޞ�A�/<�^x��v8��싂f'�h�����jW]�2�c�X��_�F��oK�Gft�.fժ�����gw@�Y�>�sWV�녂����hV�RB��A���z�ogg���A�tq��m۲�y������}��P^L��3*e�+��1�)
���Q�w���&~3�%H	b�� v��ER� �-�y��[��v�a1��� �����:{ڇ�;�	� ��.�P�V�,۲,[���ef�2�d%��e%�d���{��{��>�l�E~�z�H���FT�w�������� ��|Y�?�����S����Ӳa58槈ԩ�&���w7���ƟL�h����VF�0J��*� b�;e/��k���qTΡ�8T�]{]
ď)0К�k�����|�g�^��%K��˓]�_�das�w=/����*4q���:�ڰac{��'���%�w�~!z ���n�����I�#���fD����ַ���^�,�28n�I�'~3`n��|�ː��bq�½���xTWt������B���F(����{F�w�K��}.�p�`�78�&��A�2����%)��F�!�በ|6���������k�v����z5j�7�ϹZ�#�x!c�B��/	U�����{���)=�W����iS�圃�y|g���1��7p_t:��\���0$><��R������{�@�^Oq��=Ca��p�v�~A�׋�H�г,�̫҆O�P�욽�h_�v+h�Q��}2��}g��8�A�Ϝ߅�k�md�{�0�G�X�nmv�Ѓy)�O8S�� d���Sv�&��d�dD"����&�#��P�$��;A^�����z>&x"����wr=s�ߜ%o�J_�dՐ�8)�����o��s�>��2FG�`�9���qs�x������<'N���M	8���w(�l��0��l#��%zT'cc��B�7ϵ7smT;���nͪ�`��v����C��>���Bo��i2	NG�i3gLK��6 3C̚=/���6�&�
�#��š�t��& P�\�[�n�9#���J������қщ_c��n<sej�?�8f�� 0̀ȳ7�X�,���2���C��7#ܘ.�86mٔB���)z������=��C�đ�m�;#��F�a�HC}ʐa,#����#�E��}�0��=F�D������ʹ��#7�@������d��1�Q9�"_\eD�>8���KC~��P�@�K����������ߞ۟f�����C���h���[�����FPz�*�LeX�P|�<<z�@Y��{�)�����m��?���d�y'=mQ���r�*��*M�
�\��4����`�#��{�Q���P�6�z��ǒ>MH�c��	���_��_|�6�XP����{���������a�Y}��M$g�8���սw�:
��P�q(� �4��Wh�9������Ig�Fe���)����{��p.^5�y�Q���jϞ��Q�ݠ��0���#q�(z���]בe���Pp�zU���A�������!�t2�?�C��9�s��5䡃�����q�P��@qv��S=}4�[O�Je����0lѼI�&�3�o��UW���'�p�������5p���NG=Gʀ�A\T ��1��Y�p��f�e(���3��x�gd{?�>q$�h�E���?������`��!��K�F��u�����B�����ό(`�����6ٝ�R�7ȀBS�G��s��h�c@vF}9q�T��0j�L�>���D'��v�̩����m����y7~R1I�衣��9u�h�|�e�=�yG�;oV[�rMtV�:1|�����	�ԨWnB�q�Z�a�tj�8���AX.�m����>�i�gd��N�
�	F�H�*�����1���qO��̩a5b���(	c1:�����k���>�6u���|��$L�|�+_kGkS'���ƌf&jLn_/b���^�����Wn���� ~��s.��	���;ߑ�f�Bʊ�z�G!�19@��CYJ���!����u���|*'�*
&4\e°�T����g�j���KW=�L���O��@p�����O�3��a{�0�Ł��m$GB������ey�^�4���
n��%�-�� U��'|3v~�W�eN�&�"��#x"P�i���7é＝�3�;rr�wz�x��1�[C���6lx6�}/M�
}~C_��+SQ��X�o��c���������u�Ѫ#@.���b�}P
iԠo�VV;��F�K߮��W�E����kËſ�d_�?X>����T<�Vܒ'b
�LO:�eY|�Ɉ��۲�������N��������]���K{U���i3sؾ�J^�����?R��*���a/.��xg�O�ԤZ���w�T=�ԇc������C��Wz���T�\=�銏��f�	��4� e�ǌ��1<�t��0#+�|�͏�����厷���Ї��ky�QΕ9�%���a|_�PC�t#�u����(ߙ��y��BpP���*���e�y��8:�"�v�x�6yl��G�]�U��=����;���m��C��۸�?�;<~�L����m�aԼ�-Z������vŪ�ۼ�6��x~���5���Y�+�D���W�ܞ��N6�,��.�{Og�[�s;��-f�`vWJ_�2-�4B�7Í��. �C'��ګV]��M��?�Z��\�&N��6n��~�w�=t�C�ؑ�axM�Be�_G�Qs՚5�ɞ�'O�2!.�W���
��T���7#�L��<����zf���0�xo���f.0�9�K,`ĭI\3�e����ݧ�;c>S��F��#o�0��1�Np(n/�J�Ћ��ܝ��s�@�z"}O���@e��؍��0>F���� $��a0� �s�w�02����{eP/@�,!���g���v(%�f�zg������+{�&��!�=G�W^0�2�m�E������ҟ;��=���wߕ��X��O���0�ixɐ$��R�F�Y'S^����O��{��˓���I��X#Z5��K����$�txK�����=����Tĥ�G�����B��}9��Ү4�ų�+m�w?�~0~ŭ�A(�
hm����O�T�;\�P�<�'#����:u�ʷ<nV�ƃ6:�Q�9�JIY�؂��?�����o�׾��jk���Ac?�я�;�qg[:@�9O�ߙ�O|.�7��Z/�Y�A���(g��,7�ї<�J}#��~�g�н.�2��+d^#�°�?���x�������4,X���&����:�:���j�����ۖ綥g�7~�72i+>RfЋ��c�P�e<pP��uaF����C��_�����4��F�m�&����ƄN���)C��쏷+V/o'No/���~��0��x��=5�^�gOm��mo{ۛ�ꫮh+W�	�fMȓ��!�W.�DaĢa��40k��u�Po����r�Ϝ1+WO8�kW�5�v8���ڍY���ǎ��9;���O����UQ�FLe��Qoڴ��{߽mɲ�m��%�,��s~���A3���� ��z��� q�]��wA/�yp�}ũ��x#a0͋A�+d9�Y@����Wo��0��h�~��y(���6ݼ%z*�(��ɸz�ڄ  �x�"�į�U����0�M�xu��[*�7'�uy�(C�k�a��������=�LO��܍�bV~��+p�0�O\��+��i���œo	�N���x�1�Fá9Mf��7����G�[(ڕ���B�p�o�o�e�ko%a�b��&e^���I{��m���A�c��MZ�Ť 'z��1�X÷VnԼ(���=WK�}�o�9%�8��1�*���J�ǩ��j3���pA~33�c[38���k�k7�pc�`xk�0�&�O��\���%~�I[qj�v��h{m�Z��f踮����q[���+��К�̅�����Ӯ�]f�|44o�}&�e9�8��i��|~g���kR�/-��u�x�w���]�h�	���b���0�ƴl�mϋa�M頷'�x�=�ԓ9�u������CFH�<-�J�������='�H9����Խ�B�x�4��Gs�S�l��|�_~�� ��<]�A�h�W[#�ݘ1
m�P��l��4�i�X�X'��d�v��h	>�_y-��xht�C��|�B)YB�)��D�:/7��g��䶹���Yt!��� ����C^�g��M�mn���oO=��;��s0fǡ?�_��7e����%��ǜ��۬�sCFM��^5��F�������&
k\g��E�����ԩ��z�;{nX������+r�@ج<��A3q¤00���}n��7ܠz�W���A�B�C �xo����Ź��]���#=x�C�;�����rvtO�!2A���RZu��o��
.��b�rq��8�q���j�r��e�yPLO=�ty�Z��7>LE�PH��{_�/�ȳ���q�����+=F%����q�M�ϐ��WvsG[��{�
���G���e���n�,��A��B�J��w0t)��iT[
��#��|��9�?�~�:=A�Ug�}�s��xh=�3f��eӋ�,�v�1���/[H�u��>�a������\��]�,���;v�>ݓy�z׳D�� ���#(�:���-ZՕS���$�˰����07R]f�;4���F�xf�*�k"��(�����}P��ͅ�G���H:��˃�`�7:DFJѐ����/��P=y�Gsx/+	k�����L{��+�m��)cЕ⦄�z��W����O�8�uPT߾��IK?�`�ߎ��,T&���K���yL���+��}�,@�j�U9fݺk�P��T�i�C�~F;vl���mX�1�M����Gi���=��<�W�ds���$w�yf}�U��aD�������U��SA��C��ɟ��<چ���hR~&���y۝okx��.k�N�U �Р6������{�0*vʢ���d�t��zB>��VK^�7��r~'#�<I�:�*EP:�:���}z�Κ�<6��(�U��J�G_��qҽ��i�MoЭ�ޔ+����y���mϾCa�H3�NYr<;��8�fL�x[ަN��f���'O�v���~)�5
?H,�3���B�"�X���f�`��ر�gJ
ZgZ�<�D�ɝ�Cx�`.��!��ryh�8�E �bʳC=����Hv>�+^��6�_�*qT۷w_�/z/���TZzI�V�QO�̈�������%xF�ȸ//�X��`����z1�%C��i`�gB�j+u��/�13g�X���	����
?u-�q�=d�~�P���s�n�Ӧ�����
�W(e/}�pS�u/���+���b�r�*oW�	��<�F�F7=����]���F�D4{g�mc��]A��ڦ�9���>�Co��.KCB:����m��ω���.�1�'�Xf�v���7={qV��oS��2V�έȳ����<tz��M���T�x�����[�����z�Ǐ�}���aP�?x���`5�^�6%��F ������Cx�!R���Y�L9$D��VT���х@Z��K��j㗂s���S�g�`���o����˶v���7�>=*.�q�[	�pp�rH��2�_CsVJ�w��A ��g��l���O�y��e������o?�T�5Ϝ�2���Mִ�v����˂�)a��\����ӨU����@��v{]�Ϸ�FՍa���B��G�E���,e� ���D4�=�F�`O����9������lƌ����o}+�֐?}u��h?�����w�AnE�I��a}�bӼ�QNGgA^��zK[��6~܄�ۄ/��vS~P:�x�6"��n�t�FL�a�4����g+ �ѱ�ȴ@Q��ҙ�G�;��t��i�X��P������Dt@y���u�Є�t��[_-�f��\2#d��١�����K���m�[U�4.���H0ƹ����%�o~���\���V��^�K�����GB@�ñ(z�˖��I���3uW �N�ryf�B���tN�8�&O�����
��#ʻ�g`����](�3���)x
@�Է�����p�]5~ũ��K�Cȕ1���6�,����3�ZƊގe��c�\WmCb~.�2j09AR¶�?j�� ��I����2F/gz�z�\�}� �n��*�4��+�M
;z>/�?�ƅB}s1|?��rp��(��w����ӃG�zd�czjF��u:�e��Eaq"ܷo{��ޖJ�@%$)?|u���g."8�@*�={(���w���^�}}�o�'�� W��E?���Mc��	���S���QWC[G"?�M�N����8�G�e�~Z�8~(y�Ҁ���S�:�<��
���q�u�s����|�.���?��v���FLm�=�5�/�v�/U�#|͈6�����}�CJe����\�di M@���rxo^~��4*ң���®ğ�j(
^�~2��M����ڝA��m����aXَ��5�ؚɓ��+V�J�l�q^���Ç'�B�e���iT>z��'�^�	����g����#�x�x{��ڳ�2p���*vkG�}(�����>�[y��^��-��ƒ�*��4��ţ�Fܟ���[o�-~�
����p5/�L3uN��\��7�b��Gc���1c�T��$<[���N��!�&?�$*���a3��_<�y53f���r�)5����g�g��`ْVÐO����#Z6h(e�0�s���9�W�Cر��|;.����hI��4��j�\��]���l޼#�iS�P�N�P��=����F�N�a���[{U��Y�焎p����CY^-��F�3j �@<"F$z^��
([��'�8+k�����ʴV�ҵ���{��=G��^�����p�H�V�4L�}�g<=����gNYas">9�V��:o�1A��������޺3=@c�AG6�n�^
��o�YoפZP��^W�BA�l|ʢ��I"��y]�3��繟B<�<��9� +O�{ �6�|�7=48"\02O�`]F��B�X�Ux�3x�8����`}�ION�[a0_�Q�B�L�@����S�+�KAů ���3t]|!?sZ�o�{��.�'���\��ڸ�~|��	u����C!����_wC�jH��m�( GG���۱텶c�m�.�ъ�mﾽmw(�=���C�{��?�8}ƴ4
=!G��y[�*p$�(u���A�l����w�!��ĥZ4�(_��9����FG=m30&{��$Qg�)�o�I�q��G4jY�e�&�l	���pC�s�=Q94i��䜷�a��I[ǿH�7/�]|.�(}(�x¾�vYf�9�xx�D�^�	|0H��~��:;dz����̾ߕ�tz�㆜��{<��N��:n\)e�������!�b���F�3�ÓƓ��pȰiIK��b���HG��es��Փ��+�0y��g���	�gs�i�>C�]<`��CI?�����{�'����ڎq更�{�k_��k؄!�~���`�����n�������#ml"G;���n�vܰ~C���ږ�[ڄ0t�9:Pw�p�ͅ3��C[��������ӧ�LJ/��I�xt���}���_�eN�7����<�y��D;M
C�h�[��w��ͻb����Uۖ�Ar4y<h�<��7�{��.��:�K����x6\g�h�h�[G������0��#��tB"�{*�gU[0z�ݩ�c�#?my(��a�1mR�z�<�͛C'G;�]�&�3�͞3?ht^�x�^M���0%rR)k��2�
W�{c����}C�p��"�(��z�J�m͈`�p��/@���AP����U���=���!��YDo���w����0�BI��F^ʪ��'�<�E(�{�q�}�T�Q�	�����ɞ���H�x�xWtaݍ��|6�ِ7�l
��^(q*]e�:]*��~��ڧ��;��uU��O�+x޿6-CH��;'��n}Wʨ��^�@|��/�wC�*_�7�E��b8�U��o��g��7��A��fϞ2��|�BsL<�����V��o�5zEk�ګִ��vs{�;�l�����@�I��a$��5w��vY(�̗�2X�xQ[|�b�em�K�UkV��+���K����t˭�L웞������\=��q3�"&�}Ҷ
�F4����W�#9?ʳ0�d~��I�����m�������� @�B8ħ�ڤ�#L�<>¤(���wro���Z��;oE����xw���k���'�ۦ϶g�}*��h��!;��%��"�33oN�4�̍v��-��-\��a��x���Dw;p�
Ï��.m+��z�Њ+�����>�K:#�w~��ʽ�~����ɟ�i��g�!��xq���~�BIyN�H�Ac^�����7�hJ'�p�w��U��輐�:3�HuZ�����6��#���z�8=$a��/;�ix�n�k�4��W��_�R*x���0�mzf)�a�1aY]�\-}��[Ƃ��������)��)V�N�2�C�!s� �� �L���]��C��e`�S����/��=���s�S�k59��y >�Lw���^j��<6��@�§ou��K�&��o�!�� Ϸx<��8�Q�ˡ���+��2��T�H�W,�Q�R=�1�G��妠���Բ�b�ctl���4�x�x��%#�����~5���>àRB �A����T@0`�R@�s�\#�z��]Az��x�JЖ��]	�=���be�#�|� Ho���,���?�I�+� B�܉�L���9W�2��)���c�� �r�"4��	�Z:���:�;a�Vً�<2}�⌄.�*����*<^�
�����U�I�W!�>\n�0F3�o�ԻJ3��7�u8q�Y�=	ˮh�Q���<����[:��ʕ�Bپ%��喛�u�]ۮ���+���k�˂T��\su[~��v�e�-\xY[�n�����������ol+�/c&wT�
!���s�W=l!�U�V��V_ٮY+�j7\����k��^sS��֛�m7��ׄ!�W'���F\��ԥ�LN���]4�{q{�����.��'>���#�&�㝓A������6~\(��L&��&����m��0d&�ub��S'ǻ�9<e��c�����w���τ��4�0��Um�U��q���&��g�N���M����Y�n���vy����u�]�gk���'»�;���v�o�U1�)n��5i<�}xey��Ew.E����v�c�7��$�������~����S�<uN��p[($�`8���㎜��Z×d
υ����� �����Q�![�1��3��|<����2�t���ރ��dT	����o�ms�5�g���.w�Y���'�1xy���Vy�u�桷8A�LY`�����j�wv�5�ޤ`��Q�(�se0�V���2*�м�\��0��	-}ƻ�ă+)�%���3x��݌�2-zF�x}k���c��ںڻ��߿T�ŭ������E�B�r�g&�u�dv̧M���T)�2�O�nۺ5'��z����l�R}i�_m����R%��Ȯ��(1����a5��t ���k�{�+�8֯OFEԾ�`�L=���Qa�l� 6�������g���.Y�n��_1��KǕB�(zH�r�Ӄy0��,������y(�qs�=)=�!�=yk�[ �"�
�z_ߤ������ .�$��V�J�Wz<]���`�����x��`(8�^Oo��g��ڹ���{�;A���8�U��������?;z���ŋ ?�������j���r����s5�k_w{{�kCi�xC�������7�����	��6z�����R�/]���
gvʳ��~O�&�u(��Ӧ��q�>)��ӢG83���Acs���s���3�-_:��Y��]�bi[�fu�by(�d�P�J� vo��y�f��\CI��� ���A���<C�̪���>�X*���yPu��'��@G��b��7'��	���09�ᑚV�p�ء�����[���1��ctpO;s�H�c��3&�[n��]ݺvݵW�׼����;�er]���0o���vۭ7�;�����ቺ<$x�ڜС���pH�G>�c9W�� W��B��%7 ���W�w�CS)U���Hj��gd���}�AI��
��pӛ���-<aX����d��?����O~2e������'��a��:�=0l �&��aO/� �i�6�JՓ�׊'���>�P�<@�!N�?0��,��8����:�9oIy��T�yGa��y��Ǵ�3R�X�����{��>י9F������s�����9ў�e|�;0�<ȯ��w%L���ɽa��0th5&c�^�w��8W� �\~�_��t�;bx����-�\x��-.0tŰ�e�<C.h�J�0�p��6\2���^�q=Ӹ�Xb	"7���\���3�<�d�@y9đ6���IYE�U�"�<W�z�,�u4BZ�ȍ��g���`��`����g���8��	�<�$��#?����w�;{��~׻�?����?����s�O��5���7��{C��D|��Z~E����P<2���܃�^	d�țA�ΑC^����y_,_����x�mH�T;ϵǹ8#����;�lsn.�g��10{o��32���4����W^1����ߏ����sU��0h��̕��Lo�w�!h��;�������5��ۂV�HC疛oj7�rc[���\)hbo�����z�B�6i(:A§�m��i��i��k��ʡ����DO��DǸ��!q$ze�QEC��SV�o+��!a6�}�8#b���6{�܎�P�hX<�9l&�N�w��<��AB�H�m?ƌfd�s���㸎6G��£��W}��D�����ϡ�&F�ҍ�>���߷��ݽ#������aЬm�^�6������`�W�Ya�r��w��׭K#�P��g���Xȟ�q?<$=R{s0L�������Y�;��淫��D�]ʒT�a�-��Kɛ�oζ늦�GiH�m���7���ʯ�J�jRn ���iي�����4�CT"r��˗,�4�W�B�#�����8�lN^�ݽ!6E�;:K�a�?�)��%-2̐�O��G�{�����G6<u�ُ�؏e�mႅ�ߍ��ô���s�ˡ��3g:3�`yt�a��PgD
�Y��.^�FuA�Zz�����{$�܋%�1�B�k#����
|���:�^�^x~e�����o��2j�l�Px:x��Q��0T��z!�M���߃�X��j�;��cpE@�����ѓ��[�����t�c����4�y������\�u�(��o�K��H���\�b��X���c�_��mf<�W:��cP�A�]_�py���$�a�'����̙5;�m5c���W�8�D�[��[=̢�����_��<��������7�M�����.�����ڿ���������������o���W5�z�K��K�����S��|(��x������#�����3��Y��`��^�ީ�ȴ�L@�Jo�� �ᶗe���,W���S�D�۹T�3-�6�r]�^`�^]A�n��]�蓰2�q�M7f>#�wf�ګr�#�fU�e�a�E�-�9(!GC��I���C�Su�ct'O��>��㇃x(�396<<c���q(ڕB:ю	!���S��#u�+��u���>+oJ3*���-ޔV�h�y��~J��39F���R,�7�~l*���6*��!��gApy�M��5�駌�;�f�8�ErD��4�����&B�|I��b�<'�Q`����&O�qEzm�]�.X�x�&�̜�M<}�>�rl+�Lȵ2���hd���x
�l4��� ���>sY��F�hx���w�����t�A�{8��N�I�:[�Oi����u�^���-����o��<
�F��u�O�D��c�����燇'��rkz�xZtڔ��I^Q�'�K�^rk��a �8�uό:m�� ���F��Q�1ax��@���\J�({�����w�����&)[�<9�+�,eS4����n��m�EǑ��D~҆3���/��ô:�X�~�}��pϫܝ��
��\�4�׵ʇ71)>��0&��c1�-��qg{wj:oL�</�gn' 9�R��Յ�a� �'Bո�c�zHh��+��V��:��b�2qdG�j�"��F��T��%>�(��1�兾��$=]xk����*�I7W�:�қ L<C���zﹱbe�N\�tB�	�~������C�w���B�)�G�I�.���!HWe��M�����Uߟ�s@��}P�����p���Ls���]�t�[��~�����E^y����F>���|		�<rJ�0T`\��5�s�MB��`s9�s�W�9{Fҳ�6쒎�����ۄ`Ҥ��6>z��ņy���
�lu�C^)K�O� �Oa�v�<��F�����P�\Ɇ[��M�g�x�{�j��sJ �S���AO����u��+��x8a�PM9Æ!B���o�Y�>��7�{�Zq-�i1`�؎?�߮,�3��"f�wOd�*q?y�6�ʲ�q�S�<*�f�/dС��]�'E��qr��8����ɫkV_��.Z|Y�)���Υ�ښRӛ������% ��
�+�)��ƀ4O�j�\�u�ҹ)�l�Ը��{&i�k�j��maH��/�B��������w��I[�l���{�h+�z�N��`������^�1)����D��l9��s82��&���+=�PN���iQ6�q��I#��1d�%����S4o�8r��d�q�o�� ��� ��0��~;������ڻ���\5f� ��WY�<��` ރsx�ǐ_��#_�읢>�3�:x�0����)2�P�x[��l�w-�W>y���F�g�вP�
�ґf�G/��ŇQ��yN�:N���C����&�8^DzQ�,�����@���T�ʨ�0����DH ��������x� 4T�'b{C�z~.�hĄ�F����ܦ�m����z��b�<�<}���Czꦞҕ����s1L�"���d�=�X���ʯ2��P$z0)���W5��72�.��?+7�/�p�5�{����ەV�-`r+sz�	iJ��^�Ty
*�
����g~�W���_�C=w����I�gA�>�{l	&¹��T��gd:*`�+��;�C���u��S9	���氭A�R�]������{�����\�J^���Z�tY�0yj.?�5��O����	q�|������!w���l�c��:~�����<'(�ь�>�ϸ!x�<Ս�&��ǽe��I���%��ΕQU�4W�`�4ib���xU�a:q
\ŗ����%�g���wH�^���"-'�ظ��)S���45~��ҦͰ!�x?&���6g��6c漈7=�$��\n���q����ڜ���r��>�=~�m۾5��}~l�o/��l'q���4D��bP4"�#�q�|��T��>&��p��2��l�n��q:@)�����R.
�;)2|���w�7�guD�V���4��Z]�����g�V]z~]Y�C��/�I��x���$}�!�Wơ}�	��1�6~��9�2J^�g�	C�/��=O�֤0D�h��>�N��1�1����[䮡�:_�\�}���o������s?����~�G�� �)`�:tdXF���(/��d�"-e�]R~8�Wѹ|y�� ͙V��=_x��4���G�O�f���~�C['�Fū}
�!�m��l������R��g�P���n�O|�)��k!S��iu�^]xU����xW����A8t�t�4�Z+�aS�F\�/׬�PB5n�Y��ϡ�7*��s�K�8�J4.�C�e��<I!���<����b{�w��Ɋ�O|��/��/�ީ������D>ƌ�8���s�EyqP�����aàRA�.(\��+]�u�k�[�@	�����}�z/H��T��wECgd<0x?�y���#�	����Go}J����@O�m��+u޻ww붳��&=�أm��!�g[ڄ�9c_��ڗ�����#��
�(U���{޸qӰ0��`{>�����B�Do0��]a�lܼ�m�v������x�#!l�E;w�k�ϽTFE�S�ì�_�ډS�ہC���۞H[��w����E9�iJ=1��c�U΃H	�З}��a������,��qp&�v ��h���!Lq�}����rz��������������z���C�C9X�n⽭�'G�1�(Gb{��h����䎶w��v�#���#v-߿w_.8�[�m[�[�-mF����n��ծ�۷o���{_h��_{(:+�9��"(����
w����$?���h?��?��R�Cd��G>��X .�(���A��J/��0? 4뛤�H_s��v�*#Y<����g�ͨ�=���Y��eAgU'
�]�S���H�A[
�Y}C�'���{z�7xq���W��p&P�e`S�i�L����i(/,�(s�oS��_�3��kK�yl�hB��׬γ����76�;����Ʒ}��φ�"��^TG�R9��+�2Ev�'��=�>@:��+���g5�Pu/å��Iýӳm4���/m��j�F�����OP�3�B�$Σٽ�:�ڼ���e�9���99�P/tP�V�
�,�7����*l��	\勁k�w�<W�m�k�E����b�j �V�
��F�� ����[�{ġ��9~¸\���>����{�=�Գ��"&3��l��*�O0��P����'����ﶿ���K�b_�pon���1F�ׁo1���ʌ�g�y6�X]*_���B�U.����,�q�.ܶ�n� a��cdl]����ۑ 4T���B]��;�ܓW���E_y	�ڰ��8զ�Y��[��M��*���J�u�o+�����U����_��ʨ���w��
�������۶?����0+Rx,	>:4�d��,ǦM��x��.ȹ��ol[�lm[C��]O=ݞݰ�m��5�!`�q9|t0z�C�=�~C��)�{���և�(���7��O�xۓ�����g�on�"�Ç�|7
�P�gg��-����7ڭ6�+!��~��C?��w��^8���	nn�tl�nb�S�SQ:O��d�0jZ7���d��9<BnTi�@�:#����qæ42�yvc�;v80uo��ܶ�;�ø+ȃAcӷ�w�ǃ����� �Ǧ�x��uh#�0��n=�PvF�Æ!ۡ�_\�/��tfb��T�YJM.�����ؽ�<� ���{O�t���������i7:���k�EC.�qT�}m���X���bE���"�Q�l��<������_����4L��&Y� v g (��L ����gP��ȟ�p����?��;SI[Y��P�򢓯E~�3�oʺ�?��#mߞ}Y�|�<h��w� *���p�������������������-#ɱ��[�g������7G�x�Z��cN�v�>z��d�ؓMy�g�WΜ|2}z��jGFH�I9�=I^<�p��Н �+�+��xtOw��s��r˺����!�sc�s[�cfZvl��Bt�rϢ�9+/�ͅ�[0�yr��b�v��j��r����x�Nci@B��`R�! ��b�j ���LN�^��
�5l]�WdydCz?u/~~GBX*z�m��&g&�>�ģ�=u��jd�W���w=��(���䭾ʫ���Xa̩+.����(A���9��6��/���zx^q+N���	����7�h�]�%���R/U-�4ab�0T~�s!$y0���5���B�˟p&�����q�ǐ=,ϕ��<�[��5�C������WF�H\��� mU�q��beq��9��w��\*e��WnsR|a㾽��ے��Z
�N�΄�5�״uk����W���0���z�`���{�=߹'�wr��=
��4f�D���ٓ;���]>Ǎ���Z��!�9�$,[�۠�0�|6)<i�-y���5:��*��4=/��r��C?�Q�gu��0e��ЂM�}A����Ҧ��c�hMO���Љ'K�'\�a���'�A4X��Ĩ��M�������
F�� q��?����#��q��޶w���۲=p��Y�y��P(O�a�q�����4��������GJ�>>ӦN�t)p��r_1V��w��s��%j/Z����j�7<�F�۸Ӱ����n��?����}#��a�nh��뿞`�):L��N��_��u*��J�w���l��Dj;��3�9����ĳ��I;[�mȬNY�{���e�I��WoF����[�&�_uպ����{�0��*L���ّ���7�����������\�â>ʬ�����My2��ʠ3��=S_��=9E�A���#�߼,����/�i����}���s�!Opn�����<����-�L>�=e�΀�h�ud=Ÿ�Rve�w�w�g20y�;����|�Gc���P�xs̨�m���WC�D���E9a�ķ�a��́sF_�=�8~����3ڢŋ��y�a^FM��W����% Iի�|����`�#�_��_KB_cjX��4��A�l�>6ߋ����w�`���`�$�h,�%<��T�M�tȟ��;vno���~����o�q޿���l�'{:�L�|I���D�4&
�K13خ������<�D�{�����=f7��!�^�0H��}7X�z��C<����3N���]	�U�ݗ��ַ�BWN�d<Xq�\�q��C������!X�~��9^g
!h�7Qu��9���U�|�-m������Ӎ�t�t0��(+74�+C�ھ�{��L	ږ`�9",V�}���G\c�9�������0px��]=���-������/"��Ƥ5�fWnq=��gӥN۩�a7cڌt��kseԕb2g�+WY,�$p��(N=�>����̻������������K0��^�pAӳ�̓c�-w��h�M�'����aT���F��1'__�0짲=zn�����q������4&ʦ���b4���CA�ӦLj3�2�Xm�ߖ�fZ��__n������84�%��݌�}a@MM�m��E�x�|��P�&��P�D|����l����h��N��8��!u�[=�?'zG��v����y7ڽdRd��7����xc����j��E���>���}r5���tB��V������rc>|k�ȪI{�������Cn�O�k�記$l�	��Cl��"��Э�'��l3��|��є�ro�o�'�g���B�-�8Z������j�_�tv
�}ݵצ7�0/ck��-m钥y�C�F։��7�1��P֍!��19�X�ݳ49�7���?;h�D��}����~"���o�f���L�&�}A�V_�! m��{ۼ.�����|1^��.��;>�K��B/�yC���'i(���|�[ߒ�׻��N�i�#q���]NE(=hފ!��YL�g�E����cN�Z�vd	��JG��q���sKNe����^D�cFm��[�ׯm�,l'�m߹��0�oS��L����&��u�?jk���u���]��v����(�>�e��2�W^�-�[� 1Q>��[��������M��C!�ʭ�ff�r�y�J4�!4��;��ӻL0�C�V��W<�N���S��`���a,Z�$��ԓO��|8ܲZ���Ͽa��c���='?F��1�8����4'�ʵ*����*pN
�mm�=�*����ΐ���?��O�FS?E6<6��ҥKڵ�^�;�RnW^�*Ǎm�����~�UkڪU���˖do�>�v?ߞ#�
6<o 7��v�|[{g(�+W_і-[�n��+�g��6S��`�OX}�vu�ܔ�G�Fh�]�/���]�w�7����Ӹ����I���E�5��������d�~��J�����Ľ��OJmi����ٽ'.�耿'�x*��S)�jr�HyԤ=�SGx��&��� �۪�2���0~������)ϙ2vn��^���;v�%��Lo��0h����.�<<O��(�M�e�w�?�U�bz;QΤ!l��e���l�o���<Ҷ�	����#d�'�>SAW2C�2^KM��L������'+f������F��e	vN������"]����F�v��ڟǳh3�Ij7ʋ�j�S�"�ᴋ^.�#�(��<�:VR���`|��_y�`�����	@��3�'�W�:ڜ"�����>|/_�,="d��Iڍ2ȓ�A[�r���)e�k{����˰y����P�<Ah��(�s6�3�L�w���]�A�M|��g�ݻ�D�����M![,�GCd��('
��^��i�*3O�=߹7���k���y�]8���*�m����|�b��W��x���@N��'���%x8$��1��7�+]�=�?�p��׿!���ħ4�	y���e���&�-�����ŋ.K���%C���2,t3���>�ς��\���t*x�l����C��
ޚҞ�ߴy{{��h��a	\�w6�̋o�͜15w�fp�s��-�Q���%3j��!QjD1�)j8˞��4hM��h՘ �bj'��� u�(w���#D5\7^�O������C���46��1���G~�GR�#�����O�X0E��b�4��ĭW����=����Ͱ��]���@Q��R���D|�7�"�L��sP���]����7_W�(w7�3�3���C�y���:N	q=7t�}y{7xn�+>fβ�uz2���������]�.�-����֋��)��|�����@���S�������HVNq�A(�yV��֞�Q��ܽ	��T[����h���B<�ۧ�Y�VJ���<�����py���VsS�ȫ&��+oe1E/�\,����9�el�.��ؙ��Hk�����!,���tDȬh��#�n� "ROiH����e�Q���(D�� Q��G��a�G�4mN��x�Q��tt8*��yL�K%i��+�����p)��q�c����0zx�(Z��c-������l�BxK�9��'���Щ��FP?�Yu�x=Z�E�L�@��x��ܜ�ft"(���i��򆷉W/�W�:���0�`΍E�3/2/�\���n���%x�p%�hi��`R����錑�e�[��&���vd�<��Cm��m)��3�?B�K^L&?<�bh2d(�Ō��3�-�{i�X�<�K6������wO�+�@�[�Dy���]w%�t��iԠ�����4�������l���ѹ�Ud���ԑǓ�"�.�됒�����/�.n�9��F�0CT��c�Y���o���I�\�I����}m��V�ywڑ�Z�hq�\��/��r�|�r�s�2��Ȇ�I�3����tUν۸��ȣτ|�=l<�n�C��	�-��`�i��"���坕�O3�.^MxU<5��X���FE@�1���o�j���$�1�w����C��=<��u�5ʊ_���S'��L����u�����xӍ) �-]�>u��J�cDLNW��~e�z���L�5�������`~�P]\����Ȱ������I��Ȱ)��F~�^����A	QF��#w��1���	�'�x<z�O�2V=�R�޻�O�gb�3��{W��]�fm���u)�ٯ��>�b��=�œO>��Bzi<0��D\C�a��V�ţ���B��4��6�Ф�'����
�he��0��5
Cچ�Тg��1sF҇a#B������u�$���I�N���F��{tٯ'��U��\�F��dwI�;u5q���m��9>3�Ī����y�ࡶ#�Ɇ���0rt�G/yj��xq�.�.��M��z4D�=y�F��gq Gꡬ�kK�jGn�8�7��4�YO�
�d(��⬡����ǣHӕA�(�U��@&O�2-�at�Nա���m0�O<Ux�����
껂zW���i��z'�E��y�u���/�g �аyU�^�:c:d�y�/�&�6����k�ub�my����p�?`��4��<�JZ�2�����cE�I�?�x�(���k�����~JW����~Vz�׉�~xx�tJ|� �V��H^<� �NNF'�o
��k�e\m���<�m��?/etn۶�=��IW�D�-['[>��ϧq[���6�Q�w���|���ݍ��y���,�<�+G�2�p[�a<�|�p�n���ؽJ]&��5�ڔɩ�_�䪺�jk4	��}^CWA�<��}>c��o�;�;��G~�G�^2�Y������C������9\]�������.��9?�h����jE�<�B�:�!~��dީ6#d���h>m��(Ǽ��3"���Y
Y#a$��S09�J��f�@\i(��D�X�1I��d4JCcbD¨ ��`yr��x~ϵ��J8�O^�]ɵ�^�^
ϸK1�c�=�=�����C�����H����p�e9�c�Q�๭)e�G����������Grc'2y5���u�7C!�.ɬ�xU�z.0ؔ	������ʥ�)C�|'���nܡ��7iS������]Mz�+C6��Ĭ��0TH����ڴqs�ع����t�3�FCQ�C����>��<箻����x���Q�[o�5����'2{�š=<�6�zM��zdUG�3D�(o�����\�7G�Pڶ�����1$�����&�6�|��J��P��]~{�az̴���7w�F�]��*�0�#ό	�χBҫ�T%|��g>��f9�xE����]�f��@�
��������z���Ln�_X�^�BL>�4p6�d
�3F��p`��j�+�wz�;�!(9tp0�ww�����g/�{� �7������z���Ej��a�?e��*����$���y�q��w�!ϐSÅ����C�d�2�I���0J��������N�=�E\���\�`�c�'��y�7è�����7:5<ц�o����?oA[��j��.�!j��;3��S=  ��IDAT��d�ա�d�C���N�l��\4ܨ������_�r�t��+ܧ=fT�2�!3���o�9H<~5q�7� EiYa���ok?�����=u����6��]���׽>��>u���\
��U%K�}��57oN��L<U���h�;t��~���'�<�6n\����a�u�}�Hݷ\?��Q�����vm5W���͜53:������6?����׍�3�tևB��13wN[0a�;gaD��`���&(�a��Y�B	Q��8�c\ĭQIĂ�5��=�o���ĉC�4&�byg3�`�6t҃�,"/����CX+��hoz��oK#_=
�	�c�'B	��o(f�1*�:�}$�H4�s`,-$��Q�iՓO�xϠ�� LCIǕu�81e�I)�R�#q|! �z����WB�B&���A�� \�-?J�[7�tC
K�^91��j�>�H.e���S�yY�z��~x��9#���T��-�����$�g�Y��	yU�sӦ��{��N�F1�ܘ�j8D�����\(��b�2j��N/+B�J�Gh B�n 0*�q���1�[�k��,H�3�<WvƢ���am9�V���z>�V@Y�W<�~����@X����Ҿ����?v>��q�sf��ر-��P���,|��-=�2%��vw䀸�������hS
Nop׮ڮP@h���&S@z���4y��v)��!!�E�._S#��椧FO�h�y���2�P���Q4�}2��c������A���v���]��gz�[A�ޫ�(3e@|#�J��p�vO٫��(!3�d&e���s2�{r����oH��X���EY��K�
ޚ��	>�ݴ��Smn���}��v�3)�V�����C�p��uda���Ocb��˓�j>�@����vE��� #�m��@�k���속Q��s�nxJ�P�.����p�����e"˕�������)+�� �@��]��R��� .F��3����[9�K�H?�:��8:��Wz�e��Q^�K��e˖�kkxGK;v��uk<����we�<�:�� �7^�1آH�.C�q�^� [�Gs\sͺvպ5��l�0j�a�eQ�����<��U����+����fϙ�����"��L+���kR�!

��ƪ�.��Pa�#t�-.���n-�ͧ(�J��3{��l�hD�'J�͑=�����L�<�J��x��ګS�>A�%=�ȣѐ<5!(�/�FM�@�1���f�:��-_��N��翐��+�ɺ���lʞ�ၠ,�[<̅��bPPL:Ȭ��@<8 ĸ��͈�|.]��-�RƐ� +@Կ��b��{�j&�_!P|���ܕJ�'�����}��<t�@����\�zE�4���<V�0,����)0�o��(�� "l��p���v��m����Q���Pb�0��0	�����YLOQ&����g�Qڄ��z���!��W\����V��3��~C���^)P/%�*��{!�h��K��|�����1��h���9*QF4Ѝ	�6��>�N@��i�S�M��?�#�v�'-��o4(����������(�S�'�a��t/ĸ�\�xπ�{�?�'OmC�F���m'l�w�X��㇗�<��0��ۘ?~����&t2��]��S�F
�Y���W��`�j�j�?���hDz�|�(?�P;�F�ދ+OJm�=�u
u,�1�k;|���� g}��#�>��O�,�|>�2�R�84�������E�T5�Z�ǈ��۶o�}��A<d�&O�����K�؃A����͛mSJ�����h�g�Ȳ���@<:�*����h�"��˼��s��,�A�Y��VH��z�\d�T��.�C����'37���Q9Q<t5+�1�J�A�#���v����t��]m١M��)�\V91�n���fц����'���a��y[�s_n9p�7�������󬘻<��|EFY}$�VY�{��z&t٪��0������m�/_���o6Уx��7ov[�vu��c��0lrN����yz5��5�@( �)���c�RG�:D#����X��������K�UW��>����h�f�A�cŒS�	gC<&3j㽌#+?,�~�;��V^�*�.H\�1���7����+B�+F0�W,L��;a_�o��(�$h�H��Q`
��~�>���������G��,yy X0��`��1�M���D��ȳ�1����{n��Ӄ $(09aDY�º��00y땗��˪)1�L��e�gc�}N�1�;�xszYRp�w)D8�-���ad]q��[�F(Z���;�ȼȄ�4�g�/y�G�2�Lu@o�&�f�a��e@8깩�^��^�4�oA��m���B�� (�`�����Q���Oz��gÿ�^#��L�V�M�n��Y!���9Gu��2Qf�iI;�Hon��>�P����	C��;�N$?�/3;�e�V_��j�rn�8�Vg1l��31��x�f���L�2hlM�V�
�u8����,��C�%�QwtVJdv�)Z���^�	x)�ƹ"*��{��Jn�Zx�8x|W-��΃4����?ī��C��1������m�q��7�7eؠa��,�z�=���9dk�,�v��k�LZ�vm�M�v�ٕ��v��@ܜʗ�_�S��ݛ�1E�/��94�P8'���^9}�������%oR����^]���U��@���{�秼��zƌ�)G<[�je9��[���4N�3��Q&��@�S�߅_e�Q2<Јx�V�p�s�"�K/xt}� ���W�RW�QNe&k����+�P�O��!nmdH�=y-m�Zu@?poH�gev�in�G�[�lN}i˅9!�E��d���_q�a_��2N��gV��k��M��s��t��m�����hj_�]��K�7gf���6nhL�4�_��/p�0��Tc"��ˍ���MYC�A|��	�L�b�.H�Mp����;7F/����8��e���9kXx����ݢ,���f߅y�'C���B��1�x���S��yjPt�l�[BGϺ{�� 0�a^������C��?��(K߬	`���K�0�����aW���>��U�A(��z�Z�+�֜J��C�a~eQo@�k#�f,]��A9'{����$\������<g?m���¨�2$y,ATw�q��3��+�H �MA���Oa�;��Yu�pŌ��x�0����p6R�GZ�U�۲5󲒃pVw���j_������� Bg�h�lB��� �'���!t�Ϳ�7�ڈ�bA��#q��-Z�^�?��+ �c�Y=�[P��7�;J�Q����²w�l�'h� �}a4W��<zZKÀ�=�-ȱ{�J����:��s5+��F����#�M�=����}C���L��;�65�!Ч>��'��#���k�|2�p4��X��7&[��#G��ɼ<�om��g���(3�d%���mtm��m�j톔;p�^@�a��ߺ�Y�~P��%x'6�0�߂�������:���O[ ��s���1\�S�-ă_�iK��SO?�t�k�shY���G�K��g���a�h7m`n�m��&�ǅ7��M�X�r��g�y�k�����׾>�����;ߞ�7�K�Cɢ�T����z���Qʔ�}�c�#�H�#^r�㫯�:=�GF�È����2G���v�ӴuFyU�CO�=��i�Z�XW�,��ƾ6�uEMp����C _��0��\
d�<ᙬ�Yⓧ:���1V?��������4�m�/3h�'��E�^=u$�\<����F3�݄?t
��N�<4[Ce+C�:�m1!�O�șB�[�^,�^����X��u���\��\$r�=�iχ��Oٯj\��0v�F�fntn�-�����{5���P�S�QD�Q5�F�w9�6@�.�NC�rO�ށ�ѫ<~4�-�/�P����x��m�PϲT�fe��� �#S�3���W�B��.�e�_5�k�cy�(p�1���N2Kԭ�	�8P��cq*���;x�0�<�9�/��ih��>�C�K����C�ڽ6}{r�	W�|�]�5a��O�x�#��P�Wgؼ����o��譹a�?�g�<�G���f�����5X���q��3d&g]x���W�۶놼��`HwE}6{���2D��bb)=i�Oe����GOh�\(���Bsn~��~,�2��<eH�k���-yWe�.U�
UO�0y ��3��-&M%L܄ci��m��.�u�D;q�p����m��`�;'T��CO�SjОhz�O<�d{葇"<ܾ����o|�[��̙U�߾��Ϸ���ߵ���j�'��$��?��?i�����?���W���?�W�3����/~�}9��':!OG;�F���Ʃg��#�!E	��뭌b��Ӭ;~x����a>��6E�&��:����?:��:W������(��P4��m�w�7�7�N������x�<�9�O�m[��PO[��h5ґ��pQ��*���S����ȈU'��s�^j��>d�N���ޟ
5�*�S�ޮ�)��r�S��+>y̓�oWҧ,�	oS�<l�ǐ9@�H�G��ed�J��sr]~��	��q���Ad�<Jv�{��z�-<�pTxs�+�:�I�|0lG8�g2�?���i��t#-��M�)>�ro�aQO �����j���RO��HdX�PN�	㕣?�n�uSȹ���(m1���t���Q�ia��Io�Q~�>�"�iǢ�:7��ӄ�x{�������,ޤ@$��\,^2�����j�%��h 
�  (5�D�p�pM\џċ �9�a="��(��4��Q<!�ܷ�"sELz�Μ�m�f{XX�8iҔ��/]�,��X>��S�4z�Q~�F���s-�� �"��9?��3�4K�"`�щ��������'� rL��"xϵ������\���
pR�		�$L'=�K�3b=�B��&�.Z|Y[xqo�������Ɩ�u�x�Mك3�A�Q�'�z��������0lûF!땤�4}j�i(�$�Eo%��7�Bc�2h%���C{>��ޟx���9x���K:hS��E P�Ⱦ����f�Y�zu[�dI�eq֋�K���WNy�}B��W@GYϨs��#���4T"��)�ݏ�,�t���!�uk��5W�n��<�x��5hJC�Ӧ������Ӆ�`�W�g;I4�˓������u2Y/�#�ۆj}"����)�����D��G���#�1����|�p<�r�ekaC��>�5��X�0'�a��h)7��gVmz2d��`ؘ!/���SCp>���/���0�:��xF��$��k��Y�Z-䷠=�#�jR��7����.��=�-�-���B�]A�l��ȶ��jM�i�D;Q�h%E	��}��E(�t��ܧ��(��.��ڌ�˛�?�8��u�wRF5dŐ��׾��x��y�=��o����կ~-�W�7���v��w%�1x�|�_K��-u���F�H����7S>:C��6W|���oe>�7/<)hH����_����/>���)��|�kQ��ڎ����ᵗ���M)o�喦��x>8,}�Όy�F��*�iI�I���7:��Y����{�w���/%�ȫ������:����xo��Gߓ�ʊv��S[1,��(�Z'�N�<1�cT'd� �S�?�[��x۷��~.���{Bv�δ�eO�)mՕ��>5C~��i��C�v�=�B�pl~��脎?:��Y��Ȋ�O��m�W�!1B��F�a�D��f�l��ވ	��@5Ta�OK7�@� �;��j@�n�=�ND�t&"+,vnߙ�`�.���k¨�#�ĸ>���5��P@L���w���[o�4�ɺp�vցgH\��mo{�Y��Qļ�U?ƀ��F;ap�
#���������l�Ew�ĥ�0Q	h8�o	�����٢��ex"��o��;���f��!8��ƨ1.#AԻ�zS����OF;��!�׾�59��%���4j(WJW:�P7zF^}2�w�)2\6~s=:8&����-�X���5l����2�`�ʕI��:(`�hVY��m�3t��s�y����h�,�8%W:��|�&h�gnԋҥؤ1)�δi��kek��3��˗F;^ޖ,��֮^�֭��ky�@�ؙw2E�Ԡ鉁�I�2&��~��K3(�nߖ4c>���Ю��6�3Td�ȩ�AM���G���N��|d���˖'�e̊6<���I�z�<j�猨۵׮k�-��ۻ;�9b �p:�{j(�	'�Qu:7�C���z�A;6���dA�r(�:q|;�+;���~:���rn�~���m���~g�̚%����'�O�y@�0���/��^uŪvUE �e��h7;a�	����r�O�F�(�4hNc#�e�2�`jл����C�/�K1�>�2���)c��+��o=����;2�7E�IǊqc#;��:��R৞z2���~ʪ�'���u�磏G�G���� �U���m�I�8Oj�@�u~�mD~; r�<v'O�_��W2�n���Y�c�]a哭�����Α՗��U�R���~�9<^���[ӻ������d�����x�"C)�M���9]C.3�z�F�P)9��e��y��~.�)�������M����ur�J�\��e@����'�ܖ�}���U�̳�s�xB�&�Ң3��M��iO>�tf۲�
��a%)�I�p���T�ꫯ:_��h�����?�\�lRı������hr�����z.�>oAR�Z����w���	��\
Ft�����K1���\h5w��KEw��l��7�y�ָ7s�H6���҈ٴqS{"�̄3�X�GS ��dZ���g�i{���l�gY�ګlx7+(f��� ���B�+�� ~���f��}M�����&�껺�ߋ�	p_��	pZ�\�/w���r襺�E`$�-���$����:H9��ú����bǘ�We�Y����	����M�X.#��b�D>��ތ'+��۽�22q�$/A��D݀�3,�E�C���>C�_��>��!�\��o A���w��:x%ԅ��P���w��=i�0���/��|��)���x}xY(�u!@Lv�'��^��v��7�"��m�x���oeze���k��[rc���\ޖ.��/��̛�q*"��K��5�͞1�M6�/p�K?���<.�96��s�X�fӶ�P�6yB�~]���w��0*��Ȍߧکc�DF�Ea�_��b�_�#f�D<=۩�̡6sʤ�&��sf�A�5�8q\z^_��;m�S�y���:m1���6F��`��=�<;�GC�I�i��]�]�ھ�;��#Ω6i��6o�Ķ`Δ0�ƇP���B`�M���mo{�[��~c�:�z�W��o��p]���]�zw��[r�c\���2[s�����cmnKr�?��h�Om$��������m����Kڤ�a�G�oS���KP�h����)ڃ�Ɗ.ޗ|���tu0y%7濼���z����u���1���eÌ|L����I�)"YguMu�Ȉ������C7��٨3�Ӿ�_5��WK1ƭ�1���aT"癵M�z�z*�)B����|
ǌ��}�a�|*�ۘ�� ��Ķ�y��iĐA'Ok��&O'O����ԝǔ��3��.��������;�F�(��-}�g����Ů�/d�:d�����N��WG�0pN�<�
΀���<�c��M�B�D;>
>�w{�8�"t:�0>���ɓ���l��E��ۮ��q�d�|&p��͛37�Rh7ç:6��:$P�2\2�1�<��F�B��B�� �`LQ��;�Gcn�]m_x�.���JEĒg��A�����V$�9��q"�p������>�c$W������|�JK�_'�3�`74$e��ԍ�6V�[q啫C v��O��f՝�U��\06(�}㹐��%`���&��Q��B� ���A�u����1Ѝ�`��ޅ1|i��9JV>���M��;�?�=XuK��p��Px�����2������r�=S�T�p��U��E0ش����YGsi��&,R@<����S!�H=ke����N\o�p��"T	~�9���F�<zi�������{]~��Җ�4>?���ɗpe�Jo���rڹ9�6�ksߝ|����>��O~�gۻ�����7�.�mm͕W�(m[�=z�a�N���|����Y3�P�MID�����]�'�ߠSR�q���hs�2�z�j����vK(��ో/rJ0#1�&�z:h��y<z�[���6��!^�ө�9��f�̆�Tl
�z*��ٳ��'E��{c�<�Dg%�C���CN
�SV��T}xkx2�ŉ��Fx�D;u�p��d�;���<A��=���z��a�\�ͻ�ug���������5���[sSFraժ+�Gh�B�h�\)|�x7\i�ޞ�oQM�,˥��y�	��Cއa�iCg��~k~?{�6>h9�?ZxY���=Z�n�U1��xЙ�eP�U2����W(�w�o����M�����	�M�f�n8�t���aP����癤t���ߏ=W�sC���~0�����/�&����~)(�(S�+/ƕ�vƅ!�/|�i0���-���?����y�߸��謼�}�Kމ���>��rM�a�r�}���� %��=o�%����2��m���oޕ-8�<���Oҝ1cV�E?*�t���F1��￿�n��d��/T=�Y<�@ͭF�6_�Lv�x�����0�/�"�Jݴ�kNψ:�ڽzpI��"bq~bE��	$rB�桀!�����G@�8T� ������A�j|���㒳����gr��HǊ�#�L�<���B�!zd,�ݻ{^6b��'��d�A��n �U��H)t�h|��~����\ed¬�x����\��L���)�W})��E7�u�I�� ʝr5��Y��jy f����g��
m�]k<\҅7`)o7L�o�T.�JK�_���ֽ�%Y}�[xʖ�,�Lz�������sW�6�_���s?�s!�>�=e�uEp���c$�~�7~��������?�Oy������}�K_�=\�EYM$T�A����Dv6��UA;+�g6��^0n�.[�8�PQ�Ya�/^�W��^��ܜ�Ր��a�4�Þ�Q��m_��\�iʤ0t�!-�u6��`�u:���!�ַ�����FM��m4:p�)r����̳��>Ҟݰ��߸��|v��ߎ��6kv|9��>t�}��_i_��۸h�����5a�J�>eB�6!��qaČ
Cd\�<�{#��!"��^�BxFIr�C+,��-^���0���8�N��u&©�G�w�d�im�es�e�93��B�ԐA'����K��9Q��n�øYm�(ڂ�b�\�m�o�7�
�A�v�,=5Y���Γ�0m�mWF�Ǥ�����}�=��!g=pF��m�îe>h�b�A�����+>+|^�����o�u���u-0/���U:O��>�c���p�����)?rF�g���7m��������3��L�6��m���?���_���<�[geu�©�޳w_{��'�`�;:ޱD}z��uïAeGGe8��`v��;^�۟o=�p��bzAG����_�rƶߩ�&G����"�38#e�I���<i�=��SϘv�%�woژܶ�ו�J�
�mۖ4�z�.g��a����߯.\�!Q EdO�\å�r��)6Q�/��	6����}�!JXc=z��ܱ�=�ԓ!p7� ���3o�2��� F��J�{��KIG�r���M<�p��2
(�r#�"��ׯ�:H��4�^"C������+~���w�P��a�/~�9IN(p�a��o�f�X�ll��t1P�,��a�9'�W��)��WY)?m���}�k�+�Q�xn�Xc�<=�Ki��*�������X�	��Ss��+o���w6�H[�x2&�#y���Dȓ���=�3��M	m��l����y���Y����w�h��lX������?�����ɛS }=7��V�h�*����ƛ^��%(@^8t��`��Ԑ�ԩ�rތ�*沘�r6��!F�fƲ �f�M�1�o'�.NM�	��IC��n|���Ń6��n�%�/Cb�ٻ�7tb�C>gB�2tV��������!$��fL0��X9q<:a�[E�ѳ:yf���������G�>�-.A����c�ږM[rۄvl��0ah0Ll��c�@Q~�Q�����M ��`N��>=B��Cl}R���I��D����C�,�:q���9�������i3ڂ药�������KG�薁c�yj&��ؘ;樐 ����?�"�o�!"p83jڟ�z�٧S��z�;��=����r~e�h(��z0�Ѻ�X��[_�WG��
���\^(�8x���;a��4����P�+���
�)�y_�FТ��_��ͦh��w�-o}K����P�9����}�k_�xg��K�V��w��5t����Qe�����
t�S�'�|��%��Qzh�T�#N��Ё�q������-�lD~ё�����.�����R�ؐ�dcto~Y�\d��A�r�N�?�n�K#�ᒀC$E�@�B��ЫN� pm�F^�
��1S�eh�J��Б-�#l���hh��8�ܦ:�IX'Z~<�M	!�@�>��W�e2�����\v��HP[���[/�'4����r��}�=оm�0�>}f���Rx�aI˄����N�_� *��Ð1a�9-p�RF��iЄ`����!��=��W�x�L(�g�ʍ	G�c2t�:����>�c�@��쀲�6�}0�]�kЃ9+���.ݣ�T�lҖVM�S�{.���+F�o�l	��'�FRYG ���jT2=������Ĩ ��dm��վ6��?���}�S�̺�>�(��3e�AݨQv�Loڲ�/��=|�
-�2(�v#y �E���x�p�¶b�6c��6nhb�w�?�;8k
�s�5'���0Q&�Q?��ŋ3�áLM�ay[)x�б�w��0��*=;=�S!O�	+H�x�k���GD
'N�m�B���t�ܙxwL�|�P�8iz��o|�ܜm����Dc����d%̑ڧ�BrȥӻOF�@��ޱ91)�+a���F޴)3���e��߄����9�h������ڬ�ss�X�39w�>�7��P(a���sA�;��hO<�d�7hC�mR(��KNAgD0��
%2�D������Cx>�|lNx(z�&l�A�R�=<Ά&	�z���y�e��⛞�f<����H���*������_0Xf����Y���<eqs�l���'p�4�jC�H��+��Ƴ�
����=�xC�{:M͙3oX�E�<h��a+2<
�|,9���C{魉k����)G�Ü�fH2ϐ��SZ�FfQ^�>���*��D�ʃ����Kf�Y���]�c�2� ��$�yᖎ�V���2��t#���|���Co�K �	Xz�WȀ,�����(�bNFw��L<�����@;�a���w xX�;B!0��F�\��>w�԰��(埓N��C ̾�����q���Oey����+*e��o���Z��;�ƿ|FQ�[�γY(B�q�3Lb��
c���iT��胁���n������*��=����p���p�<pԫ��)L�����wkG������������x���H`��d��e��(F�����ӹ:�����/SJ����vo��M��&e���P&is�CJ�w�~}���}�S��qk�+C����P��YC�%4���U�����z�C�+zV��۔���ӫ;l���=��P��ٜ�Γ���y��`߳�`۲u{���'%.�3;��D�?��(�ɓ4���M<x�8dO��14>�K��A+:�^�i�ԃ�NY�MF4�on�>����0O3��w�G�G���s"��?zhr�������m�֝�XD5v|>-��O���c#^��>iYc��m��F���t��C��А�e��uZ|69��6o��$4��QY�}��0��c���]{��9�2�L[8�q�'-[6��QۡqF����E���RpQ���*s7h�#�"0B.2Pu�����@Q���6K��n�嗧���0�r�5��my��鯠��f仗�-�O��@};�{��7��z?�[�=��YM>������B0O^x��b��Q6�#�D��^G[<�`��(�:9n_�=a|=�e;Z���>�C�VoU=�m�6#=81�FV�dH[=�<D��Η��apk]�GD'�|Б*���� 6�/>�|�b�W�D!��Q�P���Z�}-����)7gϞ�r��J>��%*�4��<Z,����X%��Wɗ�f��U�K��@�FD����--6��3�2ZnU�����aa��r�y��5;�2hLb#<�Z�y��ڶ��;�P�!�|�{��졮��3x�"������y�Un�Aa#�3��0�㖣�L�c�������w�m���ߵ�~���.��D�Ú���c��ِ��<Ed�7��}'��#��ӛD�<z��[��`n큰�;�0N���tCE�7<��T9	z=V�9N���2R�S/��M	�0��U��ܹ�����3�T&��(J��s@y�_N��)b|��c�&/�c'P8��lҕ�$���t��6�'��C�W�i䩿�˯�ʯ����{���᪽�[:�i��-F:����$ݢ{8���NPV�An��Nl�e���P�K/�ɷ7nʺY!d��3�͝b�۲-�fuȾDҳ"İ�)T�]�<t��xj^u7dz�9z�=���?���Cm�歡���G욫���Y����0V�3a���^(��^Ĥ�(O
��rUE7�>��b؈��8
~!έ ���5k�i�v���{`�ٛgڴ0VaЌ��v>���'��8�}����p�e<�(3����[_��rb����5p�/���p����	(��3�GF!��Ї��.��)���;��&ߒmp�'�?�2^pcPwWV*�[��aeq2����e��yكhN(��A�������F��-�,�bU��A��r0�b�}/鍄A9�R��
Pwx,9+$=K���B�סc�{��0F�P�B}+����"��!O~�+G_���4���Gx��{�IynU�������ߵ������lzx��xN�/9d����k�kW��:�>�9䙠U��c>�LEy�~�R4ɓ#� .�Q2��!J���d*��}��V�-����}�����K�M1سow���z��3���/�+큠7��5��l�%�y���m��E�5�ߒ+�̭�3w~�<yxG�p!�_
��F���Q�� �r��,��`��)XJ5=5"@��k�YM� ��3�A�h@BR����E}"��`�tE�I[`kp�Р�p%�M�dp1jJ)/!��@����P@T-�;��A�ݻP�����j����Ѡ��!{g���1:q@q�d�;�;���Ի�A�-��˾,,j��s��\�2H��e�3�0 al��c6��0r���h5�g����:EB�)�F��*�G��/.&��zA��{Kb��|S �4��Ñ�£8^����oN��<�;�x�f���'ۿ�w�.��n���C}��P��;�פM�#l���O�U����G�yn���������3�:��2� �@��6�^�ф�	�
�`ܺ}G���<���<��C!P�K�ڷ�`��L&�!����<A��QF���ڤ�MᏐ�!gƤ?q��y�����(��6k֜�1�1��m��`��ݰ������'Ӿ��{%ⷶ�oț|&^\���0l�A��}�Cfl�9?��U���0�F�ѥ�L���#C	E���S�vG�����ɡ8NE2!�8yj�F㷾}w{v�ƶ��m���CY����}�m	�3����M��޶!��[��n�����o�.��bXu�ڤ�~�*��/���>�1c��*Y���T:H�Й�oB�m�	���9I�&2�J{��0fC�l
���1	t��e���H����W
���b�~�i^^*��a��U�*���w5�LŃxW�W�/&/���Ӗ�v&�3� L�J�6U)�h��@����w2�Q)�������`���uߪ�O�5�����yt���rϽ��l��*W���H��W�L��3P?�GQ.qxjN���u��j��ء��E�7}���E���%KS�"��>�C��IFY��M�1�?��/d�
�0��m��(t��D�3m�L�Q�i��s��m�q.��o�$F��W\!��M05%�9�߿��CQX�&�:��$H�|c	�Ɋ��$�gyY7�ʐ�n��g}���z��F��[��c��ƻ����WV���s�N9���x6�"�zgCp�H��STL[ �Ap�Hy�@�z���A�V	�*� T^�"6q�WA�d�s�ڻ���4d|O�2x]�[��{�`a?n��ۿ�@~�.�M��#AX
~Y��|s��(R�#��`������EY>�r3
���P�:�v���)�G��(��m��~�?��m��D0�q3fЍ��I����#�	�6��( ��>)tR��\'Jײk��4�0ﵙ�M6' ZT��;=~=���>����jS�G~��=F4�w���S�<1<6;p��>�s�39�^{6�/dl��(lZ
�ciXٜnJN<;jL;tD��l|K��]�ׇ���"_�dQVw�ءXGڔ��X�О
��;*�w�F�~�Gu�]<� Mr�_��9]^��C��[Pf(�I���ys�۷�4��ۏe\*�/�G�n}"��Q�c9/e�U�>�0��޳�=����2��WYCqQ�,����8:<���'�����lV!1>~�0���m���F�vٴiCz�^��B{>ϜZ�v�ؙ)C�	̘���醉0�,'ߎ��8��Ɛ^y�Lv�uZ���p4J��M�*���/%
���o�
�Xx)Yt!��7��+;�O2j�΁��Ý�by1��w��O鐷���}�q|�|�/���9�����e��kB�H���wtxmu�Ө	cJ'����|���5�V�<��"ّq}/�^0�������T�S5�&c�m��B��������q9|m�{j&�������v�\��<i?^}x��������es¨�<=;'���_J����`LA��)��
�%�zfR�#N� ��}",Q�xOr�+~DbC5K�Ǝ!��Ĩ8�Cйj8WyV��QSSd�D�S��}���'�eyz�U�_�A��0�ag99���p eq-����z&�����u�R �o�<5�'�񜵯���1f��qrK|Vw{z'\��J�0F�Útk��t($+V^��*a���qÀгb�X��|y����R\�ʔ0� ���d_;���N]0����fxV�����k3��ԓ��V��W�ڞ����P����REed��h��{��	z�Cp��%ax���&ç<��e��7��С�UN�����A#/ƏaH����<FAI;Z`_|�(��(�)ȶ	��	��P��wt���0|�=���$�m�(۷S?��Xz&�A"ai�Ea�<�yC۱}s�a(�r zr�.Y"��1���w^|�/Pg��^wW��Ѩ(��~�Ϝh3�Nj��zc�����}��h�R^q�����N
O=^s^)
���}���0Ө6~��fB-ÁG�<�g�?���0�I�J�#x�F�|at��sR�'����s4hޭ.9�j'u��v���O��#��"�B/ک�}������#0h�s"���Z��:n.���d�G����Ƀ�>����[W�#=e��K�J�H���@�|�Ri��ߐ]��>��39$D^xn^�����W��*H��]C�=����0
���u�{Z��x����kZ��̙�A��sH�~T�|� ���{۪�/O	9��t	[L1ސ��{���Aӆ�x����_g�����w�Ln���]2�J�;v��6�-��	�hXy�	3c����i_���KF��{���Yvma�(y��Xt�:on5Q���*hR���WaN��o�W�@���������
�;��l���T`�h��!���7צ���W�+���M�ң�ΞթA���Z��d�=H��ǘy��_לtj��:�l����Z����䏄b�~嵰��
z;̔$&п����
��q���A��+�`��]i�����=�ˤGF�99��٧�3O?�J�!�����0=T�oNE�;�)yw&��/K����>����ũr1T�1ܓ`��n�g+bl��{a7��w���=�-i�Ք��|������=�9�����g�0:���A�����x5҈eIX
�@@WOyP��@�Ʀ�<p��@��{1��h���nx+M
��#x�-mW��׆qV.uF�'��v�B��p�db,������~4�e`<�eJ�(�F��{|��V�����d�ñc'��-[�OՕ�pἶ%�~��O�rhgq阘����D�y�#�h�˲���rU[{&��1�����M�6������ɓ�o�AxbP-C��=q2�&E����AE�=j��ɠ�0��-Hk'��J���Ė��7=וP䛼�夃��q�X�c�M��s:ޓ��xO+��dN��r�Eu����|R��`<�W��U�=9x�wt�2��QK�d�:� ���͆}<�j?$<�L��@����e⌄��՞��~��/��w�]&�]��/���_x>'��?��wJ��\9��"��D)��3����:��Fc�|�}���z.��3�(S�//�w�Qcަy5d�E$��]!�o������]u�'�;a�ޞKT����0W�t`N	��0�ݚ�G�^�l�p��9�G���p>t=y*������5W�^��v�}�K_��{6�[�hA{::`&۫�9;�d�7Vz����;7��i3"�26/���OxU<5��>��Q�p(X�̠A��t���4 �#�@�0aH�D4���Q߫�O�46h��Ҡ,T��®� M�(]� ���N�:%̱t�~#�"#E΅ ���ԙ.78��w�UO^(2	W�h0CA/׋�Ti��{y�ϻ�.��J����1������m~�3b��nX�!{������q�����I�ah۷o�ޅ N@��q`�|���bNFC���k?�p�V}�����K��O?�l�����1��#���b�;�ȍm��FqrK�y����S�'����6��1���b囥����BXݦ=�W�Bo�X�`u 4��=�ޓe+�Æa�=C��wF�~m����}��H�:Ek�.Ѭ/2JC��I����垧��?�]���J�jSϻ1��01R�A`�=������K�`;��x�?#��M\�8=|(��
�IA��ڞ]{rh̙Mk���-�?�=�c[{&��X��-^�$��*5��Q�AW\�!�R�^�MΒ�PLbR�`|9+��}a�?��Oj���ns��o��/h�	܈?>xr��~>���!Ҋ�&]N����'
g�И4j��ؼqs{��=i��3�lB~���y���l7j2dC/m��?����2��g�t>v�g�N�����o����������c�0��r�*�G�ӷHbB։�[YV��.9����ލqK�H��`�#�{�q[�_
�u�x�ϴ:H:
���dw����|VP��n޻�om]F�4�习4�v��0�F��(�YЁs�S|#�J� �ǀ&��Sc��g�H�=��N<��9�����ܤz��>U��	û+5@%𣓒�y^���K`cg:�Q�>R�Q���@Tu��x����W,i��]�.�x��}z��F�U��C+���w��(˄F7�͜9�-]��͞;�͛�0�SL����p���5����H�ұ����4'���D ."�»�կ=&��cԀ���O�ӸJ���}1�ȹ�ц�ȉ{�D�/�ߜ
̋`��	��x�}6O$�JAg �V7��\!�w���
!�,��i����A��ʫ`����~bܸ�(�0t^����yDN+������O}�:J�u�,�� �a�!3L�4�t���mZF�|���b�g#��a�<d�����e����8���vg{�{��y�;#�#5��(售r�S�pb����¸b0��0d���hDygx[|�������^��C�<\�%�;�RSg8*��\�m�m��F]�N��H8�N�)��t���v}�Mp ����0�<���M��0�8&�~s���}{��8���be�7gN4۷?���Z?=����k'����"���e��E&tt�-�z��ܸ��}���8eK�	c���Aks,��mF�1��h���|}DR�c��q�1��8nB_5g��c����(��;w�p�2h
(�F��U�����!/���f�~�C����z7T{B�@(������*�M�]<I#���_8��*-p�����;�c���oxpE?�޿Ҵ�oK�o�o�lLZ� �"�o��'�SߐK�2��JS���L'i���{�#cN9�C�k��!�,x(e�cu̙#Ü�/M��Ώ��Qj�����u��3���&��a�xǆ�w���㊚�#��(���K��̯3��_�j�������mh����O����A�x���9�#��67:&���h���W.�Q�W���0��Q�H��Y��96�^,A�j���a6z�Bo�Nt�]�� A��6[�U=&z���=}�6o�Ҿs�]��@��E܃���z�+J\���{���4�t���w��|72��+V��:0hxl��ZsUΏ��1�s���y+���殈�F��x}�<�\{`jw?�4GH�0��a�w�qG*W�at�H���om�}�kr�`�I<���ݩSӘ�^"AOGچw&=���6)\�	�PVt����/��G���'Ca>��4`ƌv%�e)��
���u,�`�z6��4������s���h�%K��CQoF"�iNx1����dͩ�۶������y-k4�u���3yx�9�ɧ�i��G��`l;5*��6�l��Qz���Ked;���N��3�$��3E�Z��Ú��غ}kS���1`��� ��:Wg�S��2�����sx�\��<Z�V�k�(T�^���������2�_~���P�.lˑ ���e�|G~W�*ޏ�,�˼���u����*�
F��J�w#ˣ܃�/���8%K�Jڈi���L�8_���C-%'�\�;���ry�$|DΔ��yӢ�/*'�D&���N�>9���0`�IÆ���i���!��g-��[5��x!�<�2��i���b8_���;�4�bhZsV\���p���Q]�C�_���ۖ-�7g[���-[ڡ�![��#744�͚=9���/\r�0�fD���}5���PՐ`�#B�Jy����èt�Qz!5"/���wu�/���U�HK�<7�
�`�?n���sz�yf �<���m�a	��GB��]�J���~�U|P��w#��ܷ@YL�q0TDi�P��6��b+<X��@ap���&HSz�7���[��42�'�c����-� ��� ^���Q�|���O�T^�dM�0pL<�Q>�J�?Q.��hI��T�.=&�g� �k�}8U>����0�S�Ջ�Q�VI1���4(T�A��
�;A��<��}���Ǎ���'��3��C'�Fm&ö�b�h�WH8�<�I�&�Y3�����|��A�&���˛=̨��T��L�6�͜37縜	c�!sJ8k���f��,n��[O{��;3��9�,�|�؂�Q��ͦx��r;y"��S��9kj�%�ڔ���}vT�Ҍog�q�!'AF��U�;�*S�+���6�_�1�]{��*PQ���p�~���T{V�~aYYPy���z�r�sa8���?6�,n\+��p!x�w���u���'��??������ٟm����~��~.���O}<�Yq���?���W�����g靉�'F�ѽ<�`��^~rH��<1+=�9�A"k�Xed%��ٳ���k��R�o��1s��)]Q���
�Յ��8��]���({ׇF;J���Rv�"2�sG�����b�0����2(���pI<5*X�w)B�Ƀ�5�I��_A!R�i+'8E��
  �ʫ�q$x�R�@g޳�ɸ��Ϙ������=�r�@��_����U>@����|�ag��J�`�����5Ƃ�H<�uQ87Lc�A08��cn���x�x(��;˞�P�qa����vE��eԸjgF�<y�|/0�xK�0��ɀQ&i�'��Ï����r��J'��}���DBLZ��t�<��W{^���p�!~�O�0f@��7x?�~�A���z1}y&�6���;m��b��`^�q�}̘q8��%�����QEok��9m���с��Ӟ��w�]�`a���;uo޴1�*�g��O=�LO(���:"
��,�����4�E/sht�g�bKXǏ��i3gE���g���aB?�������]?��Zib%�zh�&�}��]/��M8w��	���ip�@d㷹?FLo�~��P�N�1����o��B��Ş_,�W
��H|^9��0_�F�_�����rP߸���|=�P9F�)���a��8p�1s��7��Z��3�Cl�\y�u�����|#�D��+@�<�Sm�av�$2U��[�g2ѳ�{�Fs!���D.���H_|��T�@��3�}�wu�=��ȉQυ��kֵ�˗f�w�uot�M��8#��;wg\"`\t>fΘ�V]��-\�(�#�_T7�"�,�����[��K�QR� ��oa~����?�����O�~&S��V6�@�q4N)0�� ���}�۱�ҙ1{z��_����w�����ۿ���6':��\��3n��癍���um���i80�ԥ��U����g5w'��פc��Wi��qL�7�*�*oJ��#T�*��]m(x����[���3�8UW��q�MT����������,�﫾U�*��������B�	������y�=2]�{����e���%�i D\�h=���@��ψ�����?��n��~��'���(��s�X�4w���-}��d���߾�}��{�\����jM{���o�뙇UI��y��g����D4��0(��SѮ�`<��(�2&��Q�c��	Jl�'F�Mh��l�O���'�+�\����j۞���ƽ���鉞LC��2�ӑ���'v����͝2������\��h��|�L:)p����Q�j�n�|7�����0�6�
���jǺ������1Pi����~0_�F>��@����o�|9_���t*]r���i�14�+��aup��ZhR�/��l#�����ש�Jn�G%{�]y��|�#?��_���ٟ�Y�1���\��n�)<�d��m[�`ڝHr����8e�?(����NO��� |�]v�C&�O_�w����G��^{S��G���7���m�����i���7�����ի�ӹ�=��S��	G�jژ�,jo��׵���~4w���W.���G��"�bh��+gqz� 	.�Z�K�f��}�����.�U^..������	�EO/"�������Y�J�a|��(����JI�#�`���π)%���?��������9��1(<T����+OP����Z9�Q⊁���V��x&��~�A�\�P9dq�|��(O�U�d��h@�hQ��IL�:�M�6�M�J,�I�VP�ʻ���H���p1|7��ߠ~�W~#i ]��Z��r[���X +��9e��"ꬍ���~�7���J{���~;#͠�x�4�0�SX��Μ:�l��|�J��mv���Bxڏ�����ؑCm�Sm�����5�ڭ�_ݮ���Ѿ���S�ۘ�����G�fcߚ�C菉��3�˻�;�w�y�/��Z	p풸��l<��P�<�|�����F���	8�&M��2\?�z���@��/_�?�{λ�o��1W�+����NK�׭�ӑ�0Jq�aLe,�,~��m<����#a�N���[i�S��102��� \(��|�i)G��G��+MO�
� m���|g�����\������l�o߾#:�w��_�җ�g?��ܝ|Ϟݙ�o� �lt֍B�gF$ȸ�
@����Cc��EC�8�͐��#ǚMM�m��;g~���H^T@���%�a�鱠��>�����w`j�f?y|���蹓�~[h�,e6tLO�mA�`�+�t�+/X��{5ỹ����4�
��9�9;�?�@��x" ���8��s�,H��i�Q�C���|.�^����.���5�Q6������9@�G����;��;��0פ13�MV�~�lHU�*�4K���%
�%�
Ua�Y�Uq+������S�LQ~�(��=@2h(?����x���4����H���	������/���V���_<�/�9s��4f����)��k�h��9��	ż���W�-��6�nH1O����.hkW_�n�����w�ٮ���x}��߷��:����1��Xt�D(�xp6z�g��`��963f��h��(��5�b�i���#��ێ�[�����;1hF����0X���p�G��MM�te�xt8�l�
�PO�ׄc�lt��D|�Or]�6��#>�|��0��Ccڄ�˄�äPs*���/_�n���v�m��dW�m�V,mKq��	��.�V����ڌ����B	�|bz�Mc�3r�E�����
o[!�G�W�7)��atXm����hb��.���/��K��Te���,���J_��0��:�~���P����������{�7������h����~��~���o�fzV8��c����6<m��'�K�{�V~�F/:'����t��a��H`gsF �I�bqG�>��H(��d�	�ى�N�Q���4^������]�C��1c���a; ��a�G��鴜ټ�PX����Xu�ꍚ�9�VhH�5@�߿�}74�{��:�������#���ye��BD#������ ~�S 0�f�������9aY��G�iV��U�Q�kR����F���
)"�ߙf�0�]���=�WA�δ��~?��ba�~�}�qA��\=���eL��HH�E@OEC��/����/
*/�}����ګ֦��o|C{�[�ȱ|��~��|�Mm��%!,fe�o�e�㛾!$�g��+CYߖ���~���M�{m(�7������|Y��f�r�a��m^��DB'�e9�����౓9WO������s�̣r���/�����?��1��-F���lk|�qAk㣎_cl��yVܻF�C���v�h_bn�˫׭���N�	�"pT�X�՞j�w�n�������h���ax̟3�����f��mr���啚�ʕ�V��/w�o�営n��ve�sI'�	da��6+�4�ܶ`�\�"�o�[nl�|�;�����h�w押����yԈ������aڢ|e� }����w�bϿ�p��v�,���܃�������y%�5��Ձ�������_�e��^���ghj�'>��,��v����E��d2��>*z÷���h � �)�[�+�;驃��"���e�J����������]ȉ�ğ2�x�HƸ0no�|��L�n�Y��Ne1Y_��Q���ĨH����GPqJ��,�/���-�NcyW�3�T���{_3��o�耥\a�������sp@ձ����Vߨ�w�o7����cД!���w婀�J��WfCuQރ�TA�u�0z^�~W�#�z%(;|&��0�h����GB�(�\�L�6�o_*��p����`~���U+��|ǝ�'����n���<�N�Β�ݳ\�Z����o����'�n����[nm�W_�K�[�.��5��V�)�&�������Z�ha[F��SsY��Ǔ!���"B�H�1:��ŋ�@��+�/��������c'ژISڄ)3��ӡ��G3V(��^&����0c��ð>qɀgΞ���	�5��Ү�vM�4y\;z�5L�	��Ԏ=���au�pSAˑd��#�Pa�̉^┉ڤPsgMo�͟��0�v ������y횫�j+._�fM������+�F�cQ.ݽ�0Nn���	<��be��ʕ�������kڍ���+�H���M)"m�[c_��[�$�9�+ŵ��`��� �����w��r֯���0�������v��%Ou��k�e�sb,�0�Q��1h�2���y�Ƿt\�g�!���G��|S��T���L���e��e�%�4L@Α�PD�N���� so%���ˁ�G��99ʐ�H��_\����6e���)�N����6����0j��
���C�*� �#ҹL�\����@ Ԍ�Ӹ	���C�UO�׈�L�r����J�-{����W�r��v8�j���6*�I����:r�`�>�+�$�5�%�z�'8����eQL� �=qi�w9�=����P��0�W���K=�}��:��w/Ҩt�]����q_y��c���a��6�m�^����gA�1���8UV���*_���?�8�)�I�?����O�I{�[�H75Z�ǂ�D�h�/�M7ޘÏoy�[ۇ?������oh��|S��p�Į�;#��63��5r�=A�'��0N�ϝ�shl�5zt�����*�S�>!�ds�+?=��G��c��.�Lo���-;v��[������i3f�������S�(K���N�3��`:}*���N�q_G�9Y7�gN��MeG��'��g�y*���@Ci��0):@g#��0�Ʒ�����P:�,�q��Ʉ�=�^��a�̍:�É�G�<��x?O���Ƕ��m[6眡[o�!��k�x�������I��x���u�^����mw�
�y�愲��|���x�1"�>�H��i�ndc�V�6��js4� ���ы�+����K�[t��R���0\�����ndx)�~�n~��J��Οgޕ�C����^2���Cڍ���l�Q�cy^:m��^=>Ƚ^"_��AlR�2���/i�۷��Q��ԛ�����ww5A����B�U�ĉ���� �{��]*:�+��m'G��g+����xĵ��~S���s��Ȓ\Z8�%.1V�AD�O�u�8��f'�X�`a�Ü��"�Ap/�"������P��]"N����<c��'���ZcECE��1B����^Y���f���-kA��V?�˨q/ �9#�U<Dk)��+W����)���)YV���(���z�Rx|���U�V42x?���T��P��>�
�P�s((q§�M�o�8+�/�X~����v� ׮/��=�v�=�ȏ|����wF�~U���0�k7�tc��[�S���ŋ���lW���]�zu8W�U+W��W,�g������������ڑC�׳aLD����EY�M��	e|*zmCAwCa�E��J#41&ӎ����m�ƭ���6uZ2q�"zaGڄI�ںu׵���{����Ϸ�^����;��n{��ڔY�����"4U��)S���a��:��D���Eo6��#�L>��϶G��>cV[�tY�?���wH^!���=��M��=�\еd?�J�B��x~w{��'����Z�s<�l���x2?h���mu�r���m�es���f��K�Q4)���_�v�7�e�s���Y��m���������S_��׶;�xs�a�w�=��<���V���ӫ�gE߃�re��K����*�`���k��ε�f�m�S^����B��Ԑ��n.
���%�Ԟ�6Rf(�F'-������ s��,r̘��z:�_�hq�ohk׮KOг�>��Oc�ȺV�;��3���x'�r�x��	��@��/���=��t�*Q�Z��p[���<ǋu$��oD
Ǘś�/` �W	.�QSDBѳ8)�A0ࢢ(x�A�լ̱�?ВHِ&2�x��p�T�E$~g����9{6� ġqV�����b�`�l��nV�(C7�#m���C�)T��O��O�_��_i?��?�L�ɀt��}=�n���@�*�ۢW���s�WU�^�?�!�8�pS���]���u_��=��� ��0*�zW�]�u3�L���Jc��>=���0$�3�GϞQ��-���u��V����w�%m���7^�������z��;k1l�,Y�+ޜٔ���'��t�Ά03�`ޜ�vB�&�`̸���:c���Ț��q��Fo����'����x8yDw xЎ����}�`;z�t	&#�0o>�P��M`t��SO?Ӟۺ�=������9�&�`t�
��}�=�D7f���<j����a`Z�d	��(�����Lh3f�i���<E��Ç��Ç���ē� ��V;l(���.'�	:�U��A{&�.`�
��_�<wVa����c�cڌiz��e�1#�5N�_�6�gW^�w��n���ks�
sr��2|�v�U�k֥�Z�3H��w�A�})x��>��{�e�_�Jx��+����"�,���;�l��nw�������MFs$u(����Gս��QiF����g���&֞<�6���/���c�c�T7���#�9w�7?��Q��36����G�����]ҝt�c#�G���4m��2V��`�a�%����n~	��K-��Qط�@۷goz`��\]�X�V*��^5�$FM!���PC�����[��䰍]b5N|��s��}	jŏT��h_��Ze��������=�a�L<c܄����� ��D�d��fpk���<�<�K��=�ɣL0���Ҩ2W���%�,O�v��9�2B^!i������
�p1����.
.��bA�*\���g����R��+�����<��X5���`p87��K5Ǎ�%;T:�&�Ǒy�z��� ��<���V�.�m�����}&��8���cGBXYr�w�ܑ���u�a��0��.n3g����&��Y��TiG|0��q�=xƎ��0[�%͎����z���D�&�aٷow۴q}{���׿���d\�x�a��īr6:È��Q���'B����-�).wu��hx��Ķ{���®=�t a���f�J��7�Zu�0Ə�øe�&]�|��H'���hb�{Jy�^tNi'�iΞ;�M�:��܏�F�!2��'L���0%@���`�®=���m[�#�<��z=�����R{�Ʒ��;<kؒQE���W��G���
�
�p�g��g#��}����ȃl�3l��ӍW|s�5״��j���?�[k2l�����v���?�;����Ӧ�Xы�;}�UP�S���)YR�B��:�V`�?;>|�5I����t�2'c��if���Q�~�$�S0c�$�����.0���&����fUT�u*�'ӈ2��ޔ^���L_fR�>mw��}�N��2���1��H�K�0u��r<.�3���r�
 Y��v���3i���J������M@=Lw$D[D�>q̲�z��o�<�5{]{ڈp��DP��Q�*��#�}�|\�����댒a�y���sA���+��Ba�_�
���_00\.��`�݅�|WWe�0�}����3��ߐF��E��g�L��Λ�fx��28�$�
�z7X�2>�~�7G�I�?f��}�ǅqrWs�6lؘ�4D[�����x������t�Pϟ��͙� �k��✧c'��B�8�P��Q&���(���u6v�9��/�H#����-���콻�o�����6}�6+���������-o+�,��m��%mi�8:�nI���]�	��2c�0&e{�_g���9_h��Y焬�X�Ȉq��!4���M��(��!PMT�01��0Z�L�٦L�>�ٵ�`;x1�64qJ;x�D��x;|�x�ͩv�h�;���n�c��6;�7�SO=1<qs_�x1���M�����o��֑*ɻ�\J
��]JPV ��傋����o*�gd^�b0��+��2��v3G�6#�U�j�mwޙ+uB����}��yq��G��nY?z�>�!��vE����J��F �(xUy�r���J���l�v^i;��N:c,(��}����z�^^���ʨ����]�@��\}��(S0F�B������!�j��'�Eyt:���b�ø��(�����䘄NL�6B��ڽ2=�bpO(P��r���)��"�
,М3�ّ�����ZFT��D���w�)B�+���}��d�����耽��K��׿��=)�F�W��ŇIXʫ.zhk��}eX���������R�*/�HP*�ݓY���qi�|�X���#��|0z�}�>(C�V��$�&/"旂�y�^Y@�����/�i��k����z?�ld>���ۅ�g�.����>.�7ܘʖa�N�L0��|����Y���3=�}$�ʾP�[�l��B��A�l�g��{��x������<�|�ވ�o�z~W����B�HK&���m�^���=�Ҁ?!����ٛ;p�@��ǎ

���Ѷ~�s9��2�ٳg��2'�����%����s��a�+V,k˗-�\�V�\�V��"Wi�gr��+#����魒�o��x�l���t��Hn�e��c�9\s��ׄ��8�@ X���D+�SF��b����pK�frv�9�����?��{���0�Lj
������3��o��u���{מ�O�a������qs��t���m����֮�ac�·x��}��6�ok�ַo~�[ў/��������h�BPtT�A��ρJo$Գz?��G�idx�Pq]+͑P�
ܿ�p!(�I�x�`�2�ֈE'TGI��`��������x�d�O}�S��]��;y�<�{�)o��6wμ���y��W���|o�)��Y�U����Ə ]�ȿ���tj��i`Ƿ���U��C8|������+(���ڶbՊ0`��'�=��Smڔ��ѱ�k{Ȱ���S�mG�"�߂�=�M�<-��v�������KvJ7�`�)���[p�H�:+�Q�-��i�Fh�j ��`IC"�ݲuK��Y�g�#yB��jH�G:E�D	C��h����v�u״�Ӧ�|�o}�[mK("�5�=H�דL�abu#��І��x��TN�N-��d׹�+�ckmid�9��Apjvg��T�6���{�ct4�h)H�O�����Nz�O�b�A(F��+|!ƾ�m��'���R���[x��
��B�N*����^�žWW�#`���m�M)(���6M���.�Y����<FB�yhB9yg�J R�Lz��!���h���>�h����y(�'�7�x���P����=qoϮ&궳�v�����u	ك���ad�߄�ۤ��ܤ
�}(�1j��=�6�>toHńj��,Z8����A�'�9�&eYy#���&��!8삿O����+cxpr���a��o�1<�#c^>6N{�[=z�⅊ȝP��x�<�yD�1��$_�}�w�wi6nl�7nj[����<�Уm��-��s�����@0���2;O>�T�x�u�>����3mNtZkz��A���:��r��7���1�� ]����K���\�N�W�.܎��*�˕w.W~U~�+���0����RО��=��6G�pz�n^ޚ�K�ũ��;W页O~�������t�ӵ�����F���k_��6���\���ۡc�	�����f������Jn�S�{G�+�j�
(_ћE-��%@� 
�a+�#����.�iЛn�>',���u׽�7�&NJ�8�A�j�(V���4j��9Ad�0���2j ���􄛆���A8͟7/�==��3)���H�/�� �F��]�Jv:�%H���@Ҭt�*=���Fº�AN�����W�=��9޸t!�7�O��N�\�CO�*���m޵n�t�&��^�����;S�<	G�*!��C��[�Ae�~c�p[�_�;��%��|G��a�M�;�0&��8�m���;�Ɗ�1P�U ?i�)O��4�7}�Q���oA^��p<��e��3V��z�ז �?�[2��(.Z2h�Zů��[�P��� ���8�5'�C@8�(gya���PH�y�.AJ >�����i�=�X*�͛7���{v_���)��(��}8�l֝As4+�.�lq�q\��s)�V��'�1ah�艣���<z�T����s)4�\<m��\n������^����N˞��Dzc3f�q�Ɣ4>xa���)�h�os|L�eġ{blyRB�&=�XL/Z@c&0��ϻ��N2ڂvv���x=.�(�k�tm�����3Ϧ��q���cASv���n���P"&?�'OȐ���ot���ݾu[���3�HrJ��!�g}��a0�]�)���{2}�.*����0gd�*��P|y1x%�\/V�����܏|�L��U�N��#�>X���@�K�����ې<���!�U�@�U{�����7c��{����s�'C�E�iD���d1��a(8f�,�y����͝Ψq`0Pg+�@����-��<�>x��!����(�y'����x�����{x���,X��o��]�����?����ǞJ2q�P��� ��16�\����6͚97�:!l��.�QSD���JqR&ϝ�����|E���Ӑ�=�֐PƏ� ����{��E��J��F���@o�w�¨��>����_��WR���e�K�x��Ҷ�o�^�4MHe�xf�0+V�)y1~Y�����Xі����to�������⏲/�t��^�Qco��,
K��k�ch��S�P<?�MfՋ�˖B0\0+�aѢ���K������X�V�Ý3gv�{��˲<�.Ð�#_=�Ya��	�Wg�����G�z�������۬x?�oE���͂#�ԃw*/�d{F�&բ���h[B��G[��gwL�1x��}	P�r_q�OŁcqz����[~�!0�C�%$z��㏆�ܘ�Li�D٭�0�t��T��VY���8�D GB��8km��W�EO*q?S��಩��=�~������0h�~fC擓�ǎ	�Sxǚ%��;-Ƣe�&Ԛ�{��)�)*�tB��_���{����+�c�a4�h���T����a|�#�a���P�a߾����� �="΄�E*��0�և1�;͛8ó�Ј���d��;n~�����2��@��q����;Sn=���Tf�O������a���h��m��ޗ����S���Pϒ7���c�Bߎ|�|�O�
���A����|Vq�:�O=ĕgE�`0�
#��-}��0�y�N|���:#�>�@�Q��s�Dv��M� s����!�I�=�L�*:3Jz�����՟9sv�����)�T��䩓Sv�):�O�e�Obr�;���&[�������fжUT�x��(/���˖/m7�rS���O<�z���/�Pځ��/�鰙g5C!���:��3{n�o�su��������M@ixʅ`F�������O��O�o��od��{=�|��6\��^7��!�A�ᤕ[F�#�)�I!�<�@��W�� �j��˿�>�������{�����/�k����ۙ�g��	��'l���3/�r��?����=�rˣ�.�?G�z���}|�;�0����������{�B���7��<>{��������s���UP��M2���)܃���%`@L	�:xp�ա��O�|x����j������ܨ� =���+V��+��y�ӷ�ҲC=u�Y����{���u��[V�X�%���$��{RH����� 3t3s�~�В�FB =$q�8Վ{�H.�V������%��H�[&|�[�������.k���n��Ԑ���^���ou�ތ��/�8��ۤ���	3O$� #�O��
��L0(7唖k��o�q�p��~P�a	F�\��0�+�[m��{p��y�(^2�H�
M���x��)�: p9��s�+^�������-�m�ЄIͤܜS����k{�ц�nͦx>!�ɓƇ��8����{RX�=m�&��I�l�!�(�&����2�>.�n�1�7�kIO5Ɩ�������hOF~�#�ˈb|�Ĥ�Ma��(��M��%(��L-���0y��Ӳ����_ˡ_��y����E'�!%�0�b�"JZ��z�p��W�[ϴAom������4PtPao -tZtS�y�پ��Է�|��xW�
�+zV��������u_e�͐@ůt�{at����}ݏ�8�s�2�-}�q<�=YMn�@�`��\A�:PҪ�5�C&�B�e�ډ��2iPG�}:���e?�?�^��׷E������~�73�j�G�!hP~:{�![��1Ew��<��}���g�%��W�]�SW|K�c����x�킇yb�V<�i��������/}a[����������mڰ)	�[�&��ΰ��#���vܱ����=�}̱�cVD�~y��C���{���5Ԑj  /�:v���~w��@��4������t�����=�����㪑�O��`�^!�7ٖu,�x�4�wێ-�~�������67,�[Ê~�￳}�������vR�HtN_����a)�a&��e"��'>؍��T�](v�TFF 9D}7�r��xa�`F��Q����������˞�`ū;��S��ԃ�������FvW�
ϔ�I�V�8/�ao�O�<���v��'�7���U���d��6��B�Uf���6J�Ż��q�w���W����L������V$��PےWOZz�R_D��
F��{�����uD'��H>�<��ă�s����N�z!�G�t n��>B���H��q�,�B��$z��mz��W��&��>6A/v^��07dor�#�F�(B�'�-i'�|B[~ؒ0'4�^g�"}�7��oh�0����ʒk�=�ȘPӳ�¸�|���i����&c��ob�!�o�)�[K�7�a�^0�o���Ɏge����Y��!w���σ��&��E�:#��u��U[J(�=or�Hu�w��#���ޖ�6p��hI;���s�Pei������X�w��H|�F��/(~/��0MP<���EK��t�잕��L�*��x�� J@��U\iy�^�C�|+}@6ƃ��|*ݽ�W�*_ū��;�}dU�N)O�H��i� ��O9�t�"�|��5���K�;�u���n˝�������W��͛�0�r�W�W�W���%��8����&����T̨!��]��|t$WǷ�z�qǥ~��/~�9�����B��*�zm���<�#��Z2�Ka�����^�}/^_����l��������9�k:��yx�7�O8�͜3�q��yd�q��NXqb;d񲨵v,/:�@$c�(�2�h��A5�xI����Sr(������hX.�9a��#;<��}|Oɔѓ�4M9�Ͳ�x_~@�J���c�i�����t҉�ǵi�x�6� z~��s_XNQ��!�C ��#��(�O��}��`WO��:2P%]����#fF˗����^�̡��G>����h�_w�n�d����<�М��OidĻ�1���S|N��g���5���[�q�y�ܜu�,0bV^m!�����\���Cc(=	�\�;�����>$p.O��q��9��50�� ��!n+��7��W\�4c��oʛ���3����4�;��{1���vy�~(=N�41����Uo�q�>�-c�1f��2B�eo��S�a��#YF
0d������Mo��sYG�^��s�҈�;���NP�Y3f������}���6>�1s�pKZ.nb/r�+��s�h��1m���A�'�0~���Lщ�{4s�]��������N^�0�3=ۤz��U�<{\U=����n�����DC��c���P���P  �7�HT;y�wKݜ]�-~�u�'}� -/�;A���M�>q���p�x2�'����t�D ��yA�����e`��������6*�W�R�EpYú9�"��Uq�P���[�ZJ�O�^څ�W^~�����;o��er��O�K�l2�a��Yrhȏ�=�.>���v:��
XQj�/��zO�'w4n��E�����Q�_�C�Y����3��s��ܝ������#!w�3�~��3fg�������QM|7GS̜>�=��m�#�9e}O���a��=|�:���y�3�s��S�� �.�Щb�l۹�-�q�ig�F����?(:�'�zR[��0�ŗ\ޮ��l{j<����91!:NS'��ҹsmJ�Ƞ9����R���SSP��G"t�C�C(˘��ۿ���я~$�bg�O$��9��c�����mjG����ʘ�`��m�ޖ
�H�����qJZ���/B1aDJ��<�fu{�ӟ����7�ys�����j�������u�<��������]���έ;��f��!�'N���B<� �#e���E>��޹"�/7�gH�ώ	��"L�,��Bq[~˅�>��� �᧟���J��K���{0 ������s������7������ٰa}0������)p������{�Ƈ������S�	8eֻ�l�KT���p5�0~�t�Z6��oo7�tS��c�i朌a��'�rJ��_��,��������?���SO?-�M�9kv!Pv�\�W�3RL"���_�j�����Y��eUZdH�=�b��n�-'����%�w��{8�̚.���<'\K)���Ǐ1c��c$N��{o7�c)�ަh(�O�[^�%aܽ�ok�.[B���Jp1Z�(��u�1^�G��0!:�D[Y�7�->D}�l3gL��W����~�5m���uz�Y��4��v���&戮�:���w�dڎGF&|3����c+.r>O�~��Cڼ�3r8h������"^-��d<6�|����ر%�;(]�vK������>��O�q='�9i�Q��.�G�êy$к1�&˸��v迬ӫIC0�����N��z[�I��h����s�y�>�4���� ��œ����P�ɫ����{�̈́�\u��ެD:9��m�۰67l�o2Dۘ����䪞�H/�nԹ2Գ$Fvz��o��+�M�6#���o>��?�k��^��<m���^��c�XtF/���r�
��+�W���ss=��v4lI>괉G/���toC��'��!?������������ݓ��Yu8~���s��~��9��C�ߓe}׻�il�q�44#�a�5|с�N��Yz�I'g�ؙdd��=xk����d�"���&�[a�k�G�8����g=;���0d���?�S��?�֐k[۟��_���c���͙��D����@�s;q�ü,�qǭh+V��]rXT�w�z8��5�VC�,Yʕ����������?���&���vs�Ԟ~�32E�h��P }�!��b�tf�#.q��������'�{DW
H<����������׶W��a�_����~�����i?��׷e�/O�����پJϬ��s���|Ӣ.z5A n=P�yv�"Re|���`�m��</��~0�W��+�9ŵ.�d�n�x&���@��������?�ޛ��w�wr��<b"�3f�/ޑG�=�NX���,�U8W_uu�=�F���^BE�g��mr@]��p T����k�%�S����{7؄|�3�n_��3߭�s����y86��Yal�����������i�|���_���dGOsZN~ø�d��ʒx!���� ��C"���$���p@8�J��� ���<N���	�Prat�%���F�*XDK��!e�^BDO!��/![��Dz�p9#��#?��� �� �'�����B�^�3����Ia�O
#}|6ӧMmS�=6nܐޞAK<=�*�Z�v��}BYL�:=$�C�*����S܉�&����l�N��M�7%��0f���b��9i�~r�ź���Ag��X�4v�a�P�a�i��(ǘl��������g>��0�V��X�����};�>P�C}Q�@h7G��i�x��C�eܬM���w�{�����.�g4h�z���B�e5� zy���a����[�)�V}Wq����Z��9�[2�6�l2�Ί�S�l�{���c�ss�xr��Ż�������߇�������r�����8#|����a��c蠻ܒ �nFW ^��	����.�r�E^os�4��� >
׀,x��1w&�}��o~���~>�߫oc #���Xzw�2�\���0�$���Gv6tE3'�xR��_��v���i�
�Ї>�����,y��lr�����Όc����u_���S�.Z�8��9|�03�a�Nr��]�"���)�{�Mtǳ�ٱ�|��y����O�_�����w�{�[rۇ?��?l����o{��pt:t&̩;���l����g�͉y^�b�OiԀK���᧾�Ɍp�A�B`)O���o�)Lq��3BX�zɾј���K���������x+4,oţ�h0y���8)��kL�KۤQL�{.�O|����=����Le|xS��wߕD<3�&����(�, H\>xQ{�s��[l���/��!c��,۶|�Q	N�d ��+@Yb
�p�go2�bS��� $DX��G�ꋈ1F%$1'/�1Yq/��ɕF��� _��/Z�0�25{tʃ���������n��vw(�����r��"w�G��P���3��/��-=��_(ﾻ�=+�iw�qg��/[�8о�=��itQ��+ˢ�����uOW�0Y|��m_���������
u����ia8�.\=����k�{ɽ��/ɝD7h��m�j'�bD�����<��Z- �S����L^
��4�F@�G���o�7]��(�ƈ�Ξ3�ݿ*h'��x·һ孁�-aT�/W��i�ӌb���!�y�h�g���mL������<���={N�X�� �s2ѩ�-���o�yn����.T~
�I���B�ݸ2J��dӿ�sggz��ĦE�r�;ɛ��
��	^�	�AS��&����ꤛMa��P�ydA���I1�3��'�{�����z��!>�]1��3:t�k�=���gC�,:(�ˋBր2J"R���PF�Pq랂���|�Zr@�un���{J��K/L�ΙUx��q{����#50��0
7m�4Ɖ	�x7!դ�������!���ǯ8.k5jC�iEgL�ݛ�%����v�&�l@�]y6x ���wpmn�J��x�,��n
?u5�{������I~��hn�) d��,׾9�99���'�{���F�������`�"?l�aXM���뮉N�E!ˍP��r��!~��^���Hwk�/mG(�Ud5>Vo�hs|fd��������������h��lݜR�l޼=�n/�:i\���K⛙��(�'�q�d�n�ᦔap̛�a��:kִ�|鲶(�i���#Os��lA��n��� ���i �C�*��l��z�����+�M)��I� ��y�e� ��(Y��;
�&VI�3KR��ԡ���_>��d��$t���_��\�@�F)6���E緼M��$��!�)žJP]���*�(P�4Wġ������c����{�1��.y�1�:���<� ���9�~N�O ������ _���O?#�蛜�[��,�W����`tsV�N��%�z4�ӣ��^H�:���f��h��R�@g�!8�;�-��|�h ��b=ٞ���SBq�ޛ$j5��%{Fp����~�p��<�ox�a��Aq�)ݾ>z�4�ac�����A�4#@ݫ�>����B�����-�����7��'�2�"�$#��|��NP�Μ�L��65���o���F�ޮa3��͐Tމƶ9�t&Mth��6c��� ��E��ώ2������3��t�ļ0P�������'{�0�X]g8e����Bw|��[0Q`EC� Qݜ������O�!<�&���kV�ѳ3�2�e$����_J�����i�28=����s-
��F�g�]�W.Ϥ#�O�����W��o�ôШ+ܺJC<��)��7޻׹2�»�~���}o��r�����G?�.8�+it�Gޑ3z�V�hs���A����t^�é���N�N�3�qv�7�eu���F(��g�5eu���_���������O�}��_h_���y_:/x����^1x��+�p��C��$>G���̩�-�N��|<:��/{�4�s���Л��ӧ�c�t�x�L����Rv�G�潘�[Ƌ�5m����K>˟��+���~��Y^�hmR;��#�IeR���-pI��=�4�'|�#3���1��cLȃ�.�"�Ή�zZ�����S��⪔)3�3g̊��5y߆��C7-��w�G�oV7j��#�z��)�(��3J!h �=�~)��[�i(��ip�h A@"���FB4��GC����`L`*CSI<�b��[�#n���aS��S/�[q6o�<���{�
�tW������,���Hz�?��?�=f�W/q(�.����^�F�}[�P��K>�t�Ơ��V��G� p����9g��C�KOM|e����3o�W�$=�(j���b��H��U'�,�J���f�q�#i� �
�جw���<�F{�!�~F�^��e�V�}��k�}M���?<|��5��h��W��r��f�ϯ|�+)�M���S>cȽL�Ζ�kg�.hM*���'s��/|�ً�FO	44�z1m͠n�Umo��@�6W�=�������})�>�n|�5	�|�I9'��Z����1�N�H�i���G7�^~��w� �΋2=�y�CXO��F�g&!�����$��B�p^�b�0���f\��wE�W#
������w�3�=y],���mL(�q�ޒ��-1���6V>C���3[܋g#~6���;�"���v(�g�!��A�Gö�4}'�}�+�O�@�-�N3�h.}���8)��aiT��B�:uޡe�.0tL���y���?��}˭7eg�{#��ɠ�sl{�9�hg�qf�$r��o���mM����f)+��PI��ܜF�C�k~���+�O/�x7F}IO���x*�<���:�l�h��kSrO<^o���Q3���p��#��!+fi�Dw��W�m�j���vfz��4�#���</W����=й"�o��lw2��hV�VGF~S��/�$��,"�Փw����-�V�W}�|�]�&W19Fe�����w\��g?��8��4z.���vQ�śDoO�6泙�3���i�R7�t�`��6m��&�2
�
����R1[)
��1,����k*.HG�����t癸��Ƅ���� e0�0E�P��)ķ�!����������h2޸|����o}3'�	������B�����0*=哞�(�׽�uY~�ܒ&�Q��[��b�U���f��*(8��K��:7��t(7O�44j��P�H`����� �<�l7 �Qx8���c(�{

C�}����q��c�"�~z ώ�� �IρS�����N�S&����9r�����pzZ >�6�qɭ
�!�C��c!����WeZ���7ږh˓O9%��=5h���Dna^��p�M�/Z��6QW^9�����˿�y3v�F[�RZh��6�b�mʶ�i��fF#�) �O�1"��IS��8���i��'���C7@�+��Ƿ����L�09+�ˡKBy��;gN�1!�wLf�^f)��*���9	6�)z���yg�O�ܦN"��E��Ql^��4j́�U��/�6ն�Z�(R
��[=���Cty�l�<�(wzj"^�]!(ǵ0�(���-�]�uoOY�g@Y؏&��g��=26�c����Q������y�w���LH�ڞ<����I��0�d��NЛ�1����_Pwu��{���+������%����-
�p�駝����<�M���*�W�J�p1�c��m��w��7�3A�:3��!;���r����p�t�.7�N<@C'�5���o_��Ҷ&:��v�E��Z�[�!��y�aD�����Z�T�kC���9���AO������U9��!���WM>6λ�-�k�}�s��m�5�':��s�����[g .Lt֎�ld0���W�\9W��o<�{W���0d���|��l#�_r���g�C��`������s��̇g������f��V�^}�Ձ�����xG���&�i+���������x��Qc�ij���+�Hy��N8����.���F��pdg4x��)j坚��<�F��鳢��?f�t��@E��2�CQ�D�a�#C!B:�� �"0�b(֤�5�6Ƥ�RчR�7�/bw�!)�!P\BD ��-�
iIX�&;͝?/=5<��;}��$ʒ!�'O�����Y!x#��{o�G�7S=
�!c��&T��`���/�/﫮�*�MY��x�N�d���A��UP����y�7y��	qc�b���lB��
�pp�őm��ۭy0ད��B��{��!|�����v�����+�|)�`X������RCOk�>�&D�(h5�{G��Mm]D���xy���};�?1z^eԠ�jBC9ճa�cp1��x�޽�E/�v\�q(4��1�!���)!@p�-�?n{8��VFxYY����$&Bͽ�T�ϵG��^PN��m�3w���K=$��p�;�\�=?z�s��nV��ɜ�M%�;G���N�;�C.�ԧ�g�w�y�6-�00rA�f8DB���팚�C9>�������@Ѻ�!W����HG�W$A�z{ʅl'z��QcL�ayP���+/�T�1\�i��f
5����/n���;��#OG&?͞=3�Q�o���������ζ11�℣�>&i�B?$�no3ڴ�w�T C�ծ��/�߽�5�	����s��y�׼��px��Y�4y�������׼:�"^��;u?�=4�@���+�z뭷�o}��mvtb��"�{����P/y� �M��6��Ua0�i�󫕺P��D����h���v���O��	��<�]�F��F��&��:ש�>�f�ͶP�zֳ��Weg��xv��g�/��4j��(�ϴ�p'�T�W���K��}i����:��F�Qْr6hZ�v_u�隌#�u-F9t�Y'�,+0�I6�S�3��a�PCkʧ����1����(�H��_�	���MӉw�!�Ȯ*3���m;�]��L�n��Ƀ��<+��k�9��]|�彳�"sj]1nt<�A��9�_��8�6���#���{p aߜ�A����g��7dC$!o� ��K+��:G�k֬N�垴ĺFAM>��4�箻R�JG�1���3e�`���I�!�u����_�=��)� 1&���9���Ð��˝�O��4n|C (w�?+�޾w���Y��R��ޓ��D�%���T9���8��ƽf�R��
�/e�q������K�;cO�f�]v�J�`��.�g�uVW	�K��%I f���2vEfN��P��)s��`�6�>�ypGVH�c�P��?�vn�m��K<�#z�G�]���Оz�2`
̄������e�O3�;������^!�F}��d�l�<��@^<B��K^���A[�E��=#�?�Y�|0����N|?���Bޖ��sL(���8��q��a�B����s�ig�qj(�aH�Ck\�m��4'���x_x+�Й?ov[0N��s���0���Ǩ�xv��^���i1h#���ch�PVGJO(% ]��x����Q(@r!�м�4��v�����$��l+�JR1Ќ^�txy�L���������+�v[�uN;�أ?��c��=�e���>樨{���>4���ė��؎=��P��ۊ㏋�87���$���V�n)FZ֛e�kC���şCP� ]�|=3h�1be'��>/�W���)A36�|�k_���~ک�%����M�	��eb���sBf���y��0T�&�Q�q�Ө���I~��z��k�\�?"�ҳ����>�7=�{��x�0l���9+�<	.I���/e�%y��U��dՔ����_2�l=1>���E�����;�N{{xݽz��|�>��~6��ϻ���Åw�q����ψ��<˓��aY��&��N���`�t��Q����&W�m:���o��}咾�!�c�����Q�t66��Β��\�?��U��V޷[�qi�F�1R�Ogӑ[t�Nci�6�އ�Ҙ��=�t��uo�{td(\�wW���?���I�Y��`����aB.��?B��11�w��4@���P�W��P��{!�I4DSؐ4 F���]ZʁXįɺ��8}�T�l�k��E���%�x�ci{.}�g���Ɲ����`@�������L�@JH����^����x��x��~�<~{�^{�檡P��ٍ�{�*w��<�z����G��Nn��+����<%�����{ٴ���q9\H�e����d�Q.e����?�͊^���ɑ���2H��*oV��	t��������A��~|#��	*�_��>������_ۯ���@�:F�莑MH��6��:�o}�[۫�"	(eC{�C���X����^�������w���7���<眳�q��ٞ�^մi6ǋ��&GXA�>�� +��|�נШ�#Aoa�NZ��9	7�C>��3]B�%����N�z��rhl��al~@�At���h�=<�	���=k��A�:	�3�ޘx������ۀ�	ܙ_�SL�,h&�}��(�
* B��998��H�*Dt;w�믻�=�~m�g�qxک'�<���G�Gڋ^��4~�y�3ڳ�yN[��67�) G������2*x?~��8W9�0w�Y �[�����,0D����}u��9!�>�|�.��s��o�2�#IgBB'���o}���.��7�^yHn�)5�t6YM�	)�7cH}�6�o�D��8���S��<7\�h�0��3v��G���;sq��<�#��'��%q�G4������T�)Β�6��2�u���NB�׵�j�µ՚"���M�w����l�����
����������i��[��~�7{��3/{�K�LB�)���[I��7�+^\�&��U���su�V��4���=x�yhlg���HC��fi��|��)�k���0X�[7`���#�����O眭j��v{�i\�0�Ӈ!Cꠊ;#ڂ�W�![��,��o8���.p@���T�!�4���0I�Af
�@
$Ae�[�!��=�ȝwޑ������}4��G\B�\~j|J+�hX֫�:X�������4\���cME@xs��C��Qԭ�sc��]<�*OJ���7b,&��q��җ�4���*�M��b������;��7�2����x.�=C������]}L�R�`�܎U���c������G���ʤ�d�1}B���K&=7�2	/�_-�^���V��oϹ���=u뢗i|Z\��a�6���7��$4���ƤQ�:�D��G��^;�C�G��9���zl��x�>��&N�S}���(>
��
4�e��ǷeK��>-Gqx��̍0�dX��ӭyZ[��a���ˀo�G���u9�6BN��m�B:�<���adϙ��3�*��̥���a�02�-��{FO2Á�B����;(���O�+<��H\�������#��4hA�p�aQ(�]J;�R�����[B0�#C''G�NJ���Ƞ1o��m�4������َ=��(�x�`xN<3�d~�;���}Nh/~I_�o�J�O�{��Г��� ����3�Cx�_: ���J��~���������x<�z��9�/��j?��������M*����T������2�Mo���#7�Fi�M��#�J�gxttBq�@\ƌaP�sa����A2��>S��)]^�W��5�N�ܹ�x~A{嫾/��҃��_nb��\�hKߐ��,�G7%k�5y�����'���JCZh�s�o���<p��Pܥkx_���0�U����1hx���03d�g-�6\��y#�*e�0x��Κ=3�c�v���l�/PF�POu�����_� �I��>�Fn����F��4:ldiE ��|�|��C]�3�|;s��4�rZ�y��̯��KG�nN���|C{�k_�Gu�<<;�#�h�:D�#u��5DP�"��\�� �3O�;�1a��05�������\z�徴O���4��5 &$,*=�Z촪�1��U�P2�9	�1e�G吾����(���fN繘�ee���'?��=~/.����\�w�N\� e�n�Sw�cp�F��L?�����)�W ��CE�q��Y�-I�1��L=!B�%08L�Ġ٣Jc�T�pl(Fy�J����d�v����͒Y���7��1ϊ�Zٔ3?#>�B/��衚���ʍo�[-����oy�[�e��~�?���ɟlo{��r8��_��(�6����uy�髷�w�zE��Q~�Z�e�tC�O�v]�pQ
H�>x����0l��f��f.̎PrAe�50�Ü{L؜N��Dl9��CO3������ʘr�����Ｓ�H;T�+= ��9�+C�a�K��~�Ƌpz~�:e��;��Υ��%�m
�,O�w鮎6Ow<OM�[КBF��#��0��O��w����^Ӹ%�H�ٺv�*���V}�^^<�z�2��lOo�j��S$ߏ�ؙ4w��%�E��ŋB�-��>]<�]�%�H({|N�9^ŵ�mx��~�p��h0�u�E�����~�3�����V�	x>y��S��5_����o��ȋ2Ew�"����\"so�o*YV�Vj/���b`)�w�'?*m����3WP�3t.ԑ��#7�"��P�A�#^:2�G��dﾯ��v�uפ�Ń�L�{(K�I�T;�W7�y"��o�&�ΑQ�,�����U���ʎ�py�_�l�y�z\y'�U󶂠#��!��2��{���s�3�����[r��z�l�^�i,�[����5׶VG��)+�㱶:S�|�K.��C���d���	Ѯl0��\������8y��\����Jܪ`�)� � ��A�+�B�j�ٛ�@���,"ר�@*a�=7f�����¦<{���n�[okk֮	a��*Q.���/�$ݽ)$�A4x�&���B9�߼5�!kܱ�[%Ni��Ξ&Y!���q����Xټ���+��KE0B���,W�c���o��h�L�#qàѫ$��]�%�2B}0[�����Q�;���(/�x$�=��o�[�V]	�idirū��F��Y>ӆK]�愒�8�W�lf��u��0�e.��rVu���W�+r��],���~0��\��RG{�f}�s(�� �Q���vC��Dv��b�#u�E3����.w��o��+�n+*�(��*mj��{߄Ktg��aA��Ќ�4r�W;���`#�dhWۙ�N�C��l��\��*/�ũ��ͧ�<5h>x5ލ�3�da^�I9�7g3>�!�n�Z޽�mXo�H;Ԇ!�"R���)E�mKuᑡ'�Sk�G��.
طq�kd*�D��^o8����+eI���+���M	���$��18�e4oo�{h�H:�6�0��G�+xe�A�l'm�*���i��L��
�3i�mh� �0r����!����P)E�;��4Շ��C��������/}�KG�-��{#)<��g6�-<ޝv����
�6-xQ��\��߈$o��~��fTx����ʻ�\��gd�k�����$�o�"��F��V�B���[]z��׶�o�3����^�q����:�k=�o�U��������?��?���y�ϟ�ٟ�?��?�����O�,��������������]�M���*3j���?�zi'A%�@g����V�<�8���XY�CT�k�yߚS����'��P��"�o��C�l6�w�=��ǣC�m��0���C�.���W�����y9G�!��bMl��4tyC�
�{�B�S̨)�0�
����-�!��%0� �f�'�"F �$,;�Νc�dj|�~n��C� &�AX��D������6�,s3O���[��y_ȕ-��^���w�#��p,eMb��GߣE���9���-�D,�����
i�E��2��Q���� _� ���az<���~�=I��-��Ê�$(vB���J���� �.�7�]q�U�̐rϕ<!�\���[�@�eo!L�zY���]I�v�{�mW��*+#��_>?�n��(cu�����}o#IJWY��;�!��.&\)5�I����V���1�a9G"
��������e�I��g>�]��6�-}�K�~]�+1�Ӧv�UW���!٦�e�0r�j�5�L���v��ݯ��r�ݛ�nI�`c ��/��.
�������wn(�y9T��ض���vF~��.�!̶�l��D{�0[<߸)f���M�Bmێh�X�O&L����Ho|�����	ų+�N�'�u#KwM"ܒ�ax�`��iJ�7°q��΄�!ػP?(����b��D�2�u[�1���� �M��[�w3유��3ۢŇ���i�ܦϞ�'�u6�Z�ޞ��d<�:�!=QAÌ=
v�zCș('�):AVfr�;@��oj�_qi���a�:����*��j�K/�$�	�P�O:�49|�Sq]��Mz���{��2�_B� ߧ� ���7hO|�-��!N�1�ѳ8����'����͛x�l�!�0l#_�9+����.� ���E��0p���`��ر�ϽcE�널y�����L����0��3T��G�|C���r3@�h3������m�7>r@\x�2�C�^��;y3��]q��C�a#0`��o��_������|���/� z�{�2�+ٹ#C��t)~ou2��0D��}K�@��R:��r��dc��xo:�('��?�i�e��YF���Q�C戋\&L��K����hU:v	Ƨ�e	\������j#C�_����K/���4�������s���	�O<K�["�p��AJ�S��\sm���������A�te�H�*'�iѻƜ�tٍ!D�'8�L�H�	7A��X��D��)q��ꫭ��	x��vJ�E�#�����q�(D�;�5�:a�G��e�}<�X�9����(U�g#+C�-W��	�s/�	C )�)]�W����#��`�Z�K���巺XY��qU�7�@�]�PB��l�dHʩ����F�����j���.|G��T��an���0�KK^�M���\ np_��o���K�ۅ.��n��T6Qc�D�t�b�{�'���]v��Q�������[�K�� n�i]�Y�r�b?]X�̞��W*��m�)x&0ԁ {�ޟma8�|��0L�-]��H�.�ߺ�[q]���qY.o��>]�~�m�^������vC����@�4�[���wݙ���MmC��ʕ�{�[�e����tmRhb߆0~6D/=n���^�3�1���[�z}[���"�uA��R�oAA1�xO&L
��66�n[н9g�7u���жMz}��F,�Noꎗ���=���nM�K�9��D���X^ �?1:"z�ek(.֊+FY�i|��b�#���IS�X�զُ&�;m欠���9��(�Ckl��5ҞԦ���qc�M����\zYR�k�8�^]�d΃������=O�jc�R(�RL��N��P��E�o��'u�^�K���L&��N�b�G|g���\�����xd�oѪ��a�<͛����2�6��6<d�|u�mwT���I���XzL.�[gϥ�y\�NC��zL������ڢ���s_�C=�-[���x�A/��)'��r�������IA�&|����ۜy��Y��
͇�ٳZ��x�Un�8�,�Y�yV���;�%��a��B�� ,Y	oe@z�7|��5D?���`X2x}�&2���}t6�N�.��(��y��g�����3m��M��^6��~�>�@���j���)��a'm n:��&L�C�[��ѳ����!v���Gy��������0u۵�^�>���<N=��l��h�[�c�+T��m/a.�N
���{<�Q��S�xأ� `
���Dw�C+/>8�[$��O�?���uO����H�{W���\�6u����h���d]��tZ'(����~ �ҥ�۶��J��vv�ӣYܖ��RPNĪ��ߌ��~�#�� Q�c̘@gǏ���������?��oj?�3?�~��~.]�z��<9ܮh�a�6��!`a.�kA�R�@�p�l�:�{�ʫl}� A]}_�.A���}o�H�����\��m�Lq>=�U)�x�䫭��U~E��e�8�R��5̤���0���ƣu��[��=nܞv�%�K�pc3l/�������w���8dd��Ah*���u��bC(}ߖ����>!�{�������{K�O}�S�C�8�|�0QN.ƴA/���v�ŗ���}i�\�o}��*�{�ڻ��wѓ�����}�}��j���7�|�]u��!���Cx:I����3`S1����)��h�~�����ك�O��g�N��	�έQN����]!�l��$ ���C�w%Q�7���$���<�q��J�S\�?����&׻̎E<�������ׇ���{�0�o�\x�(͋�//\}���߾�}�_��n�-h���>W��]і,>4zڗ����}a�~9���nk}���\��>�:�!���y_�B::}�a�k:|�=< �H籠ɨ�%B�'w�~�5�`u(ykٱC4�0@ȓ?��?h��R��;F�y9p��h=����"D9����4jb��1ǽ���C��|�M0h�0h
/��������e��C�қ;f�����9�S����
[g`���m|`hjUY�!��F��v����U(ϙ��#�|�g?���gB��n�S���-D�<�̨bT����F
(��*�n��;��	>L��{�~����k���|5� ���r����.��=m�ڇ�u�0�!h;*��1i��|��rEd��>Y!���� F@���|�6V]:?�|�-��
8�V�$�;�(̧�4�3�=�-��[~ݝV�C8s��6'��CT��nJk����w����Fosu����9Yp�������zʖ�a>!!z��ѐ:g`D"�ˣ`s�q
߮Њ��7�ʧ>���'oĢwn���Fjv.��P�!�I�>��p��_
H�/��7�+��B4�O�(�t����d�(�������T�c������,�-ً�U+A���o���M�=�4����6wU&���Qq�!��z��ɤz��)��rfP��1S��u��0^�CK�s�.\�vtVw�JK/��eTHm�4:�z��׾.=B�'E�\�)�0��{_�)�r���jq�饞w��W_}Uz�(E m팱�uI����0X���/��|䟢��0��Wqw�?z�[��oܖ��=wߓ����&=o�~��ZvG�(����l:���9x����S�`��6/���x	Y����ͥ���}�C&�B?<jg��]�������]ڿl��^h)S�r�Y�{�3xR1��tX{����?@C�b��^�.�5Xm��\��\O��;�xS����x�g���e��ƛ���on�^ri���}�}�3���x�����\y=>��O��p{�_�{NW�ߩ(=>#K�u�8�>mg�c�eir��p%�6i+��v�/��� ��~��p��?��R�-�C�ϭU��ж�����wچ������5�!fg<Yt�ɧ���w�yG�<��}�xpי���D&���sה=����u$��b��<�uix�[�:�j)TrGG��1T�hk�u�����/���_񊆇e<wձ1��SN�y���r��ա�ƌ�b��FE��[�H�Y�$mϊN\�L��2"��o"M�yu�����#�&���I�Qw���(�3�a�e�/=zȊ�N���c����Rf�˾dJ�)O��J<�GD(�H���QS�%�Q!P���[�di�)� @��"�0CL��z ��	�I`��&N�&M1��Jw��H�2b�(T'��صɍi��=��(l�}�<B6���1���+~JԸ����&N�EL%�	��л#@xj���)L?����e�$��;�N
8�UY��+x�8�r6\#��0���g\��ƽ�r%R�\��h��Y�ކ��!��ʻ@���2F��uOq����ੱ[���rm��3�!b8�X��`p�#����p+= =���=L�3���#�ty�(F��:,������1?�#?�������7��9���4w��}N	�{��=���x^�L(�/����R*������\����]w�tpw���ڍ7���weж���aG��蜸i/��N�\�W^yu�?�v�j�5�e�Y�tnX���>3�c����� �mzJF�I�;�9f͚�_kB�_CJ��)}�BmR�=�V�R������	���O��tPi�����R�=Pt�3��������y$�4�,�x��kR����^���w�;n�;�o�oE���[B��M���#��;�t��]햛oI7<C���.o��օ��K/O7�!�k�4$��;o@�ſ�'A'�� 1F��{�߼;���P����ib�F�ٛ6$�[��dl�Kxw@�?��?��2:���u꺡`w�����C�zf�2K{P��Y�Ga
hY���0�~�]w�ЫRђv7Dk��+��2���;�C���]���4��8	���?֠\2�ś��uJc�#d=���	�랎�z��N�+Ra�^�U;��{p�~�uɬ���%;tz��.�?�@�s��K;���e\�Q���L�6U~e���-�M��H��d<ѝ�-X��6o��oJ9/��^o��+eж�X|g�(<�]���'b��m��oN�^:�w��ݧ؜�B��c��*���c�s�i�D��}
�R@)h�į�J������֐�	�I�!16�7��1�� ����TBFOZ�%�Qh�QG�N��Ғ���2��m����6!'=q�r�����L9�	�s���y�g�;g�X����ؚ�fq�R�z�&�Zfw��ʍ�;��$�U�/��@q����
���y%�������#J��t�chc��h�Ǒ�O��_�f}VJ�x��*^��P��F�Y&/-�*Ɣ�0�0��nEB��F�l\��[o��������=��=�Qf��qƙ����N���~� �x�D��K��΍�^��fnsG�ip�&��^[ͻ�xX�k��$b�K��s�����7�<�v]����fw�uOQ��!Ǡ��� ;�RY��7g�@2l�q���.�M�]�nC��y8���J&\R<�y�N�#cř;�ܼ3��h�=��$��`B�:1@L$�+mʀ�ҍ�
@�����#��[:�)1s�L�g����Սr�y ���(qiÏ '��NH��C��a@�#Bwʐ�"=�5���{�7�P�O�=a���T$�2B��<�G0��bWWA��A��!�2�pQ�8qE��,t,��=�;���p�+ށ/�O},�g�I��s�a�(�U~x�)#g��,�V��KEK#m8֑�MC��â���6�=��6g��,�!?�ó�t�]w�Ѯ����nI�����7�#���m.��׻�c�,�ɳ��(E�����B�d���ҙ�'0��p+�[��)���򐗎�����
�@{���=���{z�;���=+%�,c<��.>���ے�ț[o�%d�#A�v�i�\ �|cN����\-��H�����$]XH�PF<�w�[t� ���]������ЙaE�H"A}��i��`�p�����aH���T'��Z9���w����:.�NO���E<�X#����Da�z�'fB$�b&�); ��$諱 �[��g������S�k�h�4�g}X$0�iHgShTLX�)ᔀ`"@����2=�����˗��7G��&�+L%a��I�+PWybd�ϵ��D����L6����^�>�ֳ�̥���4��p���C!�-�/f ��* W�Ҽ�`q�^�0�kY�q�ù�2\�'��	�ŋ�^��+�pHgs��w��F���4Z<���	m�g��y��!��0Dz����xm�O��z��^\��d��
�$�Ա�Emge ����&��H��P&�3�B9P(p_�"���z��t^9�E�-_0�`�-@0�<Y�KЌ����tL1�e�8� ����h��r~Oѵv�����ۊ1K4��)Ƈ��v0v��|7>z8�䭨S��<�
E��QE1(�)�M�
�Y�g���6�)x��-5/��3�01x~�����D�*��vVN'	o��=<���-(�����S��qC�ݝ!v�l��,(����wh {��B�;=9Ϩ�᭾�C˥��4x'��'8��ߠ��w�Qg�lJ��k�MG��4��K_�R��G?�q�#?l��ַ�5���m�}��uŁk���i)����_�O��n�Uxa@�i��8m���^��\-e%wS��Q����u�r�`���Ky�s��ū�*/�����WX]�#�4�%�"�=h����j��ca�#F,� xzh��_��z7�$�M��p�y|d
ق_ܓ���^V�w�����U3֪��x�,X�i�Q�޴�UY�n /I����6�Y#�ד�K���d��)=���7t$�ΐ��S.N:�J�B.�(|m�I��׬�+���S2ub;"�:�lsBf�
�g?�q �5U	H�̂�(S� �p	O�:y[u����2"�Цc<1�/ed�=�N	�M����	�>¸&'"��U־'ΖT�*<4�4���.��פ�����P�FC4�۽��I )��`d�4��������|��A���2C@9(w+aN4�`��H��W ��y!� e���������<	"���W^�{�]��~c0+%~�}}���y�������U}	���@�������=�ළ�{A��{OW���lᭌF�����)J;����n��=T�f�/M�����������]v�e��+�L�G��������Y=�h�N(�6��G>�C�63C��p��C~�ה����0B����?���8h�>�AV� E�+�������d�77|�6�ҽݭ���"t!/��9���Q���Z�*qʊ�Շ��=%����S��h���s>���
�O��샢��ӹv��v����ۯ�{��K�v�H�Evr̝@��s>��Q?ϫ��y �}�ެS�L;p�b����p��)�'��t����~�W���{��=z�H�gD�����,�������VN�wC�½vG�<4:Je�W����X���y=tid��y�,��<io^�i3l�xP��2fc8ta/�x<���9Zr�W�V�q�p�{{6���vF�K��qPv;b��EZe�O�9�:��Xڼ�ʏw.���v[��!r�G���/���ݻq�����2�b��AÓb�d�!7���k0#�!*�ݓ�o�\C0]tqv��F�8x�a.��1LG��{�F���o�7�w�%{��;��3�S��{;�[�ƨ�[����r�)�3;۵��u�k��|D��i9��P���s�qA�����-^�%���?���#�C1и~3jX{�����D�&��w��_�bװ�f�� yf�������_��	,��������b�ux��8�̕	��d�(�#�9B=9���Ɛ˅! 0�98�B�#������N�������7FT6d 0{�<E��U�����{��S��VJ�ဉ�ߕS�rOhX6�c"8�W�ވ ��0g�X­���;����{R�0v��Y�!�a������)c�a���޾���w��������=0��3V?�!0� �'��ݒ�k���{2���g���Qr�g�2�(6�J9(P��n��Ɇ�������L'��d���>���En���RG�{N<w���ʓQ���M��j�ye�jW��Ao߃���o(���iqbD{���U>�1�ekS�������[�̉��QmhsS�=�P�"m�ܺQ�o�	E�8|���~5Ԉ:��N�Q����������nڦFӣ���.�v���9���Ð6T�w{oЦ���x̣1t���
`�������H~{m?����k7�rI��1�v���ږB�vs/-P�FC����<pD����}��߾J�v&�Au9uP�*/�_������2d����%�8`({���?�`H���/�}|{�ݎ��;;Q�O�(/�#{�Yu�qǶÏ8��8�<�cٲ�B�ӎ9Z8*�yc����?��u֙�q��i����|�I��4*���l�tH7�x�Mi�O��;̚5'�?���gL�ўi�-:�<&�D���͡�(�\�0�^��������~�7Z(�7o�!�2\�����;�>=(��:��;0��������!�x�y?ʨ����
r��Yއ|��H�����}:g�1(�w�z�_:�G�7����r���h{��@�\��+_���ɶL��3)=���5i���pἶ<t�M�ԭ}"B��G�h8���h�"�X��2�|9EC���J�{.���x�{\Z�]X����E>�wl=�4Ҵ)�>���a^`���h�L`��׍�Ý��F��}٥���o�!�ޘsY����[A���Wu*"��U9>����/����8�w��C@|�ܼus;�����]�M�nBe�TY:{9}èѳ�S���B�p��S3\ה��驜u�!�������t|l�b�f|W�G���4�����0�g������)$,#<d��vX
�e��a*�������O��{>'D��HEJ �A��]s�5��{N��w���C�(� �x4��� M�ũ�^	���R���cE�PD�Ջ�	v��� Pm �a;�n�졑���c�d~�k���hUC<ɸ�0�ҐI�;OJ�`�D�j�_�7M쓯�~4G��P2���:�Y���}hM���1����Ұ�����{��9�8x4]8�F�21bM��]Un�"�a�|������Hw{n�y��W�K.�"b�Q����^�蟢��{�����WƎ����6R��eh��˗�sAxN
Cz֬�iP�%��x|M�_P���[>0�
���|�Ӊ+�r3$;O�9j<���a;���бUNz��Rm!?��x�^C� }�:1h��h���s:|c"~.5��4/�����-�VGz�漐3�����z�X�-�ݐ[��AAV��������H�Qa�oټ5tŪv�UW�k��6;s+Wޛp��~X�G��������&�[U�X~ز|'.���o�U\��g��V{�9���h�>�dN�5��0 ����g���4�|�}y��9�'�w`z>�	{�q1�
�;ɡ�66�2�&Ҍ��g�}n:�1�n����������Q�k9�M�g��'A7�3oV;$�^�$���5/�qFp��5E8 �r�K��0;��7ǽ���L��ȣ#t�'��?�h.\�rk0���}��@�n"�\�7,x־�Լ�c��3*�gٰ��x�>G��~��m���SI��0m��S�\���T�^�.����U���Q�g�fn<YJB1��'�FM03��b�^o� +�����0	����$�L��k�&�y��<�iO1(��N<�Aq�!tV�c6�1R�"M+3����V���Q:��f����ǯ�w'�{n];�2\N\qb�օ��`��Yօ|�Y���aO+/��K-��^�M�_.q�92 ���a���S���+AG��i����
��kݗ�����~w�İ�8����z��c�K2�	=�{�3�l��&�*'(w.�B��Τ'|�;l���.>���T�B��M����y����}��wE���t������!���>���p���/n�������8撥�/z��^s]m��ԡ��2p�ӎ�y�#���F�����?7lƮ�y;�(
�M�73�h��l5��$O�3�_��+��*i��ι6�aiKhT����۶�hB^�h�x3��0� 0��r.Z� w�Fw��
҃�}�C�������'#o��WG�\z�e�h/�n����y������k�͇���>���g���{us5Y����<�6�NcM�ۢ�����n����R7�������� 8j�Ə��L6���+��7���3�ugzO�8=�Q5w�}g���)C�����%W�F[����c�B���YY�VF��^�з8}t�ya3�Ny�����4م� �!�2̘6#�������Qc'�� �2~�~���!��ˇ��p)�пr���#�|K�0��͟F�)ٖ���0�-���tC&���+_� ;}.Y�J�<�~�è�=gF�3�3� ������"~�l���OV�_�P�Ns�
���L��s��)���}������i�]�|AHٰ��HӚ`31�sG!�\Fڽ��ڟ�uk;��cRY/�f���Ksh�Da�/������wB��0G��
�c4� �a�m�j $1K�\�)���!L�n	?
�`)#������B��X��GȨ��t(	���0E��-�$��
����]���������d+u"��[��E��%0���"-�a���{�R9�����>Ve:�T� H�PUfCb��y�l�S���FA�A�d^�޽0��7�@�a7�j�E�^Z��O�'ӏ�Q nů߻��	���b�]X}���!��d��	(tC=>�4�Q@/~B�{��ZV��]oS��셍�sF�wܕJ�с�����v]�֕W^��.�g���K�zɥ풋/�x���)��o��)�Ç�dz&�j����cu��d�)BT'�t+;�z�aF{)��ڜ'�<0��I��G� ?3����T�+VJ궔!"�"�7%#�+.�v��@����SP����~E7yI�.����;!�EPF�:3n�O�M<�C_�W6�m�P�x����RVq?�EᔌP�~�e�t./y���)藌��#�#�]�$sf���0���K��������}#i���q��ul�
��~;7�T7�k�OcGY���z_��Y�+��L�0h�L�?l��#�n�n~�#YtH[�lY;$�%C���c�"�)uu����Ki�����wޗ��{��� �g��� �[-�`��>�,�1y��nX��{\�7�M[�/Cp:v���1'Ϸ%;�2�m�_�ȃ���!�qw�ػ:m��������=4��c��6ÏS�M���y/Ho���ܻ�}��e��)O	�{s�16�����I:r���Os����qF�;�0&*9`�'*Y�P��42BC@����(տ��w'q#�w�5&�E�-\tp*JDhywM����y��Vs�N��3Љ�;�������>�^�򗵷����g����=����~�����6k��>wg���
r��`)W�8�LO�P̳���ʠ 0%+�x:��]9��ͺ�ܹ�	;�"D�=����ʣ�@ݥC13S�أ�8X�y'O��Է�"�x�U1�B�mr�-.�J`�����gu�3��Є2)�~Ѐ�h�}[�K'��	��1=t=$JӒ|t!���FpQP�xC�oF��4ĩ�]����a������@���?�a�m�7���+|�y��<�^�R�{Kc�Fq��ĭ�#L���K/hy�.����i���p�P�{Q����w{(��2�[��W�X�g�:=�"�3�:�3�_����^�yq@�G��cm��#}������y���)|-������d_�w�q����5����?�s�5CP��n

��-���5�u��R�w��i��k����@�x�=�cF�;�7�ל'�W�:�����N�6��n���Ր[�0������u��vxV���'$��p}�!�M47ǐ��	Þx��M~�K^�ܑ�CV5�e����&�g�Q�G�	\��p<�fPzW��S����3��?��b������w�n��r���\m|�K��K�e/{e��A���i�m �`�(��(0c�?���ۑґ��/}�˳C���ko?�w��;ҳ�����g�o��o���v֙g�N�g�1j�i��mm��Ia��?-���S�^;!p������Si7�/�N�1t���8$��"��j����jH�m�SN)ZJmtCa��,�����?=Z̾t��v�I'���N��m`4��>�dr�fP��n�����z�]�C��f̸b�%a-w�Țl�a�[S¨p�|<H��ࡼ�y)��ǀ�A]�x�D��������q�e7R�\�{�ن�^z�䥼�歸�钶xP�Uy������F�@�&���*ˤ�ݛ�σ�F��<n�\u|,(|Ե��.���7x��*��?w=���[ؓ�kV0,�8h���n������W�,���Y�� �Y~�i������W�@=�P�U}�7e���+�Yo�POa�kϏQ�+�%p��%�\|r*P|g�}V@}�hP�Խ+��=��K�Ⱦ�e�x�i4?a��G�W]}U���k��J&V:U�(u^}�!;�:��4�ƛJ���f�_�OC�K�.kGqd���4��22t|�q+��jF��:��mvHv�#��|�V��:!��-�@2��C�`�s�qN;��3ۋ^��v���泳�9'�J�H2�A�XY��S��4u�����;�x�EV�G�|��ɏzVx���)���3i	��ղ&;��Y�`���1r�;��c�x�=���]�������`H[U�*S����oB��!�}#-�FҊtyf�Z%�l����=Ӱ�1Ǥq�&���0bƌC���������RD��Y�r�l�(,ls��L��7wA�Zx���p��B8bԸ"0D��aE6��kpJ��d��x)��J�;�U�a���a_ϣ�B�0�n�EJ���u$K�;����I�����W�@nu��?��y��O��O䮴oy�[���o}kNĨ�YR��<����oI�Q�H}w��m�/����g�3x�[���7���{8�N��
���UY�@�ʣru_x����̋!� O�	s�R`�� �����=�4�Ty�aY�Q�{F���G�� <=^�:�<�)����z^0���ǂ�����t����<��p���h���z��Ӥ�2��)�ޠ�t���3T(�iwq�3t�ؘi 0lJ	��ܮ����/�Un�UH�ѽ6:T���C���lW����&+��a����S����1�?^�p��YvmH�\�Q�A�g��?[4�ʿ��26��wް5��>��,CH��9��㢃�(��=��3\���1���MN��bL����{���e���\�s/�ܸ.��?����&g�X&�;��W�T��������+�����V�o�ߍ���� *�������Y�,Kw��gk�U�ÀK>@S��2��C���щ�"~�O50O���b�8��+����C! j��r�ܭ4�1!I�
Kc�C�wa�#Q�=l�a9
<���`�3+a�$�|�����2�A]}�邞<~r6c~��F�{x��^�~�M?�{����|5�&ԩ�&����Q���ᄰ#xv{_"c�dYւ�!E�y%�.5�3����;ʘ���/`P���~W|(�0��@�3:�J���v��������dü뷶BkhG��q�F7���ǁ �V(�[YF?{<u}"x�_�[��P�	F�uo��|���o�E���R$o��N���,]zh�=�]1$���U�G���T~ޣ�w����+?��!T�}/�PN�_
�J}y8z��<��.�g4�
��O�6���1#-+��eo-�����D~����*�:�}��m��P�ĕ�g���C^�&�+��ɤ���4�x����0�9I���ip�{G�ʃ��56I�>��'[�t�-,�������c[�-�w�Y^�������<�Xr�?]OS�L�2�=�Ѓ9Dk��H��g}���e˗��A�FV,&p�q�jΩ�1}Z[�,\`��!m�L�����q���ͩqf\�=�j(ħQ00�+�$O�o2��D5$�����F*3D�w`X�z6���95�ںk�g��sj^��������>������6k�9?��	��t�#0V���xfG]���"����P ����?���o d����3�8�s]r�%9!sO���Cջʱ/O� �=�1�^P�3��F�<��+�o����[m[��gމ_�R0�7w��h(\?Z0Lg_q+��Pu,�[9F�y4���U�z�?�+�G�?V�OF���޾>������sj�;�����=�}��>�ʤ�FAM�<��hO���~w�6uZ��!���?�C4�G�}Aկ�C�+:D�hi���!}W��#BA�\�B��*/�,��>��]}S�9B��@ZϕҮ� �F��=π{2_Ү��r���a+��7��T>��fX���*~�Wq|�;~\�M�����,|�0����ݠ��O�<�����|{�k^���Gͯ�ʯ�!�r�a]�\��;�o��/�ė���M���;a܄쫯��͜9�]q�������������?��[��;m�䩹��}���c���w85}�/�#����b%멧���>�6�s�{Z���w2>"�0�����6Vb#����y0^�W�RG�ɳ��Is��r��M�o�=�]��<O"��#�G�'2ϸU��ye,�����63���:F�^�j%�����HxJ�5_8Zq�t�+/�����U0?�΢��M&�g�u ���~{�]x��ҫ�\�K��V��eyG���0���SL\u�M�1�2��J籠�Y�Ɇ��?Vx"��}���}�eH+��r4���e��#C�K�;n�۬K���.��U�!�3��3�K���qW��xͳ�[P����%m�t�˻�τ*�|�E���AZUf2>W_��e�{��:��.����:����|���7,�x`t9
<�P��w�WYяgʩ�UgCo}+�����[����ۍDD�s].up_m3�!?�!=�/)!r�tɛae>�e��d�<Vi�6�O?�m癩<�)�G�&~�$r�'���}g���;�D( �W�ȼC0<1�������3l������J �B1`]+/Ww� �Z0,�wB<OWZ &��$*��q�9l���Xl&9���x���M��o��\�����\�������k��k����;����;��;�������~��?Ov���?���O�$���jULi8����}~[�`a����S��lW�-���
�(ߍ�7�m=w_B�p�B��~�*��iW�`�}�S��	���Z�O�V�}���?�rTه�ɀG+�0�'3�����ݔ����贋f�V�x2r���$\F��~g�Q���GÐ�G���ʱ����I<Zz�J��~�]=�'gK�V(�::�a��s�Vy���w��PyW�0L�u�����7��r�E��~WY�h�x�sIZ�0�?�V����n�\���3��Y^,��*�!�Ɨ�C��~�1�)���W}�EU�z窜E�fu�yolW��>E�eZ]�I���e�T͹Z0�H�7���&{���)���O2d%Џ��!V�+�{W�1M6�;$�匋�#��)O��X�G("��4 E����0�<���j��Kږ�[���`��%��y Psbl�� 6��Z{��ߟ���S��w�ޡt�=G��{��O|"w�4�d��-�c��,� qO1V�yå#֮��u"���[���G�ޞW���B�~�A������ޓ�fգ��d�s_0,�0�/�[0Lg_�W`4��|{�*�h��lI��	��o�79�yDd�]��k���*�ѡ�6:mP���ǣ�0�a����{{{7�~�%ˇ0�����:��C�gU�
�A�a\���@��i˦�L�=���=�Hc�v:�jv�NHW~����!�yJ���<�Q#-:ǊZ��sU�J�$c�q䪐��N��6��Կ{����r���a.{�<�3WC�Lx��
���}�)��j���܊H\��  �Bv�0�A��e�$��`b�9#����!AhĚ=��-x,"�Ia�Q� �|���2�b�E����Q~���_� �T�����uk�a5x1�������;i���TلFV�t��c ����1W�y#�m��yWa����0�a ��0�-��g��D��~?�e��}���y�����-^������Z�{���o_a_��w�dBPl�W>p�7+�ꉎ@��}���<!�+�|��xgtx,_����8�m(p_�at^`g�nB�6(�6��;d�+�?d5��4ҍ������9�>����;�ߟ�	C��o��o�;e�H���@w�	�9(�QS:���/m��n4���Ȁ)�%N���*�U���X�M'v#�����m���F����Л���H�����ި��0)Fu-L?E�2/����4�{�]:ǾuG�zWnJ��0m�M.ڬ�;��j������4P�o�s.����	1&�P7u��;s�71gя�`i���<�LP��;ށ�a=�g�����g
�?��7�h��?��ݔ������O>�O�}��������Q>�Q<0L���{�;��� �$�2f��C�z�<V�UY����B����?Y�����˓��t���!Գ���U����PP8v�B��#K]��#���7�׽�u9����Nm�zիrE�}�N=��<2�T
�B�,�uOO�9m�gʒgF��mL�t� ���H�� S��O��0�;5w^��?CCwC�>_[۶�a�D���4eܜ��P���sc��;��5������,��_���"=%p@���PVB�0!��Wi�5�V//C)|�7C<F����۸��kc�8KY��W�7,ִZ#�ǃWVfN���:HzA#�Ţ!��WyZB�^�7Ue�N[I���n�5��[u�'�k�ou�V� 6��őn�-�����P�=Y�^ðG��{	����y�uz"��׷O$���@F���^�%~V�x��4���|[�]���G����';��P�
�C|<���d��Lݰqc[��}ӛ�;�����w�-�����W�W�O��O�#iՒ�{��{�w��������.��*yɳ�YY���0�7�uc7_�ܳ���C����mj81ӕ��
x��f�}��ҭ�Q�҃���߅�'�δ�ӻcT x�(K�M��Me}E}O��K�ψr˕m���	f�E��4zx���5��u�<J�}Y��	9�jН#�!���dL��3��yf<S�jDJ�x��IѨ#� ը�F�i��	S�M�c�� 5y>��C�/LƐ��u<����3=S���U��{Vi)��]��  ��IDAT�Y�f�� ��첋��|�P嫲a�ף��_�����[���w[����뽯�x��W�z>���x�x�y�a���[<�F�Aջ�+���#~��x��
*-���" ��컁�oP��FC�Ox,x<q�0?��_{�F��{��ã�m�x�[~�0��a~��{����Nh�x���K^���[�
T�
��<�sޤ}��9fgcs(�y�W�C���u�����2�a�t����6;tJ�Ay_8���lx�7om�&Om�g�Cer��|��"��}wF(�W� �����|���H`9�D�t#t}�|�G.:�6�hH�+�#<1�]��ReY��I0 �":g���3,�D���"8dEJk��mmҔIm�Ծ�"�S�N����/�嵐q�!����o ^i`�ȸazkƄ@c����*7�<C�!?eq��x#�0��p�w��7�F��`U(
��v����;�2l�o)���G�!���q�aawoi�~V�����z ���W�8�K0,ۿ7<U�]����^����{�`o��͹�+��{4ƭ��O�i��:��*��ַ�])�v�= ����a�����]��HF��z/>YJ�0b�i��W�27A��� >9Mf��(�H��Y�.w2�ַ��V�z �8������4�m`�wVO� �{�Ƒ)�e���0:6��ؾ�\z��Q�L8#�|NGQL
cG^�ȸ�r(HKي�#�����3ۜ9}�1]e��Kt��M�k�䉁��Yd:o��i��4ħ;�����.������a��0�0Qa��&ŚP�_��Z����ba9K�;��5�[�yA��;BȎ����g�^�	ꙫS�sX�H?�7�4��=0�UV���r��*�{�;C��oߝ�o"��vq4>kKpiE�	Vu�G'��Ҥb��%?��%~����3F?�{o�
F����{���v����S���g@��0�	�u���~(��:a���_W�{Û8�����-��* �N�g����ޡ�'ݽ'��o;���J���W��(b��t�yZ~��~,q����N�ݒm�aT+S?��O�j��}�s��l��S���_>�����*VCA�O�-{�Q�
��sc�MHz�/��7dB(��rx/]��.��]���v0�����	'ߎ9��v��Em���m顋s����9�_Ͽ3�M�Wt`6ze��Im�����_���ձc�'���`���HB��Ll;x�ש�!�����	��$�֮�&؂�R�4��!���;c(�͊4���#��ev��|c/ʝ�'��M4�PҘ�\o�2D���G&�!n��Fz��W�^0v;�m�T�N�u�[yl'Ұ!�Ƥ2;2���c�{�?�c����3#�>����/�0�NY�ag�E��U��\u���~���/�-�h�}A=�|��P�W�����J�ȫ�b4]�o�l������AY��*�ЏIX�.���):#�9ohu���������0����U�*����j�[����B��@����F�W��N�8�6��lo0��?�?q��ATOm�7��|����eiਇɼ�]w}�2�я~4�1j[Ƌ� p@��ر#�{��G7:}6����[-���=�}����v闿����3&�~�w>�}���O�s)��9��SC�8��a�̉��c<��qǯh�qD��'�x�lhZ��(������6s�����V*&H�z�C:'���+��t�`R�s�x�rd���N�����g%p>̙5��'��;>vb��ɰ&��N�1F4Zyc �®<pMc�0�D,O�P��Qd���h��;��
b@ �_Ʒғ� 4���r�[��(����2Ap�h��>lnd'�bl�a���xƌ^����9͠wd��>�sLz�T��>������Q(U~y{VDS����{iU�*�a�na��c�7,�0�}���R�'
�i���Z��ν�w��}D����_�(|<��ȧ�;�;�������ݔ廁��d��P�䳕MN 7?$�b	�����}�ӟ������a��:K쮻�ʭ8�q�:n����P�w���[�m>��d�&LL]Ǜ����C�F�^�<5��3�h�z�����N	�{I�YmѢЧ3��14�M�21t�A�_^����ׇ�9�͛g��� E�˃Ȥ�^,���0��lޒ�?nB�Cf��K�Cg�<nJ:P�G��q�代�'�;G���P�)i���|�0Zɐ�2�/Yc�x>+,?F��~�~����/�#`؆�0��aZ��x�	��^����u���@ �q{94Haת�8E(""��X܈�I��x$F�2VP_W�8�g.�C~��=e�0u�,����e�߮������U7���w�~��0��=�We��7��������[��?w��*�h�۳�(Pu��R��r�= tQ<S��w�G=����*^�VȰ!���}A�Y�����z��|����r_�9��'���w��eF=�8���N�ԤO�u܉7���
���S}SχaUע��<E�u�<�T�����U`ĔgCY�,2�si�1�2Uj��2��v�ѵ���X���፛�jj�4K�oݺ9�{��޻�þz͚�R1��|�7���r����"���7s֌6gޜv̱G���>2�,X0�͚5=OU�'=ti�>�ab5��0R&��1ѸO$���c��YgV�:�<�6w�-�1��u-�����P�^�ˈ��=u0R�ŨeL�
��-��c�6q��l �5�n6�Ο����w���^@���)㈷�Q�~ֳ��q5&� ��1�ۼ�"j�k|��3�L�G:�`w� bCԮ���A����9ܒ������ܑ�\�'��rQ~�_�dg�5kr�g�^sM����G`8�3��L�����<���[P�U&0��|��Ӥ�܈���Mw��x�{O���eغ�m�`�yHރj��g���i	�.��zV�s�V����3a�rmݒV9*=�
��e�!����tG��^�*��:<�[Z{�ہ��u]��Z
��{tWi�z>���2��C���,�`�υ!��*� ͪ���[
wț�o�s���{�����u�ݳ	(PyU�@���w�PyT�=���Ăg@|����^�+����7�A:P�{���'U�����{����&��ˢN{����e�7�_��|�����Ҟ��3�G������̝�s0y�>���{�9�{sÍקd�����)a���([��A����V����6�7aC�zl��M�������j�Ǆ��쏴U�V�vd���ҥ��SdNMT��k\.;���҈Ʃ��<7����� IY6���S�djh�F��Kې��G������+��� k�+`�p�10�I<nI��J�iؗ]qE�ڣ�=�X��z�������ڕW]�������v�e�����ՕW���#�y�}M�᪫"�x��B@�$����Np�X�'��P'���<C�vCfi��A�u�*�w�Ig�n�	�y����v�d8�]� (�Wi
�V��9���{)\�w~��D/�ڊWx��h�0���]�����F ��H��;�̲WZ��+m���Ǽ��&�kN�x�V��09d�:&S�'Ǘ�����0��=�����=�Bς��/t��ii�>���]A=G�#�������J�3��z��+�k?tCG'�ׯ��(�ß��T��g�:�W.e���+��w��O9�ۼ�������%����19�dU) ǆF�ߕ�Rjv�{�:�xm�)�g�,:�xNO����a���z�9�����=�S�7�ƨ��B_��Ӣ�3r`���u[��Vr_߷V�JW�7<�!���ݒ�=tI�[�<��zz;,�^ܕ+WEG����v���ڄ����^7b�uCp���m��C�<6��.�='�Gh����Da� 4�M��l����^F����)qH�����[�	+V�S��
�D'm���d�b�ԋ.�(�A"���^���@s_�@�k���rd�(�4L��ّ���.c����9Ϫ��	���7�;ﾳ�rk�q�}�λ�>�c��y�]�� @�֪���<3�gW^�� e�
ie���:d��q�u���ʡl��+�~Ym��X��u��G��?c���-"]��2
��x�|�G���Sh7�Y��rj���]����9=I��l�DZ3fό�!�6�c���o�X�e�L�I�e����W����Y�ĳ�/�8��ô@�{/߁���A���,�贞�t��G�-�����s��n��D��Oު��@�9ztB�ڳ �Q����~U��/���w�F;�E������؁ܫ�����V}��z7��z&]����(��%OZ؀��&����ߵ��oq��|�x�(��0f~g�����YFٺ���=��x�w����O��k8^���w���,��^��ϛ�F�2�����l �K.��P�u�9\�!��}�1�?�/YrH�8;���.]�+�8@|8Q���i�����F����W��핯|E�4��wޙ�گ�\�D�V�Z<�y����?�zM�{I�����{�.x����7�A��iaܘ�K.jmf��o�����i���AG[��VR�
�i~�L��[�9瞛CY&��w��_Ð�ܖ��M�4�]7b��-�7F��m�}�s��Fjs �7oA�>���@Øh�G׎���p�D���IW%Xx�,׻ޕ҈����s�Ҽ�5�I/���e�P������02l�����ڄ0Fŏ���g�)^��`�*w�6�&a�}�����]�!�sP��L;&W4ժ)�3�0�	e#�����7�̐T12���qH����A'� o��~�f�S�g8�:�o�W̮]���Ņ�bl��~ýo��fM�g�������!! �����0��t�܋Gha��C/�U�-([���
��ȒK��<96�^���}Ȝvи���8���;r>�_y�S� ����{��:((�(�co�V�ޡ�������$�=�wL�z�O��T�fU:��=:���o��oRaY��!h�#Ac����'�[����!.꺷o�4)H��êA�<���s�9{����x&T�+/��;���UO
�EF%^��kXF��dF�&�(�2�S�׷�k��JMi��|�,:�d�D����<�iÇ2��f�T���T�{���B��g��ץ�*��*���􍕩�f�����:�d��0��-y30�\p�W�y�}9����;�G	G�S������x��翰����l;�ē#�UY�w���2�W���SC��t߃>Ԯ���4p����~��N�#7�c�l�l�S��!�SO;3���k�e]5t���8�L�xӑ��{�_:������;ok��_����/�!��.������b��������	���OKO��]�6=ܖ.[����W��5�w�	�y^զ/�t�4O��W C�ryO0B���
�S��<7����6�	���
6_�wܖl�r��uAT&�˛�1��#��i�y�QI$��� �-�A��'�!( -D�����u�X�a���/�|��?'��0�uR<#0�#P�ogJFF��3��w�DF�A�@N� <`f����}m�U�qUW�Q%`ZW��fΜ�f͜��㣂6�����i0"o������[��Ԟ��gF}�̼g����v���p�g�n3fN��fe�U�7X嫫8�{�
��/�̽�[���4d��)�G��+_�c�& W��'� .:���~KO\�i����2� �ax*`_�ˠ�;>C�Ђ�7=��Ԭ߰���|���� ��gP�_7��{�8,��+�'O�� �З������M�Lނ��ٸ
��g�]��k޳�\�Z��qq��G�u/�F�����u�����iP���ɍy��y#||8=��i�]}�U���:m���N�!�GrO����e�#�j����v����[�#�8~��*âE��P�_Kȫ{��Ѳ �mɒC��c�5�^�n	Y4u�8��>�M�|����y�Sԓ|!3�Gu�.��/O����oe��蔵�eu�-y�9q�I'�s�yN�^zy/����vk�A[���w� o�I3f�ζ�>��o�%⬍o��Ǿ#1zG?�BxglѝU6r@�����a(&�Q��ӈ[eݕ�r�8��,�����qz^�e8lٲ���YC�-�462��,5�u[��ࠑy�=y����@�ߧFc"Lʠ̪����h�P2�����q��I�Gud�d��tH��x�iE�]��pBț�j�����ltʇ�ð�#9��i��rˍa ���pR'v�Ȱ`p x�M@���|��`�?1����������+7+����;�]�wƱ�����/L� ]��#�j�������`��c��7�S;	��e�f��~��J��|��x4#�<�:�?����=d�>p��曢�!�{j�1�;��6o�65zcڎ�iú��������ܤ���	���/�{��`ȇ��D|���&�Y��щ<��v1?�+L�|hͽ�9�ﴟx�2�C0y���)>��p�oa�U�̵���ݛ�`���xÁ�ʣ(�r|�y��OU=
RAT������\� �7h�Ѕ92�^sm�{����t�F'��"��6�N�a��^���L�\�V�u�w%W���%~��C	�h�o�Ы����)��7Mvz�N��4�W�������<ז�J?�gq�l�E.���4�\�����6��<�u�ֶy��1z�k׭	ŷ)��N�B���2�y{�c��EW!���0>���	�6�w8�,��C<�LZ�G�x/�"�oR*�CA�G͢�;�O�N�E߾��2�����w��d#��1�v���ˣ�m�s/�(����r�w�F��+Nl��qz���o_|qt��2��V�Z�G��͊N߲��Rg|�_�������R���	Vi��7�6���{�]���A#�'OL�x�]w�s��C�ׄ��A#˓FW��`�җΏt�Yr|j�����vs�"o(�1�4yB·�4|�l���,�4�95u��4�ƧT$�h���F��HJuƌi�Kٖ���a	O�!�C�>�i���`2�fCb��)1*�D�0`.��+���B(���:}8��b����+'ÄG���aT(W�/"<c�ꭈ� �veaA�	�5qUo��!��ܫÊ�������a~�򹎆""�ܫ���w�,������/��G����l��#�ʄi崩OCeu0��s�C�UO�)l
�k�a�p��v��u��-Z0�ٶ`˦m���Ś����5k�ezi�� #�Gh��k�n_rq�3���/w�2˫�M�f��Ûd�$%䝺�<��L;jwsv��+����ǘ��]x��e��'�]��]i��zr� O�M�(FA�R$�s�x���v�0���F����� J�Z�'!]��t��r>�kt�{��G��A�����O���(dӐ��/�AK�p ��?��,��Hw4��lH�ה�^���4\����v�IY�,�;��{'�K�Y^���o�+e��c� C׌w^&^�P��\]�ɰ�tՇ�:���s%&Y��pE$:�w��~̓aX�O>�q���D�2=�[6��&����i������jۢ:s�̶h�ܶp�ܨW\.h���vP4��W=�*�gU����ݓ��z;�`et�V��]���k�j�E�.�tI�����@]y���e!�u
����_�Z�C�=Swm �<�b
���V:K0M�3W򅬄+kC�5���qMȬ믿��v�Q�uAE�h��sld��SO�=hn����E��pyd�-�F�,��)���a�+.�,��Ui�08��#a�؜���h��F[m�����j�ԝ�i`#����q�0�1�FB��ў�S�F��	c'�Q��}�_
��p[~��6e�u��� ��̍�0.d��m�=���vǌ1�?5��̩�-���)=�J�_q啉`������`@hL���tp������?~EN���[ڶ�;Ӣ��y}C�bY�'��"��!BysAkp��=�Do#�N�a��ӵI�yn���o�����H��O}�����y*L��n`�:Ƶ� Tԍ�U�^ވU<A�xkx�X���	�cN�͠!�=��%X�³�����������'.�u���Q�������<�Q��K_����׽��8�����y-d �;n�������Sb����V�m&�H��H{L���M�8�M�:=�&RV�C�0��c�XI#�ߞ����p�+�����i��������r�������?g��[��@_�rPC�����I;MfOA���nq�������Ғ�?��?�J6t�Y����kAݏ�3�j�'
���㻅!��N��{��}� �J��-�,�8��ț����w4f� �����ͧ����Q&������G>�42:���h\��3��}h��/yi�h\�0H(Ӓ���L�A��t8�n��=���=2�}K�X�B�R�V���/�r�x��L'M�ce+�R�g�qz{ֳ��N:���@�}s2���y u�Lvv7/���iㆶq�Z�C��8z�ɓ���h<('��l�B�[I�+}BYM���@�a�uE��i���z�+�/�<�5sV�������� ��C��T�����3�+` �C�hm��ą<��5�����C���}�t��#�2&�~!qO�����z�∯N���	�&�]�O�.tئ0j��E����m�ك㍛��T.�{P���v�yцp��7����q��0�f����<:������[��^�¨����k�i?�s��V�����������>��϶��v湄;w�L�6��v���կ��6a��v�Ƕc�=!�����'.k���"�Hz��)3��&,4b��uB��-=ޑ�ʪ���{�{���˗��,��htƑ������C�eH�`\�N��z1+V�� ��m1<�'�OC ��$�F���#�l8E�x0>aB���5��x��zK�(��4���n㧿	�Jp����������1��ĭv��&R�w�uD/�;Cl���pFt�9�}��Ƕc�;6�2���o��}���k�k�F]�
as�U�5!0/������m3~c����o�<�nwE���{��q��[s���X"�^Ř��� ��Q���#�82ǯ�	xt�`����g�ćWtS締7x+���'z�5:�,�o�	߶N�3JB|cɮ��Z�H|���0Bw�w�a��ڭ`x_��gO<Ѵ���O-�������\�J�;;�S���M�D<^6����&���o|�0B;`t��*����`�?(s���@7�w�v|(>��{R����B��������r�+�04��/Yc��I�z�h_g��DY����#��W��SN�4�24:�g%}�C�,��F�H_�Ɠ� �G��y����
�~_z����{cV�߇G���0P�8e��'��fβ}��T����ad~�m�!Kr5�9�<#�0JG����k֬M�ν�QUG2L���jW��¡��ȓk�w;��ڀ���S��XrH)��Gd�|�ژ���\KO��£�ƴ#�B��A�j����s���B6������dlb�2yf����ߨ;�󝴫���s*��,�X�Ǯ(k�;vW���vđ�=̈���/�A۰�H�Aid��ofY�k8kٲCڒC�dgw~�k������ɗ{�bԔ�A0� �IC�QâŜ��F5�D)i�A�N�69���ā��˖3mL)B�掼��^���H"e�r�JEh�V6������$�[o�9�5�!M�� <��7� RvL|O2l��X�(H<ĭ߂|);�c��� � �'��x�ឍ�]{)8oJ�}�AԻ����
���9~���!<�����0c`�<��9���ĸ!�����s�/n~�d2J�kS�Y����g�����������-���M6�s�i0؎�!X7���h��9i¤F�E��O�p}�.�0Ο;/7�"�X�����ӽ�ĕz�|�-x��ZЃU'4�?���hDmօ�#)`��g�9�HG��� �O���@9�Kz@};:<<��{���([A���۳G�F���!<�oP��Ӯ<��������_�g�p��U�ՌhO=q�c>�:2t�ʨ��*��|cr�t�=�I0��E��1NM���?�&>zD��Ԕ���:ÆgX��AW���}������-)~�Ӟ���<�/t8+e�4t��W8&�2^L����3Y�j��p�9}H���m�h�$x��(��|�:�~��=w�����q!��ޔ�S3?J]?��vjGD�0�ǩ����
Ìw.�cu|y��Q��!�vP'C8���V���s���)b�x�S�:�7p����ox�!���gG{U�o�Q��Yh�7d��.�O�!}��n���۴�-?lY��t\��h]r�R�<#a���W��?�:�C�	OX���}N���c۴)3�}֧�k�ڇڄ�/�_�6��1�9;wm�nA;��g�y�礷�>5s#<�F��t�@�hDCkT@``P��a1�#�K�i8�4&����~�_�?~���˿=އ�i�V��3
��5O��خ����^�1F��r��E��z��Ř�`ʥ;��!R�ȸ���8w
���C�?��ַ����-oIx�:�35N���Ӡ�f��6����Q�g�F�$�a(�{םi(v���*�콡��Q�-]��s0��Q�B�sww��.�	$�4��c?Fκ�.���1cƅA�-�0p����uϔ��&�`�˽�Q��+gq0��F3�,�b0�+�0t|ǀ�5�����ԫ�'��aW"z$(	{n\�sQza�:���9�Ȳ��˿l��>��g�� HS�ÑvW��fð/���₊?��oa����}�w���z�P0�u�h��G�4�B�������(�2Z�k���f��Z�ò=V ]�Do>?�@�%�%Y��F!���d�����K�9C�!N������0�JyF1��(./�N%�`��L:5:���S䂼���G��e`��=05�kL,�s�aހM�iѡQn��ɓ��o���n��:x9d�f��oO~6t�xJ��Ð�/ce�CR�|	<[:2��V��3�5�]��3�N�3h;����#�[=E��ê��ꫫ\�-Wf�s8b��oȶ���0���<�#_�\+o��Oۢ��3i�sEI7��z�m&������*���Ke^�]�ܙ{��Ųs�N+���x�]��B6+��g�z�ٱRm�����V:�i#9�a�9V������V�Eb��渚b�@P5��(KrK�P�zE��ͭ�jdi(�`D�
���(�O�a��4/�C �@4`|0�Yg=-�=<6_�`I�8ʤ,�=B��)8?
RT�U]�[�9�г$�F�%-����3�R׋�NϞA����;b�7�S�"�a������Ad,p��Y^e��8��$0	(�q��x7e�\�e,1�V�"�����s|[���~������Y&/o�.Ƶ�̈́Hw|�m�:cx�e��!��Ysf�3�"�}'�]wߕ��˸�����i�|8�����9G�9<�����!e>!�V�����l_�����}o~��| �-��?�GbԼ�г����4�:�/�n{����EsI�#�{�z>�I}F�/�{�����q��T��U}�����ڜ/�2����T���Uny��e �;�����cGc�T@w����%�zħT�Yb��A�=9f�����Ť�ti�-H'DY�����ׯߐ�3��".�4��h$/�W팗��<��3ڳ���v�)�����ގ=����g���<�4 t'/:ز�CC6�JwZ�a���9��h0�V]�ו�AY�)_��ٴis[ƗN�-��e�V�]��������<����ayI��'S����:o�&��E��M!rP�K[~u/�.��x��.=:�sq}�{�+}Ż"�g���(���n�)����p��鉷rբf�i�M���jIS�3�4�d��!y�r�w�na�k鲥Q>4�_;�oCH����'#0ҡx��;�� A�q 
hXD�9dҊ (`�i3!R���ߺ�}�3�
�� �c#-C2������f�k�,M8=hC'$y0� ^��JF��F���Rev-���=&���hCH��s��/��/��9Ƥ,.�ɇ�����=BG+��b�b ���*����Z���ƈ�FU�K�sB�UZ⬶T;�������y/|��[��������=���ͼ9���W����m�u�{}[�|Y��s�)��׾����z[�Ĉ'e�Aѣ����r����)k�q�h��ȸ���ͷ�C���r��z1<,,^0����)]�꯽�K��E���D��x��ߝ�y���T����ʞ�v���	~ijP��Pφ���g�G?�磃r�-T���xp1:��{�n��z=mז��a�@^#�Z�� ��W9��K���S��{�F�PU�t�x2�&��<�£�;���� ʸ�d�>O���~A��gF΍C�6gC�ٳ�6~��^��J�W�D4����{�������.���e�_V
�rO&�r԰��e�`^_���ɾ���8�k����Pݹ�|f�s����0�<�vƙOk�x��g����A{�k_�Eg"�"҃Z�޾��Ю������Pl
Y��WVߓQ�S�S?q�ߐ.A=Ƿ����0~��L�]yw��@�S��!�\���{�/qH�Ʈ��gp)��;�?Z��;�D�BÏw�x�{�����'}�k����[�����h��i��k|�}[��Mʹ6�ƇC�G����ՠ���зt$0���+�q���Cޛ4>#h��f�<��{���1�al����w��Ĩј���һe�hp�� �9��� c�:6&�s͝5��
���7��K�X�z�g�J�G�A����_����g��==#/a�0�H-%�p�AdƱ���f}bp���|4x�{骗:p���ho~�s�"��p2g���ۻ��])�� r��ka���@�Fս��gHX����ab�_�2���bj���a8�!z���Uo|��A���'��^�N<~E���!y~n�v�Q[�`~[q�	9l��B�k��\�/?���;4R����O�1th�|L𣤀!$� ~�@���X�	�C#�x&���:�>����>�~�w~��rf�I������6������9���;���(.u?�=
<+��x�����d��Ew�v=�Cx�4��!��[Ƌ`�@#�_�Wܺ���K�����C�AyS�9*j�Aw��rLW|��7U&�����ʡpc������JK�pfr0e�Wѫa�N�=���P��|�_H��?����!��#@0��I'}y��: �D�d2��o%��W:ӦvoC�
Q] �Ƈ<ݙ�����LCkٲ�"ή0
�����ݾr�W�ҥ��G���sfg���i��;vF��L�����M�2�Y�MK�U�+ìYs����Gg�!b���e�Ԭ�g�l���zҁg���|�������o��o���?�Gv8���w�����ڟ�韦��G�G�������::<:A�
o���K�����)|�]������/�1���NV4]�NoT$~�"�^����P<ﺣ�v�7��P��m�~�ɋ(�F��H�.�ư+gC�Y�b��c�,9���:�r>հwm�A�O
� �i��ϹO�(�����"��Y4��u6����C"�a�l�����������@t�����۷����g�5�Z��1iR?�C���X�\p���ն1撷�NbW>�&3��)����œ6b���ܙ_��_��3��R���#=*�]6ed̛?/�L\Fմ�ӒP�6�'�F����eo O�2T��2)�yI���ߩ�'v��=�e�l	���k_�Z��`��X�q�&�ݒ���1+���[on+W�ۦ͘���e���!(�1����ч�6��	`�Ԕϒ�H(��P�&�@�(7ώ:{�N�K��!�
w��q`\��L��Vδ����_��䮨%B�T���J����h����^�a=�~4�����jK�/x���k��v��R���#�9ު��xq_ ^�ld���*S�(�ߠ�Sv������Qu�3�+A�}��K�f�
�>|���E�p0�JV#R<�)ϣ����W�}�{�[� ��{ ��mW���*98%ʪ͔_0���)Jq����A��0,��
'F�n���Iڦ����W�0_�ot`��	ѡa���L��(3<ohc��%��:B�X�?�&�rX/�:(��s��J	-���L�^ ^x^�&�}��a�QC9�%���b�;s��u�9�����a<!U��~�A婺x.o���� ���?]�(���#-2��gal�Q82D��w��|��7��h��5�I��1�͜��|Ѫ�Vr֮0PBޡ�.;���(׎���M�d�٥Sm��n�❲���п��W�lxJrS�l�� -�h��}S8�T]17��pѸ>Iv�������ri�F����X��ͯ焸/�f;��/7{��1��?B���WH�T�<�.�.4Âq���0��G�w��E��7�1��`p��|/.!a������0��������孹*�Rⷼ�-�����K^����'�-�e�G��=<c8$��1�:*���m�v�����-��pA�zP��rI�u�Q�T�� ����d\���H#ұ	�?��M#i���i�= �M81[�bz hE�o�6�>�iS�z{�$m

=�u�@/W�轪?aK��	�#�_�1���H�!��J��ph����5ږA*�~��y^���=l��(P����_��Y�Z��	|i���G+�>��֎�c4��o��t*-qR�����~,�8W����C�|կ�`t��u�_؝�H�ݴ)E�d��uC02(�~ pߑ}L�x�U�gni�QM؇34�3le�@ΠY����s���h��:"�mD��׾������'/y���Y�̏��(s���<cƄ<U��m1���-3gM�d.�9wcCi��q��N^�[t������E#����BQ�l;�{�~��3�^�	~����/�����*W��ʘ�F��߾�t|[x��W�3�Ǝ�S����>t�,H��KGV�5KO	��[�1:y�X�����-~�7ZVw�2^��'/e&�gF�*��h[A�[��x��L�@����d���a�Ĩ��!d#�@�+��P�����a�vwoB��ْs_���\�8yҔ�fA pB���[�2㰘��q��%�̙;�͘9+=�@�*Cp5h/.�E�=E���`"Wv�*g�=iu"0��zBĤ8ixW��Ac�,�J0hh���h3CV?����YO;+w�U�!H�����P'��2��;��&̣�QٔS�շzY� T���0�\;z�7iR1c� �}2V���`��3�!��$!��2LKi�+�.vN �똈�A(�%K��ȃ��,�a}��ʯ��c7`���w�kfN�9��鹪K4��6'� ZT���P�7���
]]=����Z%�ᠽ{�]�xV�Ɇ'����aò�s�\�>�+C~yN��C��P���=s�hG�V��>��3NZ>=߉�~��ԁ�ɼ�w����l{�F~Wy���ޞ�FǑ&��h�ª����:P:��,9ĉ�
�T���Bf��J�Uچ,,'_�a��eԁ��)�\h�˚N���Ϩ��:$�f8t���<<6r�����w�yg���tLl�a���G�<�< ��"T�?��E=6�bʛ<�|���q�ǅI��=sj�m�n�C���	�I/��F�� 
���|�Dx'}��oiIN���5����:��ir+�Dy�Qy��s��h�Gv$��~�<�T�8���?�i�`r7��˝�s��Nǅ	�𨝢���ആ$�>"��#���P���)=�p@��Ѡ�(/U���F0NS��?!J8� �o����5�=�a̸_q�	!LR�ȓC�����2���Hыg�h�ި��4&�
��� H�%�­�+wݻ
@�0�����{��2���0m��@����;�HCY(b�LٮzU�b�!�'��)�E���b�2��SV�����c�����D�!�^��wޞs�n��(��4u�µ!_.͌?'�N�����Č�;�2B 
j�71��	�0���v�C�Dx��rț���^���0-N���n�Ɵ������6��B�Ó�s�G��=æz��G����7�1�4-�,��m��n�E��9�E�_4�h0����@�����y�\��o�ԯ��殴vH5'�7~�7���<�h;��=����4T����o�_�￞�~��~-����1���Vn�96�͊|�K��m��q�.�;�*����}�P��'y:5|�>x��Ei���Co��\T��׿!�
� 1K�U�6�W�)O�9ew�Ѩ�%��2��P)�(����a�+�T��%|Y�;�5�a�A��B@3�Nk3�o 9\4nb����$:S���M�w�זP�3O��ɯ�W&��7s֌<u�e&�-S�L�Z��2��	�o�O��f�z�S���I��P1�p$�ow��wd4B�'�"Cppf�'q�)�i��7ڧL��?z��u�1j�N��&b�Ӯ�D��x��X5�1�ѭ�.B\�X&Ͷ�a�E�Ə|����y�\���\pa��ј�a�Aq��C�3�zSۼ�\�ymm��ǽDǐ����9|z��F�����
��܊�	�T�[�a�r��Y����#�(^�m�:���)`�8@ф%�`>%k�7�rnJ��U�������X���:^g(�SH�CD[����4>�3�	D����8��;/{��m��g2��&�a�v�Uc�Ɔ�e\�����HlֽUƠ�# �bֽ���K�:<c܈���w�&�6	q�2���\���E��_�W��9�����x��.]�.���\�q�g���<*zRKګ^��m���m��-��f�sv�,�M�j��Bƌríy>#o�a$�F9���􌑨7K8��o��p*�=hN<�d��Cii([J_+L|�.�V &w��K��Q�1A�J��i�!�S�,���/x�w�P�3�U�:�<)]�׼	J��G���g�'�'�N(\'�}����/yz|�~kr=Ϛ!i�_�פ1�����f 6�#4�;��:��a��#��B��d��4S����{t_�J>2Й�gC3��i�����|�7�h�iH�9A�C0o�JsMj{�����U��zg�k��{y(_C�:6މ�<���Bo�hs�w��D�������=�̧�oEy���Z�/�p��v����X�v�����øQ>'�vR��[����Dރ���,�5ySz����s���W�~W}Ɏs�=7=��Q���{�Q���E����e�"������J��ZN�1�Xa*@����1���<�&��ۨ�Ay�Р�mg�����vlS�>ʱj��{�I#���5P|��0'�x�"�1��o*d��U�{W�ܭ�nH��ɓ�;�6� :@ſ11:�������vK$��H\ŲJO�c�P�(�iPJ�1�l�Y>K��/�ƕ�3�]B@\sD��	��b��G&��C\�I\�(�*k1�@�Ȭpe����^���qςLk�{�TFJ��sa*IK*-�̞8�2z����7i�Ѕ�z�%�.���+�%��KP�a������zk�P7���qǝ�D����>I� 3|ģ��m\������9��c��p0�on����^X��\�=Ӌ�o���MlɸB��]�\:6�bP2ƴ��u�~���D�jA�/����ojs���#���i�+��5Wx���?���O~2' @9�o��+"��£vfx�D�ѝ�ҫ+zUoy��sP�"<��d�;:�����((�6�N��\��+�oh �
h���"r@<8�-J�w<��f��x���s�2�9�C��1^њ��\PL��z�!�Fu_{��!~�h ^�A��|1>l�"�4Vx�>���w�I��>d�::vWF)^��g�����YB��20PeDW�����ǜ�|�S�xð�8�Y�0����Cfu`A��5ksb=��͂#(e��o��v�UW�cږ���k���\���)��GI��d^ӂ��<��]r٥)�����=��n���6)��x�,��oH:Rf��6F�G}-C���eR6��]u��:J�L�5�~�CJ]&}�m��Ða�;���M��p���y5�Na�)#ݳiK�۶D{m�a;gAm߱%�W��85ݤ�-[�l�;W�v�̣�e���aEG-�c���|?�ǷҐ�����ږM���x^�+s����Qy-��9sz[�lI�6D�h��6wނHK�1p�l�S��O S�"*�
��b�"D�A1�F��7�%�$"l�%@,��p2pM(K��d�������ҥ3�-}�"¯�0�{q(v��G��Z��C n���4R�q�P3;�oqCXZI�2(�<	t�����������:��|�LC<���W&c����!�I�O���P�F�����
���̆~o����s�6��EQW�!_�2v��G��L��� Oq���y�#tc�#�!�,ɞ-T�	s�|#]�DhD��eՖ�AxW
-^d9�='�$É��P,��/��{i/x*�V�[y�����{��ò�+|�����a�j_�9#�k/ϋ��	�f�v���������]�zW�XÓ�A<7�vZ�c������vU��n�T<���������Eɔ�T/2̀*�0,����bug�
�'�yEϋN����s��7��?)Mx���cU� 495x^�B{��z��3����P�E�߽��o�YB�ʭ^w�~G���+�-7ݴ��n������[��/���:<���S����&���B�ᅱ��t��n�Cz��/?eW^���ft������W��1��l��|ƈ�e��!�x^�hc�-Z�cF���b������qP��ٳ��Y�1coŉǵ#�:��[0���v��Ok'�t|[t��v��E���OlG{x�6kJ�>wZ[�h~���	�C��0@i+�;����o/}�S����;2�m����wZ�h|��Wu�y���;�~��jڭ���\�nm��S	�S�� JǸ�[�^2R0�cd�}�Q��~\<�H�ғ��T�6@�GE(��|��j7I{''5��Xn�!(�Е���7I�����0K/�B�go9y�^x��Y���[�Rַ������g��p�i��^>z:��r�!��*C����϶�==��g�B8b>φ�#< A@�8��BR/��[n�5Wgpm8�	+i���j���� �u��p��#z~��-�6�TQ{y����F�`xe���ŒX�~��7\x������,iL�z*/��Y����Yy)a�wc����)#�w�D���&i6Ҭg n1��ɔ�����ɄJ<Ѵ}_���MB�탮�
��6���}r�6p%�����sbi2��l��g�2�]�5,��P�.���ڔ�E)ZqTZ��e��ylzܾOOM������U.�tKASf9<�F���1Z�E~�o�'�'����(%�|s߽���E�p�))(o������"y���9l@&+ϛ;/��;[\w������|i��wi�;�=���1 �7�B���Ia� :���1޶�ʦ��f�:8�s�W��%2���f�Y�[P�|�n��p�6Q~|N�� ʸ=��)ad���@��de��x^z�ӫ>6�ln`�����WF�M���	x�!E��rOO0�l�1o��0Z�#�>2�f;*�q�!�1�"��9m�a���%����o�|�3۲�K�����0�C��}v�9�SN:�s����O�z|_;��Sr��w��G֎_q|8��ٳ�7���ݿ���C�ׇ��|8h\�/�9k��0��_-�Y�0�e������
8��O�&vV�!.�\�˵l̏B"@<��.��,#��1��0�� �@�V��
1r;"���(�/[��R����X�(@D��[rO�z����@\�_�[�TZC"6T2p�&��ž?�3?���~rѓV&�Hi�p� �~��@�*�Iw� ?��#␷0̻��8�N\�
i5�DA�J��e/K&.���뵛%����kS�Ս7��n��Ƭ��คF�1�IO��L����8��ç0���ggZ�V����W����r���*���T���h����=y���Y)����l�="��g��K�c��E	yx�b���.B��ŀ�;n��t���g~kC0l���={� �����
�ڂG��a!P���F������g�0��{�U��t�m����3;�����M��KK��^��p�����>�c4�]mU��p [�F�vmԈ�^諆�<;:�4��������;�^�X-�cx }��1ᐋ���1�(��PĀ1��e+H�X�CW�YC%��~U~�>zf��O�K.� ���R&߮
���Q#>�	�-�<��0�c뷼�]Q.���7�����M:O8��P��CN��#�v�w�i�d�8�b��?.�����SgT�uh�Q����~Q�*�������1F˗=��EG��-y���a<�1t��L�OC�7�6�>�G�hN�N.=D0"��;�ԓ��ώ租�V�������O:1�EG��s�9Mi�q�ϴ�Y���9�����z��SOn'��rܱG��/le8�������"�vکI3��{�؏ge�5���A�}��#��iaH-���-Y���6'��V[�40��@E,�wE��sģ�� +���_�
E��Ba�H�G�@@g�yf;;~s�bj�����1/��I���-���}˕�;q|�X*�"� (�@��/P'�	��<F���1�I���w���z"ƈ��l�����Ƙ�r�?ƀ<*�Q��y^e�u/_��u)f���I)dD�[�lJ�����4��	��@*��{�D�S�҈�*��,S��*�P���#��F҆���E�)���x��e��Qt�31�Sح�#�e�h?��F����JGqТ@k'F��Δ!Ue��2j>�*�Acڞ�� �v�[�y�7lÂ��@�1:�a��+����V]��&x�^�F�10bL?�U=1p(kW�B�����_mw�}g�����>�ɏ���$�R���WeB�=P���RG�x�t}�k<;O��yGIG٥Y<5�C�]�w���7 �1$<WG�S����D�-*#���:~�	��.�#���r�G�!�槐��i��9Q�N�ҭri/�z�Sr��o��wb?��s�7��δ��e����m�*�r x<'�N;�;�H��C�=/�?����<538��ʫ�J\�g�����Q�#�]�6;3t|�/F��7\�^��x�xS�(e��<<>k�b�/w��Yv�y�Q齫�4e���վ�Nm$���� �0�����,3�3�,f�3x�<H 	#��ERK�+�mfVzo��/΍7o��Y]-UV�͓���O��8q<r��qc:>ꤸ(���I�5������?=�3�Ac��|��@XS�C��z�����(��x�3��!-�����酸H��<.V�N��ݥ	���`��ru$�kҴ���zS@��d�N��Lڗ���	���}�����i���ڗ��6XMu����ֶ\4��DʯL�{��(5+��$ǨC���;*�J�g�������׮�]j(h��½�����b�N[%��j�i����PZ<B�^={��b��"S�-_��j�	��'Od����	"���� T�ÉX 1�<qV�K�1B0#
e�?Ƒ�\��O�����Ic��
�0M1�~�!n<��a�R�@�!4�Yaf�*=$p�b����E���o��K��x���[�U1��?yٺ5��fǐ7;��YS�Q/���P�e����=%���4�R�C�L����� �K�2�M��C�4&()���uMm���Vv�AO����# mQg1v�5�8������| ��{ ?,�?t�?x��`#d�=<��9
3z�嚆��p�b����%"����C>��@�z�N�(,���DϿ��6�N�d��A��,J5�/���?����Λ�e��A���)٭۶z���>�@v��,����ހ��_�7�Mj��\iDҨ12�� L�:$��"{�;����6|F&�ᬩi�l�2[�|x�Q5����͎�u�V��?yZ����)o�\��~�1��@��^MO�).�="���9q���I�uz��q;��߃���J��e��Լ���C�<QN\٢n2�@�	�#L{B7��q�mQޱC�B	�|�܂ghZF�D��I��e�0�p�J��7���'PTJ�K|ԋ��c�����ꠍ��1���+��|����S���U��Ţ�cSv�\:��P����JN�`�-ۜ4����GF�E�L{����a�W[u���S�Dq�R�����Ҷ�NWj���()��b��(5THT,O��`�J�;�Q��T�EÎ=H[��a�$��@#}@ |�ø������PH?1c)�ff�@|���7�@�&N����!\���˩�lo���ų�L���F�=��}.-�C񡷋8�N `�T��x�2; {��A�8顡@  ��pN��\���!D/^LG�# Y�O���y�<S'^O�o�5�O�q����	� x~���}G�0��|��!X�'u�
"�C0�x���1d��S	�K<��|�(��B��/8&.=�	�E�F/U9w��u�M�7����^�����p�Ѱc�	(��Zp%�~;i�)�G�h)��)P��7uPnp��	K���B�9�
?��:�����FW�3pO��C�OD]-���yܢ?\�~]��҃�<O�'�P��%��ШAS���2���+�y��o \�0�M�4,�z�����'�^Q�)/a�?t�"�?z��0tǴx���:�	�_8��&��rDC�h|��G��tx'<x��	�FLN�:iǥD9tį`���첡~�C>�+�GVp@[R����
|��9Ә�!��%G=I��1;y�+5��9�ÓRlX������C�!F��u(5����.�Ҧ$ٓvR�G�Ag��zAQsM�7��a��+�	��2�4F���~Ζ��/���NY�O�2J��$�Ud>�?r�㛝f=z|-j~��_����p�{�q�ƃ�3O?k������^�GN����s�<o�H>~�k�ÒQ��ώ����7z�z�a�	v�q��W�+oz���x�]��S���f��P��U�m	��5��rknb�3J��[Pj���%��9�*Qch�h0�@�wT�M�@���,�!��� �`:�iy�ߤ �S^�q'qF#����`�i����ye�-��D�{@�M+��ի��1�/�$��!�H��a~�~�{���������iЈ��0�Ʃ�|�ٟ��q��O>�&���v e���r��c�#":�Q�!A�>��S����		.��G�z*��F�]Q?�Ɖ�w�%�wM��e��#<~��.~y�F��7q��`�#�y���{����/�S���z[��s�������]`�K��o�!�t��'g���V{��uv�%3z�A`�:Ǥq@�40�3i�g<�'�p7�Ƹ�L�S��Ղ�t��,�<SW��m�����������x���W~��)������:�5�	=N��[4 4��˔	J)�C�0��E���a�q(�y���ӕ_�����~2R qQ)�JCƄ!}vj��o���ӌ����~FB3�o҈z��z� ߠq$F�o��F���.ɂ�ճ�#�(�y o��gذV�/�k<Ҁ���٣8����8Ҧ<��/��|U���6��_��_��<�< ��sp�<f�>���)�*偭��WMm�z�M^.��G�dOc��H�`�:={F���!��/�p���W佷�7щ�!}��5Ϋ�R��^�:���a��tz�I����r��K�ÿ�-@�,?�ٟ�Y���'��=�9���;0,��'�t�G�GE�B��0�Ag�A~"�%��x�m�H"yUh���L��'O��C��p�U���*��Q���I��T[�p]Y�b[�y>w�o	��E��)�F��9��p�)L�pl���Uu��������2p2!9�j��q���.�h_i۶_'��Y~�#P�5)5&J���>�1W j� z�0)���d B� ��� >�"n�og���F �1�Q��a��W���I�3����9:ʄ�7�'qm\��OAEۧ��������@��ρRCc���!@���4�0�O��O{σ|����;ʜO;�C� ��w��gzL�0�O�!�` �<��a������E�C�8DK�8����m҈�Q(K�>q����d�2���w�0����C��߄!O(-�;�x]��!Yl��&��۶m;�a�h�t�"BzrA�2`b�t������=C�\�o�2#�P�&Fp�a"�H7�v� �B�F>�}�0y�����(�Y��m��SV��/��/��w����Ĕzޣ�gL�F|�+H�X'
7��H'uJx��/��/;���y�!�4`~P���>��S~6�{��nWv���)��N��[o�ٮ�b��O�b����%ҏ��? oO�|��~P��oӀ~Cr�������5�$�e?)p��H)��N�цn�{�`j����F�-<�y���+d�ƄE	 ��G�(��mii����PL��9t��sH�Z�/���/}�R�_J<+��A��|�q�>�`Ά�F5�s#&�ާ>�+�<��(r	C���"���esIE�:<-ͮ(@?(f�����|�o�C��|o�[e�9�7����Ṁ��-�;�J�ů����o��N��K �O��2�[�1��i���l0vA�\�@���MH�+!\������)#cЉ��
��ߧ��oڥI'trzB�,�V[):�{�:;�ۤ�~�
�Q�8��A���~��*H���fY���i�zko[a۶�(�4?���5Qj�4�"��$���7_a�ذb�^��h�T:����W͸��&�;�����'�@����P���x����Έb`O幽��$|�O�<~�^ G���p`��#8`@��������/ރ�ip�~ɧ��LJ����QH����݁��a#����{@ؑ?�G�Τ��AZ�aϻ3��9�	���"�X�bfY3�L=&E$)5Lr�3s�4@��S|c��&�L/��/�#S=T#�b�M>��[dU4�aH���L8a`,v� �9��ӚQܘ_g!����Bă�DX1z@C�).A�/��M`�������k��' ��k����v(��9'���|�k���6�/����n�We����K�03�D0h�z�O��)�b1!�9*�K������F����Ç�3����'?�<��:ȿDy����~�#�?I[�v������qd����}Ē��(i4���q�G��{�}2��J�^.|��4��R�+W#�TEc�52h%�A���oڧ��(���(ߑ�v�1�e�5# �:B�Td~�בCt�Pj��N��R�g�����J�G�RLx�����qs?�Mtn�b�<G~�rByC���Mo�<>#ߌ���RN�Ma���*W(���p�	��<9�I���B��P�~�w�뙫(#�:gpɈ���D%,����(g�gtʎ�S�i��}��k[�H���%)3�������}��&�����0��A�= ��6��\O�(�A���}Ѳh���_� K�<��fECȰt֏���D-��Z�����i����%����G�e?���J_tMޤ�=��͛׺L�Z�VJ�.�Z�Qqd���r-&\���h�D�����R ��Q�i�gDL4*TVT6���{(,��W0�����x�NGrg��x��w0�k>��2ʍ0��W��D�?��e^�� YKC�w�N�a��xc8C AD��7��3Y�Ɋy�a�f�4��凐?u�/�<w�[��þH��U��yv�Ns��sg�W�%����C�&�� ���:~�	��I�������Ͽ �{3o�B7v:<�ܳ�����ǜVN�:�F��Ꮮ���G|�y{衇��r��
�!�H!����?�n9X�\���Gv<��팫�x}KH�X :A��2O��F�	��� �\K��!�A�A��Ġ��{��B�;��Wp�;"���G;����ˬՕ���T��{�gD�,pdD놛n����._gB�|��)���;��_�O�/p��w���<b8�:�;�۳55���ј�\A�@��8F\yb��UĽj�*w��"L@����ppg����3�_fuj$�U�%�wYK��_�������N�]���FT>dJ9�(�'h-�nB�!q��R/�� S������0Jx��@�.�N�eh�Ӕ�聸E�	��7K�oJ�x
7z������� >³�	w����j6n����іI)5ࢩ�����������5����v��A;q�������%?�v%Y�<��)+���G ������Ǩ�g������ڧ?�i�gϾ�=|�e#4C�,����6�W�A����	>�	i,A�@�$*У��<��3��ܦ�	�1� �R(��CK�����(+
_H���U|�<�����+g��M�&E�9'9��[�Qx"���%��Xk�֬�F�j�6�_��BI�؉h�ᚌ�@T1R�����o��k�4*0B�5	�KB��&��@j�]a���]����9��P�'���y ����!H~��~�O��Af����O��qqCO�� �<F�XІ�eC��r@�1]�q��C������[>��)34�0	x'O��G� �8�af��p���YUU����ì��܅ec�uB�z�p�L�L�}*uψ�3",�2�G������M)�	���;\�!丨��P�~�C.b'%���]���aaS��ԧ\1DN6�0����1��>��g ���`=)�Y��Ptxǎ��!b��Ҁ��k�� /���z+��@��HR�oz��?�_��{���^|�y����+��� z��
���;��4��@R~��>k��{����yǝ������r�-�ޞ���/�+������>�#0�<bׁG��:z��Eư �����/���pA'��r/�L��^���ɟx��Y ��|���#����)?4��q忩��J%ҪD?�m��m��.��7�M8dnP�o��C��������O蒼�n�^)
5�3��C�B���^��#��A�{6`�JyJ��7�$�#,�fT�E��M�p��0�@�pg�����HR��#����ɺ�Fu�*_��g�x��T�E�N�J9�ݒ�[������H)P��jH�����➵Ύv�h�����贑/ֶ����ap�7n�cĆ��o|����>J�.�TGm@����������������q�+�2�?𑧕b ב����W��E[�q�a�/��",n��Gc¯�5�MA�<#�Qo�E��v+%�I�v����Wo���|2��LM�I!/���ew�y��]��v�ޫ��E�6[$����#5 �5g���"E��1
�b��GN�]A ?����J[��&�N����A�G���?�py��Ǆ��E�+�(;*��Bh�3
�-Z=�e�(?����#%(6�J�'O0D#i��sC���J
�JaP�8��z�q�����[Q�8]�U���SFi�Bgx��d���~�ZL9����]C>�>�%�=��]�1=q�W���j(ϝ=�8$�XPϫ,�bAP3'��k��EA����������+�z�C��gӅ]9�g�����`ф@���P'���<�% ���o>�����eq�w�Gy�����A}RfF����C�e�׋8f���{�]gw�s��|�M6K���>x𰏰UU�؇���}؟��p!G��\0���r�-Y/z�*)��?��@�|S�`��Q�믻�z�z����Σ�ΡwF4���I�3R��?�!�Cǎ�+�7a2�3A��p�T	k�����
#{��7R�W���^�����cdC��H�<�eRt�ʏ4����f�9K��O�����_x��z:���<y\�٣�=l�=��=����S2��SO>��=��3z>�a�|�I���8d��?꣦�I� �)���+B��C��Zd	׬<���2|��1�����������~v���#r������,�W��UyE�=#?Lw�~P&ڒ!u��7�W��� |a#[LSC�18D�a�)�r��� ��@����K7\w�_i@�1�D����4�����I]��ħ�V�����M����!�K� =�x^3��0��{�#��ˤ�K���{�{>�(�m����iM��+���U��`NQZlH_D q B�@
�m?�����0a��@X<�:¸M޹>�����N�wI�r��7-pc ��9��k&T^/��қ�qg7�0��I������A�;i��0y?�	� �:zfza�������u��9��y��3m�Da9w�[
�z���Ѿ��"�����Ks��;5�,�*|FA��Y�u����`X��c��'k!hH�Ճ++��z��S۱}�/tL��u�
JuQ�4�=��0��9w%tH��o|s:q�C��߁[��~	���ɛ�
��&��T���˕	�`m͜?ԗ�>�D;4�G�O��O� >��R4�������������CRhh�~��~ߎJi���}������Z��w;Ӡ�{��~����/���b?��?�k?X�˔��
5dYV�W�rK��o��6)�^^١h�s��<b�!�O���Zx=��8��;�Ζxc�����{�_���Z���lX�
ړjD���4�J�VӅ�1�W���:�dB���C�~Q�'~��W�z�&�~G�bzc���Q$P����B��Z��wF5ֺ�������:k�\f�ڗJ��O��yF!��;5�۷o��n��en4��a�.W`9�E��P#%�Iq��"D���>�ZW��� �E��FQQ<�5#-�c�����}(�< ���ч�/y�;v��p�L	22PO.���#�� ��i��$.�-�+4�\�.(+S��7���i! �@�d�̬���>��i���e��o��M��z�#�Dp�؝��� bԙ+絀E�a4��� �w�\f�>�h��lh���*?���� ���+��ϻ;�5����y�� JS9Lʙ4���ɝo|�|��)���|����(?�F̂Z��xi���bT�F�4������[���D!0�e'�?Oz)��F��"g9�y�v���j)9�/5��! �E��8�+����p�r����z���I�ư)�Ip-C�9p'��)�m x�+y�L* G�!��4�Q���xC  ���|#���䙰|����%-���_�<�?���ȗ#h �����/SC\TlC��1δɉS��w�Z�%��L�*ԣ+S����������_��=��=���m��-V%2U�}�k�hSq�@�š��2��O<�y`�MH�Ũ�b��e��	���L=҉@مv�FP��P����^{|��(��W
�����2ҹi�FW�a4�i���o\��3��K�i��F"�� h���"O�{�a]2�<3�C�D<A����2Ϩ�Om����)u>g'���L���u��r�P�(�[���/J\�a����e�۴i��[�ڶl�l;wnU�a�56�Xg�2[�v��SǂKf/���(ɬ�b4����|@ciZQu�w:W�S��>�Vv��r�<~��EY({1�Q��xǡ��h-�p�_pΙ��^ h�q,C8v#1�C:��e�i�ܤ������C��|�	�i7���%���h2
����4�(W�G>~��`��p�^ ����'�������qfذ�"�3jߥ�Bkפ�ǎ�8Q8�4�c�`є�@�B��4 B�aX{��F�1 LA`���*,�7*f_���X宀�����4y�8�(I�����Pf4j�aJÁ�e��q'��,bd4�|�`p�$s�`��R���O ���q�ȝ|�L�����Pg(�0����b*
AQsgC�,�dk.#Ql��wǜ=�(*��	o)}��Y��Wt�駹\F:�3�@����R�F̷S
��==CS��!C�Qn ��y�rp��<P0���ąp$.�k���=�I����N��<���+6�D���r�D!d]�`#���
ӊ���^W�>)qL'�+��R载|��O�|��i;z���Y�ƃ�_��_�3�<�2#et��lD�84`=�
{��u�Fo��^5*ݒ	�6 ���鶯=������N-�1�����)`=	<m0��i��4����JOꑆn��>-�;Jp9�&��aA��O��Z~�啾��O���J��Q%�X9z��@qf�J�|��wвÇz��m��T:Q�YҠ̄�2����0,�o]�.����0R�p��'9�s��D+�ѹT��:�ᦽv�m7ح��Ѯ�q��޻��]�[�l���7ڦ-Rl��lڼ֕�u�l���u�&)#j�6Y�[-�������:��=oG��՞u"(�t.�=�sW�O�����׫8�}-��QfdW�����E
S5|�8��#G����\+Fkq�=�X&�\����x��X���ŝ��~���xea�b�P�u�!\���8�S�!#�aG��#@l�䒀��#�D��ϟ�N��R�(��*�ݟ1gV�X�k�8���=M?��+6�xu�&C����&.���W�R�`D������8�O B����a��
�yD���ރ��%8�wDQ����h4Q�1D
q0�+�}8QL� ����+_l�:� jL�-�#����h�~�I|rFC~1�A��%������pQB�N�fc��@��I��y�c��Iߊ��NN�5E�[BSiN�p(�����b>Fi�����CeP�_�\�F��.h�r�_�a��K�e-��"ʃBD8��! ��#�)R�Ȏ����#�`��g1~>�ZB�����]]�я~�oF��( �>�����Җ�s�4�0{�#�NY��յ��'M��>������v⨔�矱��xԞ|�{�����c�D�\[]i�e���E;{�;r��������v��Q_G´;�8Ȑ���/��bv�Q�(�,P��pO��~`�4L�h�xg���Nh����7R?��(2�~�nr'dVb���:M��8��~g2?�>� �(\�I���b�L�p�H$����I�`��2bRQ���=y�a��w�|��{j˦M�9b14e�Ѧt���F\A��;G�zph�.t��L���BܵR8PZn�"s���l��s�V۸i��\ŽS-��4/mT�1���$S�5325�V[_e��\��pkni��(�f�*)=(>k�6SӢ�t�f��
Je����wFQ�D��w�?�O��m��O�?�ϴ9�����A8�����4�t:�o2�N��3�f�Y�6:(6�vp�l�j6R��0�[����%�/��ueH���ǎ�E�Η���%~|�4"�ڴ��tYbRj�-�j����4R�T��!2��(JM1 � T�l�" p����I��'���!*�g���z�%����@��
ӹ"M�����aN�D��A6͟7z�4�?���d�?��?�u�A�^)��>��$_��F��,�x#a�`yɒ�?�*>y�����g=,|KA*��`\��R�=�Zkl����,� �hM2�-��a�M�U�pJ%�l��QPz��3���W?:����j}��(��g��(�25f��8�^��1z�,�^�b�� ���7��={Bҡ��g�����ɕ���J�1�l�$�QN�EqݯƟ�Gl��х©pDO����t,�g�
;̶m�fKU��c6��k�z����nU�T&���찕��m�u.�B/������6$����� �/Qo�_�@��82�)Y�buu�w�8��.g�4������ذȞ:D�f����Da*Vj�;
��3�>�
�qC�����G9�g�(-��6���T��@��COy�=GUlo.�yJg*Qo䗑M�P�������T�4�(3t��[�/�)��w�)-���s�. xx��{�N������1¼[��Z�\��'ܲ֍�%���p�-[�9T��+��0=�I����UyRg%���MJ�d�z��R��%��r�a

ـ�a�����M}��͡]�5}56�20=x!M�������#��u���&�s���k%��e����,�|R_WL/�� �E�Y�à�����'��4H�rE8��o�<�]<�i�g.h��Sn?|o��ʤ�z[�Bm�R��w/zR�����D�H@e H8k$Fj�x�\|Mͅ�N�� ���rD%H/���F*�����J@a����Ay h4;�q9,!�ԓOz��Jb��{epgH�������bq�J
q��<c���C�!/ ����]X��4�(��[�ٝD��/H��6KYi���q��Z���5k�|�|�����v����nܫ�Գ���=v��v��f�wrq�j[��KH��$,T+qŞl������2�[�/�g�4�LL�1�]!$YH��A81�RH
�E���`h4�3�=�C��@c��3"6l��Ap�����)e%O,ݵs�/�����D�����>"����_N��ܯC5��i���q�[׵�:���tCW�m�s����u�z[�j�m�W.ZY�:~�m\g[6�����U+}!pS�R�����6���*�� 1��i<G��ꪴ���21�A����pe�?�tV����9�^��1����	�p<;�w*��4�أ��u;�#\C"�OFHb�#4;<�T�:#�v��w�����X�=3����E��L~�E���e°�������Q:+�(x��Q))���nw�y���������G��3�����^5�S�ʁp(Yi�%U�]z��7�����w����ؔ�v,���_��Vږ͛�4o�)&a�f��jk�������j��R>hg���f�@~����e({j�G]q��m�ZHF����;��0�� �w�}.K�'a��� �c:1���ͫ�Yn.�\�� ��?�+�@b|Q&L� 7���a�|�m!�hy��=�;��(F̒DV�Z˲[�n�O{r�eS��qW�ˤ )@ֿ5�(5 D������A����Ї��Vj����'~Bf�_���M����OY�h���*�S6Q^��ي����Rd�q�2�4�l_��JP�����p'/�� �A�ߺu�+��+f�s�ڵ^?���aG�;��ޡ��&5R۶o�{�����{���n��n�e�z����Uֵ��V�Y.�g��^�R��v�Jۺ}�mٕ߱�={w؎�\�Ya�ٲ�V�Rc�B31��Y�E���Bh�h���
�yg��I<N!e�)��`��	���6e�'

g�����I����� �x��ZB�+o(7@��=v�ѳBQ�'��J�P�=��g�pk��n�M4������^M[k���L�`���,�*�[U����U]VK1�TϾJ��C�ʬFv���V_W�Br���ݻ����Gk8�eÆ��+�(`{���Q�)@�6m��z�l�gT��m��0B#�����)WdQ�CN�Ԡ@k�5S��Q����a>���_Rh �U�7���+�ޙ#�
ᇭ�[P�]����QF�|���	���)ِ-F�a{3� ��/L� (��+w�<,_�j7޴���ۧ�IK�ҕ"31ŮE�ʧ�,�o�ilL��5%� w�����b8�������G�x�utza��z��be��Y��{���2�u��9�V��f_�qJ��z)cg���/؃o���N���('Q��ut0i��C�Y�D|�#<tF?��/��?���bC饎�
,|�������?�%�'i@��&k�p#߅r�D����bȻ�Iܐ��/�cd�3��!:���2`a>�E�ȴ���4�(4����]��R�l�D�0��<7�vTCV(5��0�ɂ�+���l�b�0��}Q�+���^?��h����{�����0�Ύ�|��i���ӈch�{�E�z�D�k��]b�>Wl詰�b���\�XR2cC#X�����iw��6۵{��ܵ�6JqY)������4p��g"r�1�m�"%&@pWVq�������e��s�۶�?�i��.5V�~�*��0�#�](��rUZ��О�S�~)	91��c��e�i����b�*$���E�R�05ζR�W)�3v��Q��������B�3�����x�z^�N��~���/�ܶm��s�ݮ,��B�a�;���ۄ�f��օ3�����خ�;l��N+��YspaS��H�9���.����J�P�TQƔ�x\O�»��wG���l]f�Ӎ5u�v��P���
s�Dh�QB�B�(��|�
)X���ݻ|���>�����!On�0�Fݱ^e��hȨ� p�7�u�:�ʧ���$�@�c�ܺ�����?Ń�7�
QuaKn]m�h���G�ԩ�&�RAY����.�y��?�!:��#�����+\Qe�|��V,�2K��E�c����=�o��:}��)�IF)���ј����U$�-G��إE�;��J�-s�ٓ�B����#�Ͱk��C�I�'�E�حZ��5�w�dVSK��S�{2)�;��R�?�
�+�L��؅?��=u�72��&#�sJ�B�B��ڭ�<�������3���b:#��9�J2�C�QOyZXR����,�i30 rC��5_���<ė�!{F8 ��&�<�BF#�9꣈8�;��4���u�$�ğ�-
�FŔ�1��\y ����K%8A�����VRZ^����.���w�+../�CV��~��(�A���I�@�#�����P�K�{�_p�D���;����%�晔��[��6��������ָ��n�m�}��f�����M��z�{�6[��ݖu4I�VS�3�2Ki��P�s|�&�(>����L`�?�I��1�)@h&���Ϛ�*)7�j�:m���v��7�;�u������mk�*f��Rkh�%���y��,<����R"���9*/�%[�Q@�.�
�Љ�������D%P�fd�����J�<֪^�԰v0�^UiM5R���=]��bé�0/��y5uw��4���;=G�A�$�P�t��F9himqE�I8�L��]z���=i&*���a��j5����^�D�2�3D jl8+��>��D�%%�9SGB]����F5Z�j8��?�|Jh��r�*���'J��Y4Lc:1>�44l��-C�,�emJa��QW�suO��'��G">v�pY#n��w p�Ƀ|�?�����ah�A�my���4J��Q�o����[��?���k�@�*N�e _�_Y]�t�0#T]ee��%�lVKy��n��ڳ޶�Zm�+���^y�B�b~?�Z�� ��)).S�?��&��)�T0���g�dK锼@����.�T�[2�wΖQ'��;�ȓ�z�dKfuH8�i-�Hǆ)�[n����]o���w�u._��F��񬼢�Dc��W��cSipVf����Q����Fi��N)�,\��K�q�P	�K6��[mU��Z�i]�VX������i���9�@��߰H�1���|��r�hL���6�!�|�(S�9����2�C=���8N�z��"��P|�i�I�yM�������A*�U�<"�@ �ʈ��	��ܮ�ȏ�˹�c�P\IW
�x��ŀ?�O��Fya0t�����5�D9���tn�.&U	�1JD��z�[O'�r�'=���Z[�j��|�^{��n�������d˻ڬ��D�m�գ�u6�j䧦'Ը X�Ƭ$ՌR�Ο"5�@a(��O",���i+�_� �115"�0��X���{�m�پv����d]o[vlT�:�AB9)�L-q���_jU��ƽ$B��B��/��nF��і��� ���J5�3*KC��߾��ZZlEG��]�^nm��T��;�� U��h�����
ɒ|M��� ON��_�jU�7�N���ډ���s;;kV�u�ܥ��$�@��R�yy%��AT�ZB�{�|������f	��=������CH賲�Vp�)���1��E0W��`G��Xǃ��Ç9��i;t�������FghXxg���s�FعO��O�$�̩�L3��S��	���_�\f̙�ߕ_9�/���h��A: ��i:~,��i3:�@!#���G��MOo��!� M��O�S�z��m�&�Ŵe�Z[�R����h�J�H�#|�}�Q�R}0zk2i���$;~d���f!��	W���*(��T�rP�
r(�`��$���rh�N rO|�8����|�K9m�;������7��p�`�J�7��8�v�di:p�Χ��+3*O�c�7���~d-�2BS����ʊr[��f���F{��ix���o��s��}ƁN�>�i��L�F:yڹ6h���y:E��JNޞtB��������exC�&�+�)?�	�#K��%��(�tT���:��@��*$4h 
M�����!�*
�qd��2��������x��<�S�ŀL>��r�<�E��!���R5�OPH).�`-����ȍȊ3i��_���������Ծ���o{v�����`��2�G\�t�/��L�@M����oBN�;v4��X&|�ɨ��B��c3��FsUW������o����[���::�t�R���`�CLE�Z�z�K[:$T�i7b#�I�Y�k������UKy�o"����J��0pGs�zv,�֎ej�l���~���mۼ��/���p0
�����t� O��D߷�|�O� �Qr�zb:�Q�c�ӑ��R׬aA�:������C���<�3#���/�Q7��4��B�Oe�\�%7ZE����Q�$yO��'�^���@ڥǺ�ݻv�T#94�@4�aQvX��4��I����Zz��' L���ʛ�2�_�#� �S�� ��O�⎒�Ӫcq�XJe��ƙoW�v �(��t��)�Ȗd5����2�}C��۸�n��:�����uk<N��BZke����*� �<fUFbJŃ�J�bROɏR�2�Z�1
���J+����5M�@�)I��ϊ�fjd_#��Q�uFʕ���&c��*f��N��4�|�K�L*OɛY�OM����(mε�喛l��u�q�I������P�2���.�_�d�#����#8�	��/ng􁺠c8�����C2����=����߯�x�}o����풛��45�	�0�N�\]F���Y�:?�:g�)3��@i!~�}��||cO<���V�8�hŉ�S�.<!��+�~�5\�i��X�!\`" dcحrQL��7����� �a��Mso�A����-�g~��imʹ�Ġ��Kؕ���l���������*f�uf"<O�'�/W��z�Q����
��1�V���`����#���5���Y[��N�͍�������f[�E/��6n�l�ZWȿ�2�c'Z�Iu1cK�����S������J$֨li�-Nw���=���a;{�:t�N�>i�#C���u���B��MBcɮ����@@�в�������2�lА����#���]-K�����2b�4�чڅ\�E�iu)�A] s��..h��L��l�_�㪌$���VS[��,�����������/����w��J���g�Y��\4c�p(�E	�J4��;f! \����-�c�@v?�P����a#�8D�n�=3 e���K�$P[;;�Z�km��ٷY
���on�f�Ќz�L�J��)�U�
��L����\FJG����J��GX��Rb&Ǧmld�F���̠�ΰp&32�Ć�0^���~��Qf:�tx�.HQ�R��tBr���3$�Ɩ�ܨA7�G%�fՁc3@�ݯ�;��V)g]�3]QC�+*�20�#��5�4��_�J@��C�<��=��s��R��6%��F�v�z���,X�/q� #���w�uNo�2j��3�M�&ho! ?���iP�J�P�L/tP�(�wL@^� ]ʍ;����g(�|���(��2�d�)\�W�qC��n2� ���&��C9�e�!��F�-�p�ϼ�/�LT��R^�(�1�	 _�`y�����*���E�3K�N}�VB]������o�~���f���;m݆V+gI�z-��f�?z�0q�1J���җ��R�
���F���#N������wXL�Q��7�E�ޛ��7��KlŪV�����v�]�n�\�f#t�B�0�����T.��D��y�P0��ހ�;6���{�X#�k5�����^s���n;w���<y�N�9�B����){m�Q��d(zM��	�.�,�Ey�?Y$�<PFeXO�<ߌ�p�`lFp�k�sQ�}�~��qC��-t�I�	O��U�L���#3��2�XQ��I��nI������g�i@P49[�� ?�� ��:��w1��~�W(��+��>�CW@����/6���(W�y���/�ƂV�?�KD�<�v2��{��ſ(���l��.��6۶c�ҒLFЮ~,��	e���&FQ�0��H�Ҝ����4a#���;l�O���^:d/>Ȏ:mg��Iy�2�#Z�i��F�]b�N�ى�g���v��)}��Ѐ�	�g���(+S�ZB��,8g��8?Ir�dR���]e7�z���=���s�567ʮ֘�Wg���B��BC>ʔ�q/K
x���;h�w�),�!>�5e�tY�:��֌�/����n�E��Ͷ���!�T�~�p!Z�.d8 gP�i�y�lFNV\�9��봡 e��>��� �.���$�yL@^����S����\4H�~�!
�{�׃h��*(�F�D/����3o�H��"�C�)�~�&��0����^	��&`�<��Cq8 ?ع_9����{-�}(�,�L�`q�*�z�ٻ��V{����ǘ3599$�a"L�lJ{�l\	���(ʙ|&��;n�q�R��RO�l'L��3�☞b����.$e�9���ɷ�����l��*�٠�5�XSk�+rC��n�K�S/:d!&� 2 �`xI��P��c֔p�&��X3408d�����{f}�M��h8p�4�k��x�� o43C>��a�/�J)���(2��(N_:PC��]��"@H���3e��T�	��:9����у���d��$(��E��=~�qޑ��7��R���G������'�-�; ��;�1��l*˜K|��p�{@!/�?�+�ś䇲Q�.Ň?��Ӥ��Lј�{�'!���URf�
oMֵz��^�)ŝ�L얡��F�R]B�Li`P��Y�Fe�B|h��	�À��v��	;|�>x܎>i�N���Rp.�鶾RVDCS6*����Ф������
{���p��x�N����#|�T+/�x�����}�ֆ�07�033�^w�^{�w�o���)��Tv�@���t75�SPr�����G�~)��k�Ν�`^�w)��w�r��������(���T��% ��qzPw� ���/��ʖ���H��%F�|=��D��7x�x1��5Y��q�?�E:�^���SYfeR\��s�:��\lX��� <"9�D�Ҩ*?m1������"!�+���<�, ?��d{� ��b�2d�<FB	s7e�_{�k��;�=1�Y�V[_c{�����]v����Cp�W&�'�=jLjdP�D�)}n(34n	v(1N�a1$s���Һ�9aB�Ba�,k�h�Jf+|�~vZnRx<=I٪�2�������u�Zk[�`�u�����A���
E:��]�����6�;��'�z�����O� c�m�ݙ7)�ܺ�a!e=	}F�����Q .�Eh��N�IU5S�R�lX�ܤ�6�2��Q�� \q"xz.,'�CF�<^9�/� y�;>�ɿSC�uNWP(�(�q���h-��t�(�[�#�ވO�J��/O�H�)�缅��~!�p��@.����Nx�Q�Qt�F���t?0� woldݳkm�FNxm�{��ۗ
w�69����O��Hi�s"�eɸ�w)4�P���R�����q�9u�ێ9kG��G�\�Wʊ��1�������g.ة�g�ıS~�A_o�����N������K��C�O�ϝ�rs�N���)O�b�� ��~M�쪒��Ԙ�_XU[j[�m����֩̔S>.�3���|x�f�|�pC+L�202��4d�=��?��=��s�{�ۏ"����G���%�����Lӕ@,�&~觸CW���i3�Gӝv�H >H��#���(,�S������8��׊e~�ȏ�&[C������,n��}yT��R]U�#�w��}n0s�[��N���*��b�p��-oB�'#DǤS���y�_���'�T�o�J�?��Ձ���,�h��	�I�JLٹ�"��" 0�IC�;<��F�*W#�����������c�1%�#ꅀ9�KG��n>Ϲ|�+�����$��^Ʒ~ʰ���T��r�o��P#E��eQ9)�N��h2�E��,C��{��f�oP#�519j+�������&k^ZkS��V�Tgm˼'#ON�ؤ��eňİ�pOo�p�~��=�cܐL�\_�d�-~�	w��J(?��/�׿�����~)��K��5���<�_䗼����#�؁6�W$��,e��^�ІFcw����ec-�'�.�96�zI��������M����V=pƛ�_��2�ŋ��t���bZ��&��Jlr�GZk༒��v�����.�W�O�x�8�:}�'xAu�ly�diy}��e
|Ny���n7l���4p��-_Νs��2����)�Rᥔ��xM�N����z�쉋Rbm�O�ɰ��	�Y�*��� >�M�}�Ο=�#'��K{.�ؠ:S�C�Ayi��]%�oR~.���g�gQnN��1>��fB~�h"��|`�&)a���Y���ި:g�����`�73�F�F�+Cqw��<�6(h���p�#�]+W��nN:��b4����;4��������߳��?�=i_�җ�����������tF�p�5k���>Os��L�u��zF���?4��2�>�����@>���Gl�aG ��#��.Ƈ_���E�5�k�4HDp�9*�k3|}F2�:\�,qa��[��T���T����x�73y�W������"�e>��ȳ3�-!z�p���"b ���/�#r5>2�C?�Q�w�5Cnk[����Y�5_3C�P�|����O� Ѩ�)�0���r���S��b�Mmj���h�J��&���@�|J�,0��F��p��L��d+Fb���4STI��|�����Ɲ��w��6lX�=���r[ٵ�V,_)�ې��	1��662f�Μ�c�X̙�f���������Ʀ�i�Oz>p��uw_(��E�K�·�}�
�i� �"��z`pЕ���%�lG�Dկ|�+v���t��#Tk���_�@p�ȊG&w�X}x� ���P��¸bL��eJM��W�hS,Q#7$�i�����O���zGX��1��Fm(3Aә9�4h�#`>]	|��.!�y���b �ػ��'x7��̕�&ۡ���am��T�(NK���&h�Z���,�p��I���3����~�8�΄��j��Z��Jn�g�o�1U��Ē�#*�x�E��S�8Hi���a�$,�e���R}}�v��Y;z���W�*�����P ���ds�3"�R��Gm�x��o�d��VSώ+p���4�|� �<+<� ݆ m��/�HN��~Ȩ�*v�=����������/���k�O}�����t�.�����i�|�F�%uZ��S��>@�b�dg��΃z��K(g|����J����D��NL�hU�I����w��ȺC�5�,�TH �T�k��`�r��J���=	)��H՞�'��@������n�g<���!���5��0Bĵ�P�s�W��{U���=8N�����	.ctlh0mq���������mVO���_�'�z�4L�(�T$D22vHS���5r
���Ĭ=6�����T"���{t�o@��l��{cG�#R���Xꑕ�P.�Bė�̑ϩ%�)�tb���*���)n�6o��\�;b6nܠ^���c���g��ě%6��#�I�C�8�opp��I�A�����N�~.�S�K@�S�i�tR�ƩIF8�mp��yM��D��3�1���箰�:��\���}�Y;t�����(�?��AS�z�Y/�KA H���х`��I��2gǏa��P�.rr3�\idĢ��~���Cˍ~�s���8q���Eu#.
�"o��+sI� �\���<I?�*����x9�O>wD�A�	�a<O(�x��b�a߾}R�Ԡ�Yv��f�WtxxLy9
���)p�x�gd?9Uf#C�����S� �Ȫ�"�k.��K}ĳ�&��իS����q��� ӘJR��n�w<+�U������4���H��H;�.���N��g��"KTW��AN_�3e�\g2SR�z��Z��;�n�A���0�~nke�������bd��ĉ�~m�ӓ�z�{DGRn�].e�?s朏̜:y����<�4�8��g}G���!�:��� ��x�{1x{�x(����)=�y�7Ph��B�������|U"�����#����l��Z¢(5�H��@�H4h؃H��Nc·�<�{F��#��d���˞�e_�~��l�e��7L��cz���2Ň;w6]�9/�����-�������iN��y� >�Lp�\sXrO�ό�i/�c�%�!t8%xl8a�C2�j���g��V=�wq�{?c�,^����ၬ&Ӯ)LRl|K�����I�?���4J�5��p?zFk׮���W�YeM�Rn�6��`Lҧ-�{��E�, ���ej%���!���&	
z������À2 8��3bt��X_{�	��� |AJMܣŜ?��1�����E詮�m��y��9=q���ϣ��p L�.���t!'Õ ^�2)��pG�M�p�e ��ӓR��'%3Y�D�B#�D�|�����+\�9xp�}��i_��W\����J���
��p���_	�>&�Մ��$�e��/{�o�M�(_�C~������$����R���vgx��}U�4ڌ1=H}�x���#3=]*u�MZ_��:DlkW�~�&m#5lFP�H>�	"F)�I��G:�7�M��1�/���
+�԰�C=�kʌst�빑�rs���9�m}â�I?�A�Bn�	%�Όd@��(~�-7��}�}][�I��Z�Z��&.����I����� �]�}cĶ����Jq���(�Yǔ(��Ag�p�
t�y���'@���c�f�{^�,�.�\��<��竁��9�u��D�.���|:I���%�K07����;����x:�2�
���r��y��p��,&�d7>�(��x��_ҽ��]�[�­�=�j� ^��ޏ�WN���ܫ�{�{�{��7߲�iH=aꆵ4,1�
6'�2��%V:4.�M5֌����l|tF
̌��)��9:0acRdƇ'mBiBO����.��3������|�]����c� I�R�D�8�Jf�m+�*�4��ٔ9LLٔg	3��I��|�\��ƍ�m��m�bE���'X[Wm+:mYG�/WE��ʉ���h9l�쐟5��j�7o�f��m FB�޺����ʈ;��+4�����; ���h!|L=L�6b:;�N�]�n��ܾݺVvIqhW�2�(��|w�_l�>����:��06�b�=�i)$F\�o�j�-}7�R�}�~\)�u�Sâ_U��G��x�F���f�Css` �
?�أRh�w7A��좜L'��SŰ_G�`�x�$�����E&��n�&�]ad�����)#u�YB
���*���6ؖ��$�x���D�T�Lq�h�xK��
��ɉOK���1�!'��z=����+�a����<�.�d�`���-zH��1�W&�p>�����ĕ����Q��Z���f�:BR��,�D2�<D�GT-�aX3ǎ.���HI���kn��۾}�_��r��u�5�'�Ai�+Ъ~P�Y�NO�2��:*e�����Dk]ڢ�S�?�{�bk5�;T6���%?��|�?҉Q&�:�|%1� ��\���0aO�3���4${�CɋB�/����)�k-)]����Ǔ��D�Y*aw% ~�{�?����k��i;�P��1g�.��j*)�J���[@|�D�Q�������thpX�S�,�c��Z���������ߣ=���Q��[��2u�B�	!�;�dA���S��fՋ�)W�E�.�5�����}�z�B3n3D�*���q	�	).R~���)�g���/�YϹ��e�#��Wf����E;z�"�
�������))e�E�������uu�y�:۲}��-o����ּ���o\g�׮� +��bq��D�E~Js�T�lIy����ZS�R�UkK�$�Ⱥcc��\ePL���+p��������r���C�����I��-u�ʕ�z�Úz_7q��!{�ɧ]�鹘������A�\G��l����1�U��1r@vjjB
�"W�Ro�E�XOO3Z��hZ���İ�NHy�H��8�=O#iw��K��2Bx��Y��;����:kniU��ڝwީ�-��>��=����Q�i����ح� <����> y�[�P�^���?a狃�Ц��r)Ia0�h���:��م�sV�Xi�׵[K[�(��gZ�&>��,�ӎ�]u��{�Q=�c29�����κ�
]�P�
MeM�/$��P.�N��
�&���^���F�f���rFeX��%VQ��KF{ʭRi��TI&��`�:G��Q�A�ǥ���et0�OvC-��L=K+$�$X��&%�ƛo����<�n��Ȉ�v9�UX�"�
�����_�qE���׭_/�G��(u�&Fʣ^1DN#WQ���:]<��	�:�"�A����Ҏ|��F��}�`O~(o�xQ�B�N�<�L�ۄyy�	��(<=,�
�)�W�~lG�7�J
���o�)�B1�̞<\�||��J�<����N]ث�`��]��p��ݻۮ�a���s��p�pʊ�6�$d���:!~��4UU��7zSJw,�h���FglD=�	��������7hۘ�9!�AO��'ޣ��V��z��A���`�~D{�L��#�Vr�+�����*R]�OO&���ںt�o�
��ئYnM͍�a�:ۼy���p%ڃ�V��3?�b�a����Li��j�浀b���\T��/�� L�rC{Sc�_����(=����g|ĆчE[�s��Ç|;�cǭ[�����I����w|�E/}Ó6�^?����R�EC��Q=G������!;��N�<e�N��S'O��� �>�������#�z��C	)#5�˖9�����>r@��)�C1n��o惰/��<�b�k`��	��P����F�:�l����}�s�N��\t;*�+Dڥ��ӗ}�p��I��;�� �����o㪋I��P:3g�_�ꗗ�Q/�2ֿTrTJ �o�d�仢�T�U���$ �cz
��)g�(u>��ʰ�GIb��S��8�0*}).�b�8�Gr_���j���5zg�Za��ʚ*�޽e�f۵{��f/�� �~n�P�t��/�E[�1�������b��D*��bDC����ł�3��B��
ڻ�@{��6�|��(�<\2��y���� {�� 21Thh� bA�y衇��h*��?�Z��AA(��J _�b����<i���<��x��7��^5�f8�~y���fppH�g��n�[o��V��4�:B010�0(7���t�c�C�;hׅ�4���T#4�htH
͠�	�4���!S��nz�,���;໩�Yِ#O�
ni�C1�H�/H�;=+�q<�,��_���܈��;8)-���0e&�S�#�4��.��ͅ!�����&�W삖�����G>������g�$@9��ڼAd-�D9`����E{��4<��7��zd�;ƸW���� E���1)�G��bs��������9%�2.��y=���[O�P2�|w�������w`XJ͈]�BĨ�X�ń�>z��A%�cǏ�y����g�sE�o�O�8mM�E�r�-�m�Vod��أ���NׄP��	��/��[\��ap�7,�GZ�a���q�wa��y��a����54,���'����5��FN�B��O��/�EQ�${����Kldp҆��L�9��}�D�s�!�%�qsem]�56�XKK�:⫦z[��d�ږ�R)��U�gZ�ʭ���""[���`�J���h 2H� ���wE�D�;�8|���&÷B�ګ�z�d��U�>��h##A((�(A�  ��FȪ�Q�����O�iQ���M�6�F=�1��b�o��#o1H��� ����|�P~Icժ._���au\�_)��청�uk��N����A�멓���b��)5 ��04�,��"	��a��ZfLA!ys%0_���ߙɓC��B�R�@!?��fh<����6]��ni��U��؈�ر�n��6ۺm�q- ۢ�!}n;�Q*�!��`'&V��=l�F��nJ��q���͕��HQA�:����B0	l�(�O�*�'ޓF����֥��,i�3	|ϣ~:R��熟;�$b��3!�U��Ӑ��A���L?�5\��`�4���o���w �wua��x�A�0g��K
ͮݻ��^z�%���Y��7\�s~��Jg��Ip3*����g3�:x�>lgΞ�s�����Թv�l��:�c�.��i�9���`'�?#�s�|���Rr�md��(S'��_��^|ѧ�P��04���3g|��i\Pм���e�����m��?���~�>�C���>p�D��c!�W7�рf�O:?��FL������F|�BNL�E��yu�u{}$��N,�e�f���S��Wʱ���a\�`���^���Q�ov��#�'!}���q��0�Mu�"e���VJM�dwUUZu-�TV[�:���~���;�8��k��%ܭ������w���������XK����ɿ�p�_�!��Q�����3�I;M@#�7�E������E�vP�����%��~� j�X�](�/��k<�o%݅���[n�g���%}����R�ޚ�D�+]��*n�8�6,�RC@.�,ߌ�@D�>����BЬY��{���RCEE<y������J���)6���j�J����	NbM�:Qb���kj��/]�.'�y�}�ڎ��lY�R}K���A��/���/���իd>J#�t��)���Tϙ��i��G9|IB�&G)�4��x��{O7���/�m����tb��"?���亾%��P����vQ 8�C�A��y �#�(~ٟ��ɑGzSI��qM;�`6�%&!˚$���FN�|G�G:��C�Q7�.O�ŀ�7�N=�IG���JO��:y��?�=`���~��i7����)&g�م�n����\��^7C�30b�C����;`�};}�����z{���T7�3���_�o�<��:p����1�&�F��hd�rΨ��ڵ˷�ra'u���~ַ���JM�/�����o��6m*�,t�n�p�t����ø�/�B#_����ݪr.W�c��5*uR�:��=F4<6eOJ/���1���p6Ф+5cCLm%%vj:Mk��i�eU�Ij����Gf�TTr�B|�q��)n�Ҏq�
���n��Q`8'��r����o.�EY",���YG�Z��>�:W��5El��Ȉ�j�K���߬�+U<C��8�G60e�p ����xG���\am����i�e$�a2�����B>��w�<���[�_>ߔ�~�:kmmQ���2Sj�>��.ׯ[+:lJS��Rj�0��R�,\ʝW�G(��b`d�T���k�8QT��~0�W��J���f���YA�#L���]��#����Q�3�(�w8�߸F�O�8.%���O��P>]��H��+7"@��YG3��bdx��X���'����(�J��G��r�A�áw1n�潲�BOzrV�Pi�u��_��yz{UVר]}��	�7��p^J�X%+�+m7g4(�X��+=��2��i6)K���ũ,�lin�;�X#�z�j�ȱ��9�q���7 ���*g��Z4����;�GO�m�L���(���m��j$�bC�
��-�(0==}η`��(0Ǐ��i$�[��D�ɘ�̱��.�ѩR�һ���%6��q����L���T���	;t��=��v��)O�i:B((�����8w���?MM���Q��������{9�_eJ�;&��x����v���C�<��~�-�2hi> �/oD�`�.m-�7�9�$0���Po�5U���D=��j���7e����VV4�?�H�^�n%���K��\i�֮�B#�R���0z3fS3#�èb��U2������q��JQ�,��i����z����z[ѵ�V�i��X��e[����k�}��L��Ώr@AR�(�����χt�ƈ2%��
��0%�b�wSS��Nߺy�+��x�0��>�4A��e-n�9o?AS>E���M�����y�R��<��w��#��N|���e��3τ�9�\���2��!�<0la <�	)�yB�� ���	��1�Q�`?Ъ�A=B����e�o�v��ݾ�&��LK0��8�+m�$�Dr��0c�@��,4:,��.���!��1?4w�𖖗��wL�������ڗ��Ҷfkh���R�L��:	���j��j\�ut6Z�Fk�lP�	KNe�)MJ��.!ɎR�zk�\�����ʻJ�eD��\��g+0Ѡ(���mY��sZh(Pt�6��ƐƑ�v����|���1�/�yR�L�0��i�,�e (@׿T���î��!�{�M������r5���O0)%�6 35Sf��S�?<fC��6<>iC60�FNJ�*Ҥ�Hi�4��M)c�s��J������S�ȆIy��`��{��m�U�5�7.�W�����F�����0�N��h�ΝK��}V���ӽe� ��J�B@<a��Xl�44D�A?tF%#��"?E�d$���'���x�7]Dڠ�B����A����Ψ�n�N��T�QJ��D�a10�aZ�5Zך�b�2k�VVPd���1��xg�G^�7�sFx�)�u9*�Kr� wO�[Y%�f��e��Zk]k�lϾ-v�M{l��U�]ܬ/ņU�6sC83�4,nF�� 	�J_J#Rj\�Ή�DZ#��*-R�n��F�@]@c���0��z�O�[�X܀|=-D��ܾ�!�N����2ԗ2�ܖ��.�5�u�0 "X�J� 2h�h�����KpBH*��㷘H�p0y(�ϻ�����'o�{�q!X���5Έ���4�t�8y��޹s�m޲�V��ֶNl�E��I%�%PHH8�D=�Rp����#�x�n�b�
;���{�����.�R8�
Y���
�� ��C�bۧ|��c�b����T9k�f�κ5�$�8�*԰������$��6#�0MR�Rc�q`���P�x��G�����M�x���]!dWe���i��a�!Fo�^7~h�H�b�N���R�Pl(�>h_����Ο	��oZ�D��;����={�؛��۾s����M�D����^�y��X3�(��5��h�oT����kk�m۶��Jlt")�S#M���[�|�o1����kk׮��/x���P�(�W���R���7΢����;ia d�+S�?1�0�&�3�gt��=�Q�]{v��]�ݍ�v5I�᜗��76�L�QO��a)�2Kѱ���.N#5�|���Ԕ�-��Wu��Q�tP�Pf�|+{Ȕ�T�GN9�^�'��9�ו*��Wl�e���)N�ĕ�e���4HACaf1�A�Lg�TסVJ� %Ry�:pC�i�i�Oa��n���~��Lޘ~b0����bC��LMS�1�&y��܁��b������ë�_����I�WHyF�9|e�K�_ .����DkvPvv��B�����x9.E�)fPS,Ƃ0Pj���o�����1�;=,��(<�0�Pl?�`!�k	��+�c���D���n��A1���#8���MñҚ׮Yc�v���7lX��P:f9�z�p��}�� ������a~]��L��Q��G���!n�D�����J�ڝ� /����K
C�~
�EC)�؊2�2.�2�0RX��o�	/�FR|�<�%�T?Y�Wح��Ri����Z���陹�o,����q��1�J�4�
��{��w>���{4��kܘ�9.�_��+��7��Yq%��o~�����M�W۷��)7�p�]��j�wٮ];m�����m'O�P':�r\ݵ�6l�`7�z���o�;�S�V�?q���3Ov����Q%�o��f�;9�R�N�#�(9b�2a�(O�<����=&�ǲ�w�J��x�QJ�y*~R���ʑ~�7o�뮻�qN��ȶ��Q��wg=ͤG_�#��AQ�I���霕<�x��i[�6ڲ�f�F�R��:@���1��y���[q�;?��R!'�C�y��{�;�+<�G/����	�1��Kֻa8���X�Ky}��jn�&]� ���d�*�YR,*.�,4�>�F���d� ^�������8���=���3�p����x�O������3�.D� �U�V:�;�m�׹UN�nΎ�`�Ӿc��r��j�� ��"�b �
��&��p�87 �T� �?o��y ܵ@�
寸l�Ұ냆����ӧ}J�1�;�3�>MM~��G��OmA)F$Iφo'H	�H��$?�K};)6�z�D������Y��.+�b4��V�F�E�Ό�Ʊ�aJO*
��C�1��l|K��`�P1ߞt�B(����$��̛���0�@�2J�^;0V�\a�Ww@J�*���r庵��KƔ~�����}�SJ;�������c����]Ny��<L�<x�E���w�}��}����o�۷ٮ��{s��z�-z�i����������'WWW	�N�o|��~��#������[�qf���g@>P.Q���u�=�@��w���y��F�.WW���`�)��A�^X�壉�J�p�<F<��L v���t`�o��#�LIQ��98Rh��P��, )�z�Ӕ��U�wx1AR��ٺ���Z;Z���Vi�(LI�0_�/�u�v'��5�g�Oq������1�⣽��Z�<��R)1����M��E���|E���-U��}T0p�g60Z��@y�}�'����S���Ձc�1�
��0�x�?=	�Ȃp�0��|\������W��@>���QP��B�i�Ua�q@��2{�s�rr�!* !N|'��BA ��D�3� ��#7�=��� y��,ip�2�@ 4��}}�+E&p����Zv?��{db�4�����M��:9 ��b1�Q��������j��@�T�WXQ)?�T�3N�E��c��";�ʄ,����$�d�=�-	�$�|�E?�?��ۼCh)��/��x哲@vz���$?דw�H���������|y��|y�
~��x�F^"�@��;��|y��u	P�b�ܘ�gx���7�l�|׻|ؙ5[������	�gϜ������)�����?d��g~�n��z�ό�u,�=�v���kE�l*`�����N��K�"?-���7e�:�Yv�D9�fr��!l�w�W�V잷'��Fz؃g��O�u�)���6��֥KE�U~�%���A���QN�8�z��S4�	EFy�]��(((4��u��R��O��)���
�P-���2ᾂQFlş�.i�s��)�O��7����
�xZ��dV�
�bSU�z'^�1��'���>�Ʀka�]�dP��P%y���hO����˰�q�@�ߧN�rZY��L�~G��/=��(}�/h������羡�D�N������������]���/[ZL�T:Ǐ�����2�^,HT���@L ����,������GGF�X������a���/�j��)Μt�rq�-�K�>��\='h�!yF*�`�t�j(X��J���9o�C�7)17N�rEg��K�B��(8�Z_e��vh��
)-��.�WϫNy�O���%���W�@�W�C�0AJ�`��O٢Θ�V�R^�g�1���HoP�&;�(c�9��¨l���#T�A1M+�O;�o��ϖ���ؠ�W��L�� ��h�dڔQ'vr�J�C�(<A�u�P]�K h�J!��N��,����c�ٺ,���=-e�o?�7����u�?�k���?�����
O%�l�r۰q��Y�^�T�mQ�Ύvўt��Q��f�AT��_��gZ�8߸Q�:	E��S���ȿ������eV�p a��#����=��I
����(�#�TAIw��w 656KT�U�}>"��'�Q<@����3)�F-�"p֘�@�_�$�⬶V)�U��p�״UI����ʌ&��j��ؤ��S�<��DEܤI���@��?k�$k�13����ɺ:u�X󇼧3ň/2�3hj�+�F�K����si��v��XC���:k�H�Ӈ�3�Mr��)���������K����I1l�Ə�.�q`�FLQ��@��3��H�)�����@�16I�-LO`m~�K�Q,s��_-/�͂@�nU�~p�heI��W4�Q�Y�@Ô�=�+��W)�XM� cb`b���yW�s��Ѧ���b%�,�˛b��#�6,D|�0]<1������a�qᆡjr�a�M�|w�/���ub�&1�$E��KT%�=���(�
��u����Ii���bSGO�Q��@H��qTzu���J%m�!����ō魬����yp���h|���m�;�=��~	��E�I{4�$M���������x|32�a<Y�Dj>��\�~`|s�ǔ�Z��k�O(�UU���2\?12:l�?�����������?��}��d�����/�������}�k_��{ގ=f�~������8/���&u�V���O
��y�V��JâT�o<�MC��ψ7o�{��QFD�8	
�aB`|���L����>sʧ��vf���꣦JyJ�^���1��/)i��RJL������d�Ա���{%{2r�Bd��F�:9i�`zˣ��=mZ�׻��Vi&���]��i
��8��ں�B�!�|�<��
� ��S������1�R&��L�S��*}����t �FgڤPo߹�i���(�[������9K��0�Į�tLE�+7��🙀�; �0 i���33����̥@�!��S��V~���b�M�Ph3�/���U�`�� J�MaQlh���.�����0?b_�J(���B���|yZ ��B��_�C�΀�Ɖ�R�gG��͛m�-�vM�����o��Dwzb(Cf�"=�۩~����	5�ﯫ����*k�bé����46�J��R�a�%2��Q����,ŕ�iJ�2
�96,V:suyK~��$�w��L���K oE��l�C����F5��ӗ�
gM�M�c�%�S9��=�:�hx�/�0ׂ>�6�]�{pMYa���-u��D�==��_��}ꓟ4N� >�Q��x�~��_�����~�7������ߪM/��^�����OI.�e���~%��G���$4���y�h_D�¼Pvҡ��O�B� W|���t*SwL��׿��-L��MuFY1(�lYg�	���t� 
 _wI�st_�@;L�Q���*�0"#B2����Hq��d*���J����:�1���-Ę���w)�C�G&�MU�G��a�!�5Rd���a���b����dr���*E)^A�z;^���ʙ�)��Q�H���R���舧ɔsSs��08�u��hQXU�=���F固����6n�Oks\n+�W�FF#�7l�T������g&�4�yA-Ƹ
�2�m8J��l9��^ʫ���P(

�
���Yy�@䁀�3�����*"�6���B�#o�&D��O0�wSc�!}nA��8���K[�ZCS��7%�K�8H�1R��G�+�BP�[}m�L�5���ZJN�ձ����bRzKf�p9�E��[J#����g��I%gt(��<��RӜ}���*{��� {�J�����/	;�hyI=Av�	���s��bj����H���#l�����D��?�i�J4t�r���-J�L5��b�I�U	��J�^ս��z>w��}��_�O|���������K19S��q�S7�x4�� �|>I7dG��o��r]	������4�|�.��KF�a��=�^.j$R91!/�5���Ӡ�p�0�b�K�ɧGj�q[�R����6�Gmd�J�|�
�o��~��
��H1.=gٍ$�4]����O$�uSPf2��_Rx���8��`�2��*��f����n\��h�iTP}��f�^>�o`E(;sF�y���q�-����4����4��u@]�1�N�N�T32ͳ�ѳW���G7^�z�8@3��n��wz� ��[����e<��_�=��>O����<2`P Fg���=9k��oފT�c^�. �&&/,^My�v�.Q�|À�H����z�Q$3��r���</��8sX=8v)�QL���rP~	�i��1I��,��l��>7�^��YSS��T�i�Ĩu����Hĕ��h�[B�fw�W~*�FQ�/�#����$_�K$0��`��Ch��/ʚ��>���=ʡ�罐&)��v���O~Ci�@����Ԝ���� D��L1�V(/Aӑy�^��;.ʑ7��CG�MX��iU��uǨ�+)�W�����4R���2<�=3��d�h��D~�>��ń|���e;����y�ۍ�-�6�q�S<���x&.F�x����ѫ-[֖F>�QL�&ġܺ7�E=��q�'����bJ����"���SC�yPO5�Rh���ڔ�qA��^��ǝ),s�sƙ�僧�A*�mx��C*��[%%����b�g(q��w��G!��3�"2�h�x3�%���l����v_`���(�i	@�_�6�"�8�q�;����h;x�����(�&�������[�q���hǗ(PFϕ���y񵜢	ڨ�B�ְ0v	��s�D��[����Jp9B�V��/9���D�F���C�;c_u�\`Y�~PT�3zor���i0@��u�9�.�oR:h�h�PhJe'��M�z�%Ur/��GF&��'�#��)�IE"ЙoZzV=�Y���tSi�!͙9S�i�Z��b�RWh��}��X������$�<1A�qzO��_�s��1���V�=Aҿ��+a�=4��;�RHA�2M ��/z�4&�mQ��\)m�V0?`f>�L�S ���y�Um��jTu@ĉ�����x�S�Ӕt���@��i���|�PN���/��� �A��B�|]8�oǡ��;��@�O�����u�� #L�p9d�k~H|�#(����+��H�x����,�yq�$�ʁ���s��Կ��Uo�?YǊ�!7Ї�'Υ�ϕ����c��܅�r�艅�i������K*w��J�knjp>�#��\�Z_ߨ�8�/��h�֋�9";NA���Z�vik�oG3�s����Z&����M�U2W
y���@6�$���僚�]c]�ʕ]�^�Q��
��E�ʅ�h��L�� 25�T~(: ������B~^	�a.�i�g^	�#ܘB�bs8''s� O�h3�̓�����ɚ#�{pAX.V�tv.���К��6�
�xv�������_(�+(j�J�hM:OBiZ�JF��V�[�LYY�t���0�Pz�_Hsd�y����gl�LO����%I��z��'�5h�)��Ӣ�������TTʖ��y&�<��JCъ��J�
���V,��C�~�>��Nx�I������`a��˷Hiz�e���=�;v�j4�4���j�i4�H�z�0' ���)�2>88`���HѸ��\� O�+�k
{�}k�P���h2�Z@�C��>�����)����ΒN�Ax~D�`��S��"|^��ƿ�>u �	C<�t7�#��/�)u<���E8!�����sv�ϣ�=uP���t�Y�n��Ϗ�f�J�bR6\������&;��zJ�¯P%:g��ŀ/��wKk7���3Si�--���{��h7JJ��5�r[?��{�[�l?��?l?��?f?�?i?��?m��g�����������������}����^���y�hX�9L}е�ne��(g��_��j ��g�=h��?N����t
8u���Iԣj�X�I������*B
�{L��=��2�&1g�����+�J�8̷�+�£�0	k1��໾��{��{�������}�C��w����w؇?�a{�{�c7�|�o��-��0�P�֮]�a>��ؾ}{�>#v�pl8�l��yg�8,&�¤"2�_oX�p���@	`��V
�7$���E�xDPQ�I�0DL5�� ����-�3#�G��%���hL2�CϜi1������w�oO��oV����-d�o����8��~ڲ�<�O�H}b��v��kW;]h8x(��t�/?�$�&��o4֌и�Ǔ��w�P�)ߘ�4�b�F�
u�s>�W���+v��Qx�iHJ;x|��Q�\��g�I^	�E��;v�@q���N�bF���{\��by���M9�q4���<!�_�y�#�Tn�̞Q6$F��ۨMͲi�O2���Q~8�ƕ���$Y���t�R(?������ɇ�P?p
��+�3ŗ63ȇ>��?�t
���?gP���(ꥭm���Fkin�ۧ���鋯}�F�*pH�v�m�������������6{����ͷ�l7�r����[�;n������������o�opڌz+�a�����Յh�P�E���Va�<,�/�<�]��w�����/�w �珿�\+H���@�h�Y�O��7�#���P�!2�1��}�@zy������J��A�ʂ�BI����G~�G����g?�S?�m�'Z������~�'ҕ�-[]Qd�*�F
��9u���k��?h;v����m4{o�א P�W?�
�!k�L䒬��B��t�"Ĩ���1��]Ü<L�KUC�(7�	�9�!���?��]�Cq�vAt���Q~�+B�&e.Jd��8�`(8��9p��_�l�I�����qr�ȝ<)?�R�d���%��i>o`��y� ��W��i�F�����F�R48̐F6��Z��MS~��*A./B@&@�������A�v�CO@��J!��a7�[ �#�(�w�DO���L��p�����%�R$��;�C�<�1�R��.\�>��8�^�-FH�4���0�<��?*b���lDR�<n�:MN��>�ՙ��	)1�e�mt���^�}�MM�f��S�(*2R��Y5�?����<��R�Xå�J3);I-Q��M(F�
E)�7*O*W�O�q��[@��C0���B��̙=�nZ�z��~��� ����w�y�wF���kk����.e�y4Ey�㌮�e��d�M�7[m���3�s(�/�S��﯎~#��̫�H;�/�G��U:(z�G!U޹p��E,�@��2����s5 q�U�<2A��ʋ�aP f����{�����_��1�@���B>�@������w�u�]�G��S�����jھm�����˷f�{�>z�{�n�	��Z�nӦ����h��-�!�X��q�Av(��)���{Yq���B�Y06@�����w:�SEB��Qz%���N�N|�tb��l�q�\:���pL)`���SG)&�?0?�x�Μ�G�'���U���)o,�c���k*��FXP���EX�rM��8����r�R�pӀ��Ďp��[>¥ 4��B�/��l��������.'P�������$x�:�3Z�����:	�+�D�A7	"�x/�����w4P�<
k��5��d��CbB��iPʣ�<��<Q�����\y�b�45��8i�x�	O[9,�/5��O5�z'o\3�MO��1
�/��F����Q�R�t����W�uΟ�Rhf���q��B�|jH� �=���ʜMi)i�C��䇩�4�595�4ESJ{\�$�|��^y��+<n��2zلd	e��Y��YEO�tx�w�0�C ���t!뛬����v�ޥ�ٍ7��y��N�<�g�8~=�#���Nvf� �H[7]`��%�5�5h�e�O�������=���@�Hm�!�`d*a�B`��)�ɯ&�+��������?.�c�%%�R�n0
AO�.�`H�poݺ�>��]:�x6n����f�0��0NprO����K'=d�v���|���f�L:;�^��l&dO/;{/U���z�Qje��[v{*\RT�a����	��r�op�L�w���0���OO)(y��y��Ƴ�lQ�0�<�bJ����!d]r�(�� %O�SbޔnA��+��b�ݿ&|���(�mP���+�۶m��a����G։��߶u���O�������������n�]�>m,
e�ʄmn}'zx~@��y��i?���y�����/c�U��y��h)��7����?~������<j�����A5��%d@cc���q��?���/��H:���G44^g� �����}���)��Ĉ̐�A��͏���L��QZ�f૔������%�~�VG�N*3<41��#626$�a�eFǇ]��|� J�ވ+�1�v�M�� k%#(4D�7�z�>��O�������~)���N��Ze�W��ů��;~�����?a��˿d��_3����>f_��W��O�(����'����!۲e��ܹ�;Jё�������N����D���&��YR��1h;U�k�a��	b@��]4<��0?8 �B������|���;o�J�BH&�0 ��FCC�0��Fa*��7�a�?��=��c~��ٳ�\r1Ø�"e=�W��2� >n=�A�Hy�d�2��N9��˖�TB��K�)��4% gf��RuH�XS�IJ��m������g4.V�UH9-S�$�[Y��Vq�S;(5�n/١��90�c�Y>2CO��,�/1˴��zm8���"4�Kg�F���D�)cR���@���E��Փp��:��s���hP�q	uHxǋ�F��������kyzͿ^�+��x&L�Ƚ'.��1��ezsl|ԅ��7�h��l�����F?ix�����~�������7�ͷ�h7�t�mٶEH3�z��}��Z�TQn�ږI��Q���<y�Hy�.��g�!_�x�`q ���~��#>�w�	9�l���D>�=P���4v4�@� �It�FH����Z��0=#?�VڕB^�y��+�)�1��I�$����4�QfTV�䟆�4E�rQ.���n��Ң�R�-�aS���l���$��Ǆ"�6��㱩a��23!�xRfzH�6*w�[i*eǟJ��_E�4PtiC��d��)ů /���iR�P�%c������Cv��;z������>ɱRk�h��
�/���{�G���I{��G��_��=��7홧�����H$c��Ci��ey�4;X)s1�])@St6��]L(���b(��'�
6}�O�6�E�rUN�l"��V�8f� ��NLeà0:����W����L�U~1��.�/��@���&U0e����O�:e�gf��{�g���������x������Ç;Κ��������g-
�z��'�+_���?��G{�e�G6(et���&Y���L��I<)������&'ٍ1l�ꥹ�X�pU��r����7����i��������_x	�%����������b#���|�p�{ʥ G��G
��w ��A��51���!E�}�Ae�9v���������LxS�+��Ig�EG�C���b��� �^��3�{�G�C��<4�	�(2�����c'N�pw��hoo���z�������}�>j?��?d��=��*���5�c�ɤ_��Y=�5k��.)���랻��~��vS���9W	`���?��&�y63aG�|\�\�/ϘB"��47d`�E�d"r��#�2 yH��q��,K�g��H�K��?X��Rc>Bꤑ�[a�R��|G�D|n$�R�=ΤPH*�4�����O�2�x^~��p$�G�RgF嘐b3)35��;�t%��U�� =ՙ
����=�񋢖��}�lPF��\�r�oǎ�޾�>bV*�V����o�i�~���ɱ	����I�s�d��(3�\R_(��5u�b�	��\�rf!Hؽ���N���|�ENF���A�&^32�V���*C�� ��
E�9�t1#�0n��@�d��nE~��/��!� ǁ��0�+�ӧO���{�s��/|�������B���~�8�� и6���7'�>�����3�����������<y����6#��  �,�[D�`i�z1�K������=������Ug�#661�NJ������9P��T���}
2h�>��$C�!�9�RS�/�}Q)>>�/A�`�;BЍ�Ha�2�2�ϢM�!���3-�]Z�̨JR�G�������
'�������ɧU�U*wRz<��{4N��i���o� �3L���K�=�G�^��k�5��4)u���O��ذF�U8d���}��|�����>��;\��{�>wڞx�I{��g�ϙ�����mӦM޸!0Q2o��F������?h7n�|�e�|�2���� Q��;&�|o>5�w���+���?4�&	���+5�̷ӿ�ϛ�U����\ mq�T�&��<�����oOY$�M�҈�+�?��e~�{� ʁR|�:N��?�A�7���.�ns�O��rA?����53�
���c
�
"�9�����2P�xCo� c��rb2�g�b��I��c5<�H�앿��=�ȀC�7�(�� �f���P:�Ƨ`�o�����2�#��Χ��c�J8�r�a���q �Y�j�:@Sb������������/"P�03ƉW
�W�~���Ĭ	y��y �L�[��y �_^�|+Pȗ�[UIǙI��3 Sp��L)a�@�ݱ(�o��o�7~�7�w~�w����[=���:�3gθ&�"���x�+�R��L�|*kR�,�xC��b#A36���ĨM�w�z	����G��.'΍(ӳTB�3%JT�lW�͜�ӻI�K����S_�@P�p���dO��('�ĝ����Qʦ|�x/Õ�����hSC����f��h4:����3�
`n��Na*Oీ�kyZz���[|���s�MJ�7�RPӨ+�v:��������ߵO~��v��i�	�d~�54��pS�W����?�c��Cߴ�jc�f��u��ب��]R������eo|�}ꕆ� {FЈ���^c*��:�.��/&ʉ[�˗?�;�%�y:Y���(& �<�8�apx���P��S��/���f::���E24���x������7�]f�˜pNWhd8�W� ֡�J���M9�A�<ٓ�(��{ �5gBn��&�>���̅d�ˤ�-hXV�qm����ӿ���z��S��2:^���	�7���	��!'��s�Ϫ�¹b���$eK4)yC��9�_:��ꑶ�iKq�(�蜺A�www{���*��Ny���W�l�Z�o����nh�5*�+Dx�[e+��L]O�.��E��x����.`�hx���V�0"��Wl�(#=L�;ʉ����C�Q�I��O�<i_���|-����^���=1e-�K����O�¢�����L��{x'�\���4n��4�e��zTzgK&��LJp0��z�0��C�H܁t"} �`�B���L2a7'LyχQT^�9����e� ʄ����w��	v�HɦU���;u����BL�A�9�N�v���@�4<Q��PN-��CkR�H����Ż�c�%8=d�<�>�*,���M<�G/��)���_������=��s�T��4������~�{{z�o?�7���?�~��H���ڡ�ԩS�;Fq�K�#_�%���=`���7=�#�.t�x��PE�����0_�?������O��H��7��Qvg�/�q��� 2�@S��[1�b�'/��Sg��q��s��ƨA(��_�α�:�v����tB�c���(����!{I�g�	(��h3�*q��%y ,�}��C��,6@�1D�Δ��,�˂d�)sK#:��_
��@J#����S������6�1p��,�$0���tM�3�ʵ	��;��B9�:�1�������u�y�2|;/��R~�e et��s�e��%|�T�.%3t�|�y-aQ�o��s��N|�jZ
�@T<�i��
@�o y���`���熹R��!/Y�#ʔ�	Olo�?��XU��PYT�s?S�o�伄
zf�-����r:��(:�ah��8s�J~_�4?�)(��0�t,QkV�X

�����J����|��c}���)-?�4߻��n�[�E"?%������|⟲#?9We\���'���p���,�c�0����8>��ZA����k�ʕ>e�b�;�����mo����-v�]w�t��~��v�7��$�;����^��
�s�=v�m���2w�q�����}'�-���;�n��V۵k��ݳ�V�Xa�Ξ�_|A�|��D�3#����4�'�}�!������g{wﱛo��oeF�s2b�Äާ�'��؁�\�ٸa���d;w��)+�ęN���!����bQ=3׬^c�6l�u>�7m��{�z8������}ڑ^���K�npwvR�;����BuW=�|�  ��IDATL���Pl�?����q�E�F��,�?h�Q �s�p:A
stv|�G���<|��!�P�u��������|*z��6���դ�lP^�F��#`�q���)����0@.��y�"|���HM�'yP�e����B,�4T&����Q�L6�	K��X���ⲍN���f=`�3.�r�O�S����x\�Iݢ� ��su�=�P�J�\	9R�6]�ʚ�p� �%�w��Y�Q��*�F�D�����RT0� ��!��گ��}�_pMB�����(X {��!_)� �G�����������&܁�}1����`������K2��������v����튝�"�Ɯ����eͯ��ڃ����	���%˻��n�'�nټ��.kR��s�z�,�C�@!I�	BR��'㴗�N�����I�~]@���
H�@X0g��d�q@᜺e�h%;�ɔ���+|b���,�����ٗ�A���4x"�9$
�Gܤ��Uj�#cv��y;z��ض�6m��e���h?��_j#����o��(+=j�l����s����ٽ�n�,$'�%#�[WR�IJ��cx��@��	\Qh�o��������t3eGû�u�+�s�
<L�I��E�4�<B��	�oݺuN��.�������c��E�Q�Ř(2č]��uT�B�|G�!���" ~�n�E�S&d���|Eٹ��<<x�װ�;��p����V: �L�'|y�&~CY	��+��qᇰ(<�3R�kBJ��5��p��ɇ}����v��I���u�/���z�@I��ӥ�Ɉ�}��\u��(Hg� I�&y���MeCtY\�|�w(��NY��e��[��>s�Ž�$uxS p�\�hC^ �K�ؕʫ�ˎ(�y�2�ĴR�E�̖�Ja��"���x��e^O����6}�F�G����~��~�֯Y����~�>��O:�S�t��87��7���O�>�裶B�>t�d�����	�/���K��n>�b(v�0���a஻���?�v��Y?���DJb��u,o�7�w��[����U��ݒ������jâ)5 QS*ѯ��2���G�����JB�Cϐ�}��g�!����F^h�b���Un���;�$`>!<�G��p�ߤ���pe��6�����>�a�A�!������Ľ$,Z��_�{���g�@��u\�@/�s@�n�`����6H@1%�TNe�!Ks�ʻ~!�<��r�L0��]XdSH�w��8�0���W�-d��w�95n���g&@	î��?�?Wh�/�R:(5&�F���8Y��������?z�Ο���U��*�FJ�פ��'?��uO,&5hz%>��;u��!�b�YL�4����G]!f�:	�J9��CQ����~�1$�����q�a$�B=R�0�2&?�<PO\v���R8Fp*9H�v��rE[?�֫ƥL��x���F�0�y�I�)F=q�e	?�@�q�g����`Oyp�2�/�Q�l �8r�ul�"~�I�4 ��;�{|���!,�t �!/ ����w�(~�l��K�����>���}����XS7l���ѹ�/�Mۧ��Z<�Sj�I������n�G��wٻ�����|�v -���ᑤw�8��F
I���O/o �f�ܡOd��Wl��2��%VS]o�M��7`�?����XGw虔�O����N�	۷�:���7v�7��������퓟���Z�x��6m��������������~��>*�Q�<�A����$��
u�s��܊��-�,�������s�]�q 2@Ϳ�&����Q�O�]"-�5H���֮�`���Nm���k���q�"�@p0G=[*����|K
ó��p��b3G�"����@��Ð�p%��8����=K>��@����t�����(?ߑ'FP���s.�z�lAƝ�ӹ)�MOLI��!h.�/�x���P TL��G2���3ɯ��8�C�	�>�&����^Szb���J&�yu!�����)�\z����� �$��zN,��н�lG�s�
g��h�wʅ�Ahh��?u˓|Rwyu- h��GP$����<ґ��I`�=MF�}�9?'����>r��~��kX������Ç|�{�⏑T�b{T�'�|=|�N�<eCޣc�HOw��m���r;{���;wZϓv\J=�z.t�q�hc#�jw�����_{0�r��ß={����Ψ�yX��E�Q>��8����'|��'>�	��?��¨q�?qɬ�<�y� MI�@N��I�Ǭ$�r�=�B#�9t�;r1����;)D:@������*�=l����;7܃g���Qh��w����0J�GC�C(�y"x�����a�a�7@��މ�xB��>{�飪z2u���I�ā]q|�޽l@�Kkix;�Ys5,�-ݲM�&e�5�uމľ�k��X�iUR�Y������1�9����E�&��F�?v9!�i�l�@� /��&�2:O�Y�Vx^�_��_ q�t�$�\���,�IZ�����U�{ui~;��#5�	-���#��o��}泟�n�UWU�?�~N�-�4����R��HA0|��%����7��O��_��=o�?��'�ibX�����_���hGq���`=@\x����e��)�b� ;�Vw����HK(��^յBB�̆G���N�CyaB����0�0&vʡ�H ��Z��%�
Q��$h�;1�-����(ă�7���d��<�=�@�/R���]2>ZSP��1�D�_껬��0m�SjX{�LYI�ݰ�z	�F�񳪟�����O��ߴf!�58�+�>��@Q$��y�Yl@@"��G��p�`>�ϸ�A�M>�=e�w͡$#|�/��4r1#���s�z���Jެ+I�&S?�E ��&K>p��e�����)�U
�+�4�t��Рo?^�|�O-� �V��|z�����f}y��4>��3y����z�? yFB1Þu3L_t�!o�$�耠Xn�x�	��?�{衇<<�rF~������� "��HA��>P� ����aCcN�� ��-�7ڻ��N{�;ަo�l{.v+�\09f�7����Ω���E�Vq�Fk���@ǒ����
����
�%�$�ه�q>��{YvRz2�Ƈ��������<�z�	./�O����D1BI��K����ǥ�b�=��Qҡ��kֈ�j������1�����;�G�G��`ڱ���߱��˿��������Y��9�}H��~�w�B����^��h�ݽ /Ѧy\Y�yG���0��@�|6.�y���zȧؽ��c��l�/}���Ȝp< [�˧l��{�}�8~��)�Ԕ�IC�E��	�?�9ϋ��@�� �@4B��^���$��Sǝ��̇��J��	� T
B�ł��"Ҍp�J�g��xϻ�iGz���Iʅ��2Û�N{>��8N����E��E��K_�2�������9�=x�)��HQA�$ᐕSF������� 6{/��j�_��-A
$bϐq��͜�wN8�Y�=oH)���A_�<b'eᕾ�FF�0�z}4.��3	kv��t�����56��R5��xRgϞ��%�AC��,��㉆��B`Л/�7���ؽ끂����a��/�`���˧sO�<�:#-�԰��3���]1�q��I��)�s����8�#(=��v��)�=��y��Y;t�T�y�7#;�\q;v�>b���S'OؑcG����|����C����_�F㈾�6{��1{�'ա9(�*���#�q��?��2y������K>^x�y�ƃ߰'�|Q9�{��A;rTi���0
Evt1����0E��"�;vښ�]��P�^�z�/�#a �9�������7Q�h�N�켾�ν@(d|�O���[�O3�(�aqgMH��۲e�+g�Q���������)$��8��FtZN��8!�9:#��]Q'�5.�d�	˞�!��N�G�=g�Y!��ߍ����7�
n���d��F�?}�x��r���8�7F��.�3��(^C}���V��Lg�l#SY4Κ�z�ѧ�|Z|rֺD~� [ﳑl��X�Ε ;w�o��v���1�c�=�t��S򄌦��m���}��AVR=���<�_��rꜰY��P�h�8�����]�=��q��nm]������.�~g�q���Yo��qg�
��PUdk��|i]m�
�:�8@!h�ф�Z�Do ���0T6&�Ā��<�'@��g��E�۶m�8I�4�d�H#w��7~"Oa�.�&�H+�DAt�흾F��q�?y�L��Ay�+��D9�W�-�������/��KlrB��T~��	ϻp�W>�yy�C<s�s��3I���<��$�/�2g��ǝ{����;yI�q&�+4n��\~�'<SI�S�Q.�Ũ�bJ]𰭛�mY8�"�$xM�]�t��B��G�O��v@�H��_vȤ'|Z�C٦��t�Ձ"�ǔK_�����I)����6�Z��/WݪFs��=v�]���;����V�-��m��z�R[��j��:m�ڕ�~y���X��2�_���6v��}�m^�aW,��kWۦ�ji��jm����A���eV>5i5���+���X]y��5�ZC�軪�6�_c�]��n��z����QQ��&?�5N�V�Ω�ﶋ==R^λa��/bG�ʹ�a�"dpRQQ�w�pj5�d}�BUX]]�G��z����� ��2����ȡ����?YdF!=�%�2-�����6%G����*W���zRT���[���L�뛒��K�C�v��za���JB����T>Wβ�d�ؐ�� � ɸ�������!�+p��M�ײ�~��^�+�ͬ�3BK�;)~?w�[O��*܍zB=��xG����~�[�:�#e z��"�5�����>���?��Ї>ho��>[�q����'����:I>U���C�C�ԭ+�1��/d�e��&nu_�Mo��<��ǎ8��j�Ȍ�c���ȏ�;kg�=��RD&b�!U��5/߬�S{/^�P�^u�'��
}��$f��]��C�h� ;qP%!t:��V�gnA�@�p�h��rB�^)
���Uh��߸��ɛ<G��a� �`�Y�6~���4�h�((L%��p,|M#��-EO���0�2?(O�H9�r(^҅�`*_S���z�Ѫ ���ᣗ��	7Za�ƻ�.��d�hL�(���Ǒ�)�g��;�}�=���,<�Pj<]�����>�\r!g(2������J��\��6�]���#G���?��'���R� ��6A)�v��0��biPF��<���{��t��g��3�Ψ��T%
&|`^H��z)37��uR6m�� �~˖��f�۹{�-mn�။R6�lys��X�l�R*���\JJ[S�-������l�wc�-k��ΥM��-��K�C�ڛ�o{��-k���f�UV���*L���h��&5"��+|`�A����Rh�mY�2k]�꣛u����Ӊz���;W���@AY�z��]gg�uH��i���ߤ u�#�<�:x,�@���]���:F����v!�b!?t��!�i����l������zYgv��y�BA�Q��Z���~�,��!58n�8� �D��EϏ+$��0d�}&u()34�x�� �t�s�xu��u��o�S9�=���İ����,��9���b8SbC��v��I��k���f+S�4�5��F�%���o���zfJ��"z�>��yl�b�|E��r�r�$�E�h��������O�Q�K��:D���<p�O�@�pPF�~�Nf�"�ti�-m]�<4��2g��_x�E�ie%"}"steq�+<a�v��ZuNڄ���OXo_����%���Xm۶l��6�ik�ׯ<�,�łEQj��I�R!0.�eX��<_9�ʞ��ш3܋"���A��$� ��?��3����rU�+�˰!S`�OE�>���8"-��	���y���thl�!?�öW��n��&_O��[q�_�������~%�P�+��(�GJ+參���b��ɴ9�B�M:�W�d<{<yd��.�vr���
�ď��N�$����?��?�ܸ��<�K��^�q'�����ShR²�p��Ɵ�!d](�����g/�����puu���!Ԣ�;����N�-u.��ӕ�wa���Q]��~y�]l���|�f��m>����Ï<��0#4@(=�/⾚��V[[mǮ��ֵz�-_�Қ%�R�X6���)��G����M�{dh�������p���~B����lT����H���{{���xqT��q懔�q�{��]8^��)��q�mh�]{v�M�#�#ꫪG�ȉ
@��-�J
>��Q>(��Ł�^amYLo$�JT_�a*���ﰺ�zɡV�/��+��~�F�)-�w����Do�)W�GX�y�� ~~�Z|���2�PWW㝜F5�D�5,j�`8�b$����d�sB��Z�3�����C��g�O>�qF<n!��c~�d/�'ns��K�h��2���0s�߰�m��;�d����:O�?��]�x}����8����!�Qd9R��jN?n�S��ǎ
����a�R�'�Y<�F]|4W��B�vN�����=n���g�!e�v��M�8���R\v��\�a���c�Q�Fe�-#���[�n��^���g~�L�q����v��Qj6�_k�=��˒'�#t�j+m�V+��LJ��V�-G�.�o1 �l�!�gά����sT�#�q��3��p����p�&&��u�z�[�j���N_�!]��r���WF=��a�M���sT�+A�o䑸0�S.򈡬��r�c�v۵k���Y<e`]�?��?��>C9� �H�Jx�)�C;v��9�G���v���I^����c���R���{��-�O#�2��'��͋�J�4�%��G�Gm���HJջi�c̥K���Og�n�'z��b�-z�����!s��k4N��E%_��SЧF��l7���(������L�p�sSK�����!!x��7�Vp��_�@~ꙧӨ�h�0��V%
_�����d��OOJ�+�)}�N�79>-%��l�����P�Gz����rr���g��)�1)1���4F�#�V�����VQ�t�m�<aߠƈ^�2̲6kmiS����.������K� 4�"�|�
�oh_��A�*�4TlE�!,���J��׹2��])��>� ��X���p�h`��aQ�yytzr�D���ܲ6�+*X�JO�S�u�R}�)��ހC>-酂�I+M;y�
<�?h�������OBZ�1x.{�3�,n��.[����0)�9�Ϗ��Q�0JI��@��X�ή�n�u/L��8�`��A�*���9�?��QG�뾶�����]�V�î�.��s����
�Z�G=�7�/�O������A��)����孷��#�L���p�w+����=-m����B��!�,���[�-��]"=�'�W>�%~A��%���Ay���H���m�)ULzRQ4 �#TQ8Ʂ��Q�\�(��/vk�l�#-3 A8v���\�d���v����&�嚝T6�^��N�O��X ȹc��G�G�@>�b��Cy8!.F�/��NѦx�n��c*]~��w|P�Bn Z���'`��t�g�s�'N��
	N_P.��R��=]�Hޟ�#ʑ����o�3�d���r�s�Å@��'S�yf���rB�p����sV���{w?�.�qbXL��Μ>gg�sc��+(݆|��?%��cct{�M]Q7Q�8��_�M��o0K}2����8��9�+c����6o��t�կU�V�
3J����Zm��{������r[ٵ§vv�o������vŁE�Eglt��?���ɢ\��Ah��T�������� e��2�����-�) EԬr��_Z30�F�eY��Q���)5�}Ο,�E�4��;;Ԡ�a��`]���<��<i  ��U]�	k}��[갭m��W����ʕ7��#r��{A�����r�:��m����i7��w~-	e���[�,��(c��U4R�fdW�Ӧ�+����B��kA�Ƀ"Ǯ2�e�����3�W�B~d�,oě�Sxκ!}x�0�d� �0��wLG<��;�?o���7@�R��_/)N��r���:�z�;SO��;{�x�ǺV��N��?�~i@��}��~�����e3I���;,����������#�>j���C����{�~�{��G�'���yԾ��/�"� �?��w�&)�LG!KPz(?<d?�TP���a:<�z<�#�t�|y��={���w��~��m��n7�|�w�Y�܇Ƒc����y�VRF��h� �p;��t:XL��������Qk)i%S��Xc�6��ں[־\�S�;w�bq|������Oz1�2�˅9j�#S�\��7�#^ ��@��Ǜs�;Cs4B�!�P�b�2=/*C�k֬q��7=�H#1b�K�k�o�q�w�OO�i��Q�{�q{��'��G�F7z
_���|�;Vd��2�����á`L�P&Eb>���#�F��J���%�J&{(���?���������%+3|��	����r�%?�~.�������{���"є�����;D-+.b:�]��ڎ9��֥�j:�+����E]r(ʥǧoF.�$�U�^2�uL&�ue!�w-�<��Z[\�?u��#NӬպ���+}X�Q���L��Vٺk|�pu����ӧ�8/2O_YUa2�R�����g���R	b�%荛������O�K�~������UO���Õm�8�*7ꋺ��n�lϾ}~�
8�SB�劆��f�ʨ�E������(�!�	��.�T}�>�� ��(��Iq�.k��Q0�r��{�ɧſ'��'ĳP��.��3�G�.n��J�|$Mec=G���7#<�jlY�lk׬�|�"#P()''a3"ƚ���i�)H�%���SA�ɓ��-�����9y�H"LƇ�q��S�^����d��{�v�짏�w��4��$~��]����d�Д�Vة��}��mR��.8_s^�D�CC4�O?��}�_�3�ځ#�fXh���k'O���rҎ9��/'d�aW�q?Lu��>҃�L� ;�|�O�EfPϘ�'<ICY8#�#!,
���4K؍u��!o��n��Kn��V۹c�_
�ӱ�͎Nyh:�йF��m��H���P��R�Nyi[�j�O��>�)��%3��P���z���Z�д���}n'sq|���P�PU(�!
�'����EH��am*�'�Ā��߉�T&kSPj�HҋQ���1�,�",�A~�FoP>$o��3W�]�3L>���������PξxFJ��Rfؒ�Rá`(*��3儀C�B���d�3����C���Q�i�%�F�V��F��ì��FD�u�	�{�5{�>�[zO�Ke�({�D������=3�d��B�9�����%����/�v}c'�P�a�����������Y�$�{w�S��������̀� `8$8D�A�P�~�T�t�~���	^����
�P�����׾ږ���+w��ӧ��
Rݽ��g�;�Z+W�\i�p���vݦ�����V�;7��G8�;����O�a�CS9>JH9%�gܬfMX=L���?W�s�i�zRr�>���ԁ�����������.�9�s�:��/��B:�]%�Y:|8)nF���.m�ܩ���xmX��Xkු�I��g��3.�7�,@�j��Fp��#�gi6���"���z���F����c�W��_u6������z�swv�E�ߝu'���nl�;�R�v�v�ZJkhI^$8HЁ������y�ʾP�����/��K���;�z�M:�[5w�Գ�j3�[(���l��Ά�f���,7o�Sk�n�R�-x���jR|,4.Z�n���WA���e��� �貮�]��Z����,�ʯ�?�� F��u��V֏�������'����z7<p5��C�ӝ��E����5�ر㑧߫)�Ӓvᥲ5 jϦ��n>�޼���m;��tj��ID}���}���"��4��Ɍ[���.ڲ>ւ��&�fsd�7��{��|گ�.�_������w�'��)J
����ۢ�j�xI����ρP��92����Z��Y��##�{�ٴ�]����K忒R�o�M���6��f�'2 ���esp������}At!<���54���M��p�_\�`������_�C�~6��LE�Mdꆳ.�K_�R����O�~v���l�)�9���r����)����%�*m�]�=E�B��d�/,V����@`�<e���R�\1��\�<I�t��e��˗������(��������Aʏv�{3��q%\@�ğ@i�e���E�BK���q�򙏓�ޕ��ki�+�7�2�ߚ�J/�A�p�t�k�oeu:�$#��X|��}�������W�G/8G�NSe�S���u��`D�\9�xס�:�����nz��o�ׯ[[냶o�1���vz�c6%!���ܵ�F����3�"�w��[#	��gNs�v�z}ɚ����M�T���.1Z��8#J��Z�zL:�ft��L�F�,p:f��Ƕ���v�ti�m߾�)��5K��0�2�9�A���,0�VR�]����i};��;�\۴�m���^���N�D��<0���W��[�@�|L�^Puv���n���^:Uau��v�J�Zw�C��Ǫp$<��}�g�3`��L�[��>�9�<�|)��*��h���Ц��-����ऩ���hZ��ǯ�E๹�����*S��C���򵴛�G��"o梴���R�������z;�("�3��>����bkdj�G�#SC��/�I����q�M�-Z��	�@q��g��r�-�,��#�U�\�q�9K��(��o�(�~1}�˟��*�������k����6j�T�'�#%�`Y���{֔j#�0�a'-�!�Lh6+�f�)���Íә�0��@��#r%u��L�G˗�WJY�\ �:��k!^�����A�;� @�E�1c&LK���S�[W����F�0��r��A�q`E����⣌Ŕ~�q��~�q�r�ԅ�����^��J�i��X��'�~,^�MX,�c`� 0�ltB���V�� ̬�P������w�q��7��0���V}��h+`�n����Y�2��#J�6�W<�)bp\�3�p��p�����H?��(yL��/�+�� �z��5W�:�|�-Њ3�
q�^���NU�����A��m���k����gKI&�������Bȵi��Y�{���5_Oi �W�̚
@�cM�%�%G��'4�gZ�3�@����*o����}o���6F�*�ߨ�������j�9J�����ov�ޙ���k��� ��6eI�e: 
Q��fq㤧�GO�Y|���Y�ھ��������vͿ�	���p��N7��ߺ�Q}[{��ڽ4�e��}��Zs���z�pҼ�v��<>���g������bCF��)?��k���ܳf8�)0%��=�Jw&�E��/N�s�O���`6l��5�H�e��[;\<w1����5�/��%������M�췇���k͍����E��X�E����$�c�/�\�|�3�G���ȣ��v�CٹU����{J��=V
	�ꕫW��B)W���\��,�W�Keo�#�o�� �|	W2o�k��Ҳ8���A��"a2�O!��i<<�)ݯ�"CC�S�a�:<*o�_x�4������?��8ҡ�X�M��~hN�h�g,6�D	�^\I:�^�-�Y\<��"$�.l�����B�	�����<;0e�D	7y+ol��y�L����Y�#6���a}�%ao��P�����ϦS�/�la>a�S�'�
�\�}]�L8����P��{eA�	[W���8B3�e�+�Ҹ��X6w	S�]��7��BW�)�p��;�^��)����jq��ݳ���w�fF���ѣ��;Cth�}K+���uF��+s�0��X
���q7^(�R8�J>x�ҥ��_�ǿ����|8�����f�;{f���e�:J�r�)��7~څ6��WY`�𦣶l�l�	�����Og�Oڣ��rS��g���B�Ч��Q��<�]��j�y�Y��'�!��UGū���Uæ-�JS��dԻe�lS]7l��n���֬k�ܙ���Uԣ����z�a�֝U"JD˫��i��{t��=��C�>�9u�T�3408+y����и���K���6o�:l�fa����.ܚ��ީ�Z����u����v�?m����=ȹz�J�CK�&����]4Gb����wc�8���+S֔hO�Q���J+ᤏ_���Q
۪Us��>�N�AgOͭi��X,���0�t��>�o ���4�(P�2_%G�@3��R$s~T¶p>�N�Pf����� K)�[C��_~iر{Gl���.�C>vZW�O������W�3�����)�k�>N����a|���g�O�����g��Bv�7���2�{�Щ�� 2 ���Du�\8*|떭NN���3mCPg`BwM	rB�k$"X�m�e�7�e��^S=�@b�f��qW�!8Ъ}J��aD%L�M��P*j6Ct�/�L3��R7�(K������F�Q�]5�����Ƶ�ڼ[�Ig�?#�Ջbc��ȑc�GK3S�:���� ,��<w�(ΨH��~�q���Y-uӯ����и��E�+ǇO�:=�;!��mؽg��vn}:��Q���?Fa����s�"e鴓�3[���w�ە�Y��x���ܘ�r���F�ډ�@��s`�UJY~��H�Lܚ~ʏPb^�L��X�>���:���I��Ơ�B�\}S@�t��T_�z�R<��[Q���T�I�I�Y9hs7��x�R����9���(��IBU�Ĺ(b�$��[����t^[��Qf��r��͌x//7+,%È�HU�d�En�^:�<��2�.��#��4��|Pa{�����+��������]���Z�t��P��M��r����޽9�'���a�]��}5����\~����6;C�~�_SDt�x.(����୘K���,5m�iL��@��P��ס=/�����⷇\�RƵs��Ǣ̟���>�1x�`::%A?C�q<E�|����^��u`a
�e|�%;��-�eں�Ӯu��S�j_I�_KeJ�Ӏ�5��g=�k#�l�p���F$��kd��ڡ��� ?�{k���@_����oS��O<Q��!'^�ɥ�gUw�ݬ��q��(���V�&���Y�¡� �Օ�t-n��!�͹o����/~!�G\�������i�~�^1��ZZ����g*�"�0+��we�y{���r��1����4�~ԁ����Z������3+�2������1�5���Sg�F�Y�jm0A`v�~ǯ�kL\�ot�f�5
��*���A��]�Ո�ز����έ���-���oM�ܕ��ڵp�����6��T�
���-�m ���Dz��['�p�;��X^	�]�;!���q��UB�;� ПU������f�D}hSGgq�޽��]� )++�?�M,�S� ��w|U�y�e�0�a���-'\CK� ��Z���#N��%NōwKǃǅx^X|�Ph���`%`��lg/�.�M�"zU|#l
�(������&gXx�^d�vE^��$���)Fi�_�d�m�W�\N����i,�'A��l��Y��]�@\��
,l�
��f�3a�)�m�0�S�/�/�c�b��v��������qmY�:���[����㾰��P���w�r��-3͍�6���f
�j/�qcF�y�����լ����v��Ӷm;�͡?�-49`!|�,B��/��:�wp�}��o�����2��Y���u�[Pf�{�n�%����O~28��Dº�w�����uk�`�2dP�>�{�z��ɠ�P��={���-0�^� ��K|��w�I���/�ɝ����"�L]��_�Y9gC<|��r�ED�ޠ[#�A�i��`9�Z�0=NC�&B'�ն-��={w�Q��_8;�Z�bؗ�'�|�:~q:S�^��6@�e�FB�O9�ʌ�Z���yw��t��3E�h(�'�X6�	���ڵ���]m4!Y�Ԥ�3�i:û��H�Z�A�'�1o��p���;&�v?���wq=,��E������ho7�f q�v�ּ��{����	^�͵_ޥ�+���Z=ܸv'
M���k�捛��KG4"����Y��R�A�z��g���,�G(�jm�ؑtzu�a)�����(��Sj�nݖQ��Rd��v��7l޴e�u=����׶)`�z��	R���6i�o7�tۣ�;�ȴ(���{��W���<*F���o��ȿ@�=']�lSW�I��������8+d��n��ФY�l7
����Y�k�C90�V�ͭKfF����[G�݉�g�Y����T5~�>K�YXJ���$�lX�BSJ��sN��po��� ��"ZۿV�tt�oY���ٺeS�����_m���G�cQl���+� R#r/ϮU&�Ҽ.�����pq��gV�����ڸ�reɹǪ�����[������5�Q��x[��(s)��|�t|{��r$/�M��l9ƺ�����us�޷�����o΀fc��~l�P�֞��)Z�W�T��k�*U]ᯓ�d�j���:�^���7M��Ȥ(5�x�'�n��x���u�XJ��E!��XH��r�\qu���+��?�t��W������<|�w�R�\=�=5��VW~�M��By�&��(A�	t�t�	f�2f���aA%l�7�yF�+v��F[��+3�9_�v��5�ص�F�-��
�� �Ƶ�XB��h�F{S=����y��p�at���U��0�2��c�pq�UXc�������W�Ç?���B�7��`c� �
_����5�~�{��O'����w`�om ����[a��c`$�P���j�r�EsX坎aź���Odv1ќ޹9<���z1��VYn,Ԩ5h�A����|�~��Yp�X�6�)�#�R����ݿ�Q�
O�������8܋�eS��Du��Ӷ�`�ÖmQf�ƮOW/_�(>�F�&��+�q���_)��u�b��<�o�Qk����)�������υ��^Kǵ=�-��K�ǝ��OV�u�M�PF-&�@���{
�zhC���ѲNHP�d���۷�\h�#��:�^�C#mn�{���Qv��?K#���l�EN���6u�d@M��k�������ި/�M�Y���`�k�����O��p¢94m��R�!��P�-������<���U�N���̄��v�6}�����SÇ���mQ�9�1Y;G��Wk�X�����S��:yN�Sr8my1���Z6zr�_�d�� �އ�l����m�;�m�S�>�tm߷�O]�P(�^��y�-��}JE��-�,t֯����ܹk{x��#�o���B�XW�:��(�2��A\�A���k_�R�gD�!,��!B'f��0��O�B�Y@8�Bj~ݟsZ����4�|��'b+��,��#�Ǵ
�#a>���J�
�ѭ�qo��`��	��������:���)�{�� es��S�,��?��?�������r��\��R:%��L�{���.o�yx8w�Rp����]��m���n�H,vU�qd�Xw�L���bG�i��?���@��`Y{�/b�hM2)׽��51R�Rp�!h�N�Ҧ�L%8jގG��oۺ�:t��)�;�����v��*�e!0��9E-�N];.Z!�� ��V2sQlL����;;��	�K����n�4�5+:I���ߨ)�(ל��۔�����~M�$�{�.<͠�բs���)��a��v�ݒF��5���j�R\a7���ה�������8t�xZ�C���ž��59×�7u�c������%/(>���ɓ��	�=𨝹�"�<�[�����ʉ��.���t���(��P&J��ݻ������64��vm^g%�N�ڼ={�Ԛ:YY�}�ֽ�W~Z������A������L��+�@Y�I
��m�מMM���U{,��4�+�`�\Y_��}je�q�p���.�J֫V�'X.�I?~bx�w�n��� ����R o��gk�%+lY)�7��9�2��_���N�Yh��O4q{���� ���<�j*������X�_��6�$2еѨ����o��Z8�6p6�Ϊ�QDjY�;��:u���kŸ���$�jfն�ei��0�G	M�<�  �F�ue�7\�����C1	�M�h��1:��U�E3�Q�Ψ�E�J�3A	���⡌eΏ2`�{;τ���p� �:�����;���֙�SX��ټ��\���l��RC�)e��F�+�-�>������]�<̭MC_��6�IQ�� ���*P�Ҳ/��1��2�V��ᗸeӨ��ݕ�8�V��R�*���FfW����N m����x����:�BZ�R�,(1}�w'��Q�c���)r�x���P�}u��>���%S�2`�F����*�^�׵֗�Zk]R���:�"��:!"$����S�K��u�b�y�vP5C��1R��b�O��G�Q��Ι1�[�#[;lش���_��/L9Q`�i�p��sg��T��c T�Դ�đ���ŪC��jWp�b��ȇ5���u�8��}̦U�K�z65���7�]�ri�,(?�^�)s�7�)�>{a��>���d�s�~��;����t��9;O)2]�!�f]pU$I�.�J�)��`w�^��ԛ�f82�)0��ڔҨĤ�Κ�[�����Q�V�Y;�]��UÙ�g��GOV{75ê��	�|�k��uG�ח��.8љ_/q��� W��ǫ*��O�3������ʽ�����d�dk�6S�첤\����Ñ#Gj �oOd�u��fA�(�M6.���vi<��2�G����?��8��>�z���a���e	��%�*g���4_����;�����c��a�C�y��Cm�v��:Kù�ϝA
����o_�}������31^�x�� ��,#y�o��ٳ�3J?_�cPntx����σ@��>	�?>ϔ6�`�ڈ4?�!�e���bQN��̶g���nS��^��E��z��@I�UE�׾p<6��5�R��Nj�IB��Q��w��k�d3�ſ���Z�l��q��p�ٙG�p岝#��:�{i�����o蠣�9w�(�'�B��m���$��h�w��	�R����Χ�43 ��N(��+���7�:�8��N��(�Q(5u���6m�ȱ:�1�i��Ų�x?�
n�{���[<���%n�!ؼ�rd.�YbG�'/צ�H��/y�-kJ4B�%к�\�ͭ%��Ȓ�Q���)U�L٣P��\�N�\�s��AW�,�~�����׎��y��[�LgС���=���ˆ%��Ϻ���H�;:��2Q̜�*�:kSJ�a]	�m��UU_��V~����-��e�c�z�ͷ��'N��F�AWj�hq�y�, ����k���`��.��yғf��8��$6�'z��2
�*�t�E��������Q��t��]��^���L���S{�����c��}�������
o���$:w^�u�t�u�����A�]���J!۹{O����X���t�����w�λ�tSlZ>�5�rx�d��_��~��ڍ������
�M�������֗�貍 *@տ��݆q�r�~�ޗ`v��o;7����.z蠡��tm�C# (vd-�
����i��p�|�#�i���^�f��;-�N�����?S�9�۷}����k����w���x}؟����_����Z����W|u�e�Y��㓠��ʜ�J��FI�rBi�W#��0���ںX��sRj������f����;�?����Ås�S���.�fK���1rL-�B�Y7�eQ�K��E�%���*<T^���t�^W�jgF��k���g/�Ԛ���^�^��v��"�|�>��'l�]�Z�0|K��L�!��P����]ф���t��Ki�i��Y@�� �#�}
�=���F�_� �ꌨK�[���� �^��kK���v�l�PJj�f���7��l���t��8V�F\���KC�s?��Z��/���]%�;;�(4x�f�?E���E�+
kRme�Μ����[�(�Ui��:�vNV�j�Z�B
��I��>��?Sn��*��F�Y��+���4(��S��Q���+�H���BL
�]1�9��ڭ�C7�2�q.3SQ�<yI)Gk�.]���p8�M>�ي�� �+8~��[T���jt�K�ES��֑�u���E��=�G�7����X�~�Lۋ�u�f:gkhRf�5k�|E���?|8m��@��cT�U�R;e����~Z���vvp8��Q�Ű����x�w`/�T��ChNv�U~��C�NڥE���/~��aמ�ë��|x���R޴�D)��\����N�sWG;�;=����5��n[�n.k��G�ޭR�)�1�:�^/�c{'qܬ�Kn�Dډ4؟?d�i��rD�@�td:��El�9M�F�+˚r�ԙ���� %ffS/��Y@>4Le$,�S| �6��Qbl�3
�4�+��Ō� �� �^��@��a)�/����Q<���5��o�����C���o?�����Qn�V��:p0��#B���x#x;����݆0���\�N�
ׄL�	zٔ�(߇���ѵ�0�QX���/�Fm�+��T+��(`M8�T��0\�zk�p�rF7W"�,��9<�̳��vv��>J�R'F-ǂ������=�\5p�Δ�0�[JV�A�9{�L)?�Ѡ��,��ྻ���$�o73a)�ڂN�{#T�jF�a���B�7o]n�mǸ[���O�<�~���E�7�����$���4\7شD3�<�i��):`�YD�M{]aG�uPb��qL;o*��Ϛ�@u(�?�c�]�߸6ܮ�t	���	h�#^�)�MNҶ�� �T��S���*V���W�
=�|���(�����a���0K�~]>�֦������=�J�����>�T�[o�U����8!�+_�Jh��0a/^�\�g�?Y����v��v���w�d����y��"Q
I������_���^8����&���ʛ�;�R��	�ء��O՛�ǵ���pZZ|SS+�QNO�<S�aL/��������\}�՟�6������T�9��>bPG�����N���h��r0K�Y�Ǫ��{)]A�[�7��,ƪZ�t��W�L}Ѕ��erp����S�O����j
��M������1��&���j6k�~�����O��WJ���z[��CM˧��2>�;�s���$m��Vw�N{};��`>�#���_K	���{�W�j֚�=DA�E�ՐGv���G����՚e�����5>�~�6�q�	����r9��t��@�3�^�|!Lq;#�U�+�#a_-V���wf��_
���3E��8P��QD��i�F�:0�*�A����%k%��c���6��w�X��E���/;#�Μ�4���;Ç�O��qD���`��Vm�t@[�K7�&uI�,a?ϭ�Y'৅iN~��pѭ=m�tZ\o�1/`�KҶ}4�Ȁ��A����1;5�LFq'���(4�d��T�m�p)4'�i��(|�|�_�yeJ>�s��8�q��, ��������e���y?�{?p��r��KL�nٲ���F�UG��¥�^�O|���Xr�J#t�a[��]G�߹7��ue5�<���qZ�k�]ۤ�	�oH	����aEḩ�%��w�p����T���B��W(9����k�c�Z�D����F�G,�$kLYrR���2?�����Ah_�nE)���n�;���/�N�E��qI�vשo�'eQ�� ��J�D��˯��z)6���Pu9~��M�Ne 胟����;�������ëV�� �������1:|)ھ�9'��6[��&�߯+��\��6�RC1!�M������O �̬K�����Ԕ�ѣ'��B������WoD�9��Bf�%b�ٹsW������A�	�;�������>��<������$�M��y�z��d���ݸq5�c�Xoݶex��'�wm��O2�������}�h0g*6��釾������^����-+�)(��ᅓ��������B�e�~����>E9����%˕�mK7 �4����J�<P����@�*��(@��k	�f��J��	�����6_����^��a�s��Q�lyf�N�w"��G���ڿoa�/����ٲ�0瞏�Cɩ�R�� >z~gq�X�w���є�P����I~F�4l�,k��O���5��g]`�f��yQ�|��i�/���(E{�p���A���an#[
J?94���4�����2Ç{���)^�3W#�м;ku����]�/�:�Wޔ��)��(2w����F��Ξ�Pe>����C/Չ������K�q[[+u�����W+$�?���?OzmJ���)@'��|��2����i4KǢK����q���'Aϣ��r)+�P�k 5�ܱ�,	�:�����ʢ��>s�򴓐⧞�~(U�v��p9�U�Bâr;m�b��M~u�1�dTfD\���/�v:o��r"a~e\����;�_®Jr��IXJ˚9;��z�:� �q����'�����Ř^ܲ٧�|�b)6p�T�lؔ��{p���v�p5J����,;�����,|���t�x�;��w�o|���Z1����=�r$_@VR����@ڹsw�58t��{��ЙR�W(�(?c�_q�=�淢�.v5 �;�wV�"��1�c���H\k�\�WdI��5�Ĺ��t|`�����+��Ƃ`��<�q�@�̙ӵMݗ�k}`��w��À^]��H~�{q
��N����@�]�����-�qg�W���v��0~v ڙy�ؑ>��ڕ:��)���G�_���?~��5i4�%܎��_c���0��_�"��C��ܽ���R�M3[�f�X�B�ec���N�M�Yt�-�o2�����U2 .�j�����h���y��� �b�p.̝�
�0�iQ��n���& �o�092�z� ��X,j��Rd����ogB�f�lʍm���{׮
o�ф5TyrŔ3��ϳn)�F����hʬ��iQh�mh� �d��P������	K�3v�`|����c��s�^v�����|x<�TGF���8#�ꋼ>�a�8��4/hw�7�׮�p�kxp�.o����N�l��1|\cQ�4xu̪�'��[F�yw�r{wp,���m�����/���aw������B�z�å��Z�կ~uؽw��VF��s9<��e�E�]9h� �����t�`�����A��BK�gA�=a�-ݫ'�hi��K�P�w����e�(�];��<dT=��:�ˇ-O��\81JF�$��Ԭ�k:���ť�a�æ�Hg8c���Pjnw�,.��E!i$L��/-q���mҺ�2�k����	g<l���&�]6%�R�3�v��(o�6�.\��+����^Z�/���w�ְ�ȫ����>t�q����V�p������iN:&t.+R�i�xQ���Sn<?��С�JA�����-�ᩓg"��'C�lݞ���Ȱ��S����a�֮�"�2��B)ɵj+4�nte��c���	���u����!qx_�+��Vr��k�/,�B۫5}(=ef���]�~m�e�����
����Cw۷Z��������ں�i���g�4�nD�������/u���ޝT��1K'X)��QR>|������L�rv����G���(9�T]���ǵ]�' |��4m��x������q�� ]����]D����t����o��-n����ê�w`����,!in1�!fd%�x-�}b��Z�q���R�󏥡v���:J�[�������k5J1?i�8�	(8��tv:1SXm���CxǢ��>u" ��Q�����ֱ�Y1��yR�Q��#�.�_� {��"W����(3�m�Cȳi�CR`��	@�5*�た�,��'h(p a�3���fL������#QZ�P�p�+�!R2��^�Y��׼[�f�X�T�V������+y�p����jSd��3ws6Y��������g>[+�-&}��w��c�W_�VϿ���?|���w�^y�'u
��~���Ʃ�k�xS�W�9���%��&��o��� =�"�^�5�@!�# l�􀼕�_�B����u��_z1ى����?��sy����ݛ�յ��U�α[���(;�|����G#TM9�J�CikjP[�E`aԿ('�=��OY�;�q�+L��\��z%F�#E��oٹsX��J�+��F����2��K�z�v^ɦȂJ��0.�#ș���؟�<�\����t��Ͻ�¼�S�����^��s�'���� �a�_�Q�a�Fc�����+(����I�˗�H������.��BgN�9[��m7o�P��%��sg�Qo��a�*�<��Q	�6�5k��Ȁ�"N9�M��jߔ��v^����y�n�a�ŷM��)?�3��w�X�(�CY��"���޽g~��_�3�v�h[�C�;�� ��3�٨=�j��Teʈ+M�5|/��F�Vv��u~�Nh#HC[A����}zz�����3Ed��3e�AE���!da�CW��}Ǚ8[�B��;v"��DrMe��+eƀ����������ɀ���w����5Í(�v,͖kiz6r�YI��3��"Ň��5��6��֯qؘ��ٻصk_Ҡ�>�jxhJ �TD�r#I�"$ fc.�h�Qjv��YV�Z�>��� �>x䪳�~Ҧ�b�X�/�:&��kW/��`=�΢������Wk.�b:�;IO��ճ�Oo`�8JM����b���s��k�S�!��_�S��[�5����ʤ<񜑀�vm�_�Pa)��I.)���u�)E^�	��=z�.^>����ۋ&�
s����q��D�m۾u��ѝ0`u�ke-��]�n,�C�(>姊�ntx�ҭu����5����c�ﱂ��C��(2�n���ZhC}�ʧ!�<o޸]k'>���j����u�:ި�%��:��Qh��􏆧� k�?��ca��3�y�}���V���N�sPt
�sm���#	�G��Yo��S@�Y<��$�(���7�~��<�������cÁtl�a}��sθ�g�y:J����ַk]֗��á�/A)i�Iۙ[��5&��IOC����:�e�Z(�%3]^� ��PNǄ',<e}��0R?4m�d��a$L5v����l���Sd���wnQd2�_�jؼað+��v�-����oJ��(v�F�G>|/B�ʰi�������-Eeu�'<Y��>�ܡ:EYy�C�{�WJv\DWj m}f�tA����:4Ru�������?|�3����֋�鈴u��(@����uf��n۾����j:%|"�"�����p �
�;`�LE��/u�(z�3�C�R^(*����tYg���������]�@�I:x���
!�o��i@��ڵ��5��c?b0��������Dm��3�/~��(�	����{ʭK!,�������?
���¿*Ce]н@ShZ��+��S��]BU������I��;ѹ5���3�=�2 w��ƴ�;��n����Ȭ��UÖM��M�^ݯ�].DXO�a�أ�y�"ΤB��X�I�V�A�ܴ�5�J�i0�7�;{��`��{���&���������ܳ/�۟2<FJM�����n�a3mt����|��j�%|�E�I�պ�=4f��yd8W�߼M��xP�d���0���k׮J#��u?��+�bPT�[f���i��o�����#��_Ψ�H}�lm:��w��;��N	g�$a�D[��qU��W��P�h_3N�s�Hw���%�{��R�`
/̓Τ���!PGR�]MD@H~����('�I��6�szn�0�����!��F�ss�K��\ܾ���H�����5f�h�$К�H`)T{��~	2��52�ݻ�8�"s�U�4Z�;�+l��0lX�1��\���)ﵔkM}ۥ�Oy),��"�o�����cU-��f���O��?�á�%��W_N�<Ys�?��kDGQl�}o���J�,h�aú���|�/[��:�V{WPޟ�	]�0�QIػe���Z�X��{5���('�v�_Cϓ�����Bu��Ŕ7�����ۯ�=�V[9M�Rtt��z���߼ið3�����F���D:�Q����kx���S�>;�2�w�<=x���ߗ�}���cݛ�O�~Ͼ\��홧��d�&���v��;�r���}�^ѡ��	�w��9d�˳U����#Tw��:cS-�~�$��>�`ݘ��={*��b��	#�}��F ����}{�ܬ���w}�g�r:�_��g�/^�y�j�ՠl�M��P���4���I��RN�����$�s�3X��Z�,H,�:


م�Z����,����>�?��|��]��4�.3)�v�=�����m�e�2���,A�(^���z��5)K�K������,<kKq��.%�UE���~�ŷ��Nj����1E�q�t̛J��yh���?�����;���n};U���֯}�Á�O����g?���,Tg#�z��D�WS�����챁��i#
�<��*]5l��'PSb���,t�����p�'M�)�t�J6�N�ἦ�εa}x�^��>���~'�Ά����[Ke�Ϝ\�5q駂�)슣�ʌ��@d,I�͗�1�;t(JM��v�칢�����w��[�/��Ұq��a������դ��x���CSjz\1+�ņE�~A��o�F�r����;w4���#em̲��b~�kJ�7�K���|��$72��]#6&5�0K�>|���o�n�wc�1�9�(b1���E��8~b8s�le�P'���W-D&�L�(B�<�E1�rT�8v>U>��+��4j�<:�y(P��0�K�~U���(!�fX��\��ZzM81����2����w��:
́��,ä����#$�Y%6o�8l����q�w:sDǮd��`m�{[�k�(yީ)9�c��lF�s�h��#c!���癞Z��D�р)LF~,Dk��4ˌ9v��-��g��Ѹ��#bv��۴b���y�,l���w~�o/��bFGk��ƛ�o�}xp��Q߅��R[x�A�$�mW��� ���F�6�Ut)��$�Ӹo����9�]���]k!i:<m���������ﭚj���5���/|n��G�ɟK'q�ڇQ��>:�>9g�J�Q��8'��buH�c���G�ұ���~p�9Le��p�8�28Y�z��4W�F+�}���J��"���UQ��XZ�Ei􍦭[��ȁ�e��3|��/�Z
���o�:l�nK���:0;<���1ϻ���ӬK;[r����z��&��򵴇Q޷OF�b�y��O��P6�xC�KN��ꫵ��9E���SGP$	�f�Y�	W�ˏ%�[\�9S#�L�|���b!��Ӏv�Yc*�B�����>8�7��4��Pr�JF���p'��ի#_�We�vP�]q��u���Rg��o����)Y��}�P�\+|�~��t_=�I i�Ո�2�O��f���K�+�)#�7C۞�v��wֱ/<�bYi)>����>�Wɝ�²C��~-ʙe�Nx�i�t*W�{��;�9e,�^#>��0~ ��d�RK��-���_�0s/�����������hk<oܴ�8ϡ���T�O~�J}����Og�9}l�^���r����`� �����%���(�$L�/~V��'��lu�����l�O;"3�g�蓗���,+����K�K��\�lS��{«,5�+���RTD������ah��?��3,��u��ĭu�ԠfS�]E�Y`yԺ��[!���h�:�M#L������pKG�5���;gNgO���;7�M�A�NyMF6���Ť���q���!pmWD(2�)�a�+W��0̎������(�)bǹ�}@&��4x�~Bg��[����(�ZX���	JP&�[�m��VK�خ�o�Ҩ�����5re�p�&kن(�" ���,����(JMa+v�ێ�ZP�+C�u��<�˟Ғr�)q��'��F~F��H��ָf�9�!�(�8#Q�V'[� �K�!�-���؎���i��^������^��$�w����w�މÇ�NO�am,i:��3m%��s�}���4Qڼ?e�3^�B�@	?��e\�`��s�]�/xkaZ�x�F�h��������/As&���\|I!��kK��o\�fʮ�;����>��ۉ����(qG�)�vֱ�Ǉ�^?<��Z�k����(������HGϟ��==a9q|8r��p�B�Z�%�'O��$|x�h��N\8?����l�?�����9�Ʃ\�^�<��H�B�L�ܾ�6�(��ՋӾ/]-y���o��{���p�!l��x�b�%�ڕt>�x'�oUw�ʍ�֍;%kv�t$����:hD� ���v͙��g]��F�]G�ͻ�w��1��?� �ď+:�/Wy�� \ܪ(���@;w�j��G��l��� �gBtx�� ����Y_䞕����na&�]Ia���X���,9)��8ڀv�:�攳�/�꛰�J�`����e��J�oԱ�[g�b��A���Od`���'���ڰw�����KÛ��1����j=��t����p:�g�i-
[�5�Ay��(�}S�Яh㿺��9ƴ�k�l�_���6>�\�B��ߔش���x�f���4FT�`R۴V�!�_��W��� O[�9%��p,xi[�)<�����[(Ӣ:�O�r#�y�كi/;����޹}sع}��;��5����v����yN6��>�v�$�J�Mb4s��E'�o����O��Vj�Կ���{��G?�q���Xo�@4��窣�|ϣ�;�a���JV�OܾmطgO)4{v����/�����Zkq��|������4��3q[�~*���'\0���e�ب���;i��3�qѡ���W�'�ڛQߺڥ�<�5�ծ�U�����u��x+�H9�#�P,t��&��׮k��^�;�HCNCX�?{��СgK)x��������AV��b�`:G�����8�m�g�Y���]8���c�NMS���)�5FJh��[�+=��RВn�MJ:�>rZ/`�SYD�԰4�eL�������E��pܔ�����A����|��m��ُV���[�/ev�`��j��#��a)��?�	[�P�DxSںV��h8V�Ӏ�E�F{B~1(#~�x\�RO�N>�W���u �Ӱ���������V�J�#Z�"�U<�DRvElHs��R���Z�&�o/Q�JPn�ã�5�u"���W�<�9�*�RH��L?�2����6���+QCxj�4|�+���	�0>�ϞtZ��;4�ؽ+�t|7jz���(DQ�l�Efm�b�x�ީŏ��t!�r�6�^�eTiM�o��׆��������������/����տ���i�J9��{��bhku�gԽ���*e�H�ǳ˿���&9���`��E�Y��ݦm[�l*ɉٿ�;�S�)�_�2��kYi�ik�ı ��c@���X2S��ʖ�YSW�I�Lma�ܪ�S꛸Mv%\�&�F����W��@1�y��|�A.�+K�O��O>�?��n�p��ٲ����kE'J�{�W3�2���U����aA�+>�k}KdV�0(�T@�#����6��i��ࣴ0��N�5���c�pJq �,��:%|����O=��p6xr������/�"}�[e�g���_K9uV~��eЩ��e����L�(|�o+������������+�����揾5|�k���m����/��B�mS�j}ǣ�Gb��,����A�B��WQ���[҈L]nX�̤�pG9Ԉ�gt�|a�"4A�������j�}ꩃ�/l�;��p�ȉ��2�;��#ǏgΜ�g�"���,�U#����#�OɜU��h�[`DᅪxU� :�V��Gv7�^��L�U�
_^q-�� ���5��3�U�<��	r6j��W��Yp��1���W��0��uO:�m�1�^��Y0��X�m���������,��TN����B�h�tհ6�Թxs�7"���K�k�i~���*�$&b��К4DS v����W��.�Lv���jt���cs��7�����/�\Ӛ��W�WQ���6B3q)�+2b#����֎��\�nmў��vnL���M�+m$"~(GU�L��[]���MZ����ot�+z��w>��������7~����(�^^~���ב�k#�gӂ�=��H�z_��ZS�ɧ¤��vϨ����%����W��r�o޹?܈����y6��*�:�k�p+��ݛi�s�zT��=�	����kk�n��ע��H�<ߵ�;�P����J��Q���[��o�5���ÛoN�|�,RW�>e�i�!mC�����s$��'��N���0���������a�ڀ#JwxUgh����*��F/;=�Y��:���}0B��`����-@;����[�A\Y
R�\Q�C���k�/�~������6h�P�
K����`PX)��;�aY�G����:��nr(���&�Q>��\���_�O�jRT�d��g���d*kq,��5+Elǎ]5Hq������_�3Y����?��p8
�݋����Ϭ��-�iO�1Ue
ߪ�0%S�65�9�&\�W�nuw�7��>zh}I��T2����b�����y)
�i'�fmkg���.K���S�RH$�:�{x�:�4�?���P��3X�&Ѡ���gҧ����nf �fx�٧�g�X�7m���+�ē�/����R�F�kd@��ж����x��?��2�������j��'��2|���/���M�����@s^�#P�b��y����"�Xd�w��F�:�"*�]�_%TyVǒ���q��(MʪI�檾U�<Ju�8�rl�X�;���L �����Ic̺�B��������j�pI��԰�n-
�J��;BȮgS<�������~�k_��Ѿ�b���k�G>��u�)���޽{j��_���S�m,8���\ݛ��F@h��Rb��)aC��^E��ު.����b��/���0�4���0�e4YgX��_�ɧ������W������Ŀ;���A��:-Sh�P���t�;t��mj��/�+m�V;�w�wRߎLXtD[ #�&j�|���XunJ�t;�Y�}Ŷ8ݍ<�V�.���eUy��6��������ߎ��F��,lݾc����f�@	%��m�퐲U�;̨��OTG�����ҥ�Z{f�i���uF�9�+��E�[�A~���a.4b��)���iy訌,7mp���R(a�M�J�5�����cⷤ�5�q.��M[6M;�7oۚQ��t��jjoZ����w�'�����Ճ�b:3���6ż6�}�gS�:�]�/�7�o�����5>Ӿ�'�/!��?�������N����e�t��̍���W�"�*:!�?;��v)�i�q��P���_�-"�ܧ��q�vڅtR�x��|�g�ߓz>w虚.�V��[����7�7C��G��5�Ѧझ�죙�S3���ǵ�}T�5�u��3��WN�^82�ֽ�����x����:�{�L5�QV��f]����d���r�}�C{g����G�WyR��
�sYq�Ӕ���NBL�� Q
��e~��t:=ի�si8@ks��@���
�ߘ�y���h��x�W�y�Fjɓ�CFp���>	��6��}�����7F��RR�k�$xga�dnr�POi�gjk����$}�_^~��᯿��፷�	>,q�4�߽i������Zʷv8�t���-�ܜ��>dx(JMI�1f�g�h�����O��Ok*�������>}px姯���Ґ��֊�0_Q_I�:��F��w%�c�5�ۚ�C׊��W��j-B'��� � e�)OYK���Vyc�\J@�2ɢ����{�o=�D��{?�qFΛLx���)�*���25����e��p�"����hȔ��^U��A�ҵ`TJ?�-!2�z���_�������*���1���N�Μ:]�D	 t����55e��>���w^O��	���@n?��
��)y�c�6hWN;���W�E���픣-x�5�Og֮� ����]�=�gI-#�׆���w���U�)���9{�, �'��ڍ�jd�(:�N�"���5�+"X����c�r*�W+�@�����m�4y��m�(�_�s��|�[���e�U�r�&܌x��9���?�/��_OV�5�$֮[?�J}-(T/#�Z?
�}�}k$��'�������FCs;�.���@&��#G��ic��%����	��Q�ڹt����5�HidcTS'��];�L��/�>.��O�Y�(���<�c��8�SFN�7����%nmF�er�_�w��Γ�d�r��2M!�e���;�Q�_��R�����*�=Z�@�оh��OY�����G<$�6�w%�tDi�-p�¡�8������]1·�^�J��*�Ƴ,�+�l�����+��znx��/�>�lF؛S�v��A�y͊�JB�3�R8(p�WȌ6����N���&�|��k����ѱ���R���M6������Ȓ9�3
�/��._��:�ja0�Ʒ�2	��68���3Nc��0�@��UZ�us�	����w�uѺ u���ss�u\#e[��{)�dJ>V̄	�C��c�iJz7�ޔmm��5�IƇ��8�ɒ��i4��k�Uz�1�РY�◲VZU�ֿ�)K��G��d�V~�_^J��ӯ�~��{��������������'������g��Bʰ!�r�8��+5@��(��R��o�ټ��������S�~�ӟ������B)AB�#�`�_�S^E��/�;+)F!�k�T�1+����Đ2rL5a�A+0�a��*�A!���Ő�bu�Pݹ�~�嗒Њ�����8�Y��:�7�zÐ+�k*��|a˔b���/ה߈�@$�0��i�y�,���r�ܨM�������hg���������7�C��ј��:z��Qg�P&����u.v���qæ�&^�'�|��Ou���	ܔi.�_eOsQ�j�^"*[�$���r�Q$L#�v��&�L�A*'+ A��|��s�s������p9�v,�/��_o��F��)x�}����Gஊ�V�RSue�ߔ�)�Ռ,Yr|ӈz��v5���׍H���5��Ǻ�7	���[Ӏ�5k�&e����-=Q�����[~I#x��8����?�������q;DZ}��)%š�h���SF���ҬN*���_�qړ�Y�To9 �$����w��M�(CY@,.O8�/V��jˉɟ�e��?t)��4L[�$+��,;����T	���K����6�[m�V�%O�W�,F��j+w�S������:���/��g�Q�6N��Wr?i�vX������x�]��W���K
����/�+d��k�v�L*���$�t(5+�A�wڔ��u��8§A���;�'�$8e���_����������S�(���m�pt�ʵ��>�h���|��nA�4�5ڠ�T�����Ǎ�QvC[��n,<֖�G���Q����z��*c=���~�Ծ�+t���._�\�0�%�U��[x�RT���K�u�e��w��0�ʿ^�_�\j�z�^t��E�Q��g�.�� �τ��/�ł$G�8�(� IYh�)5E���p��H���"*����Hzi���+��(���ܧ\�Ü*\�4�Jq�J'Nx��6��-]Pu��2r���ۿ�[�~�#�}�)X[S�s���������0�����`��>}aa{����*5���R�Qh�0����7�x=��?��o}s؟�ҏ^�����pشms�0V���3h��m�0�L�)��,Fۨ#�{�	�����Ij�D�Ha�ОY�r]�au[�����&���*j�XL�:�w���Վ�����p)��͔��Q�O�jL���ΔK�����R�!i��Z��{#q·��FYTR-����,���?���o��u-�h:7�.�e����	;4e6�z��u@֦M�u��u����U���C�um�\C����haW�c��z(�,hd�1�c5�'%�N�~��8B�����/��vD�>�i�6�h�Z�
��U�:�#�йWGa��F��e�ԥ#E�ɹʚ��aQjl�n��֑7���J'ޔ�M@ɛC�:$��5Յ��;	�S�[�����W���n��w�����}�k����������A���:5#�vƑt��(�?e�_-�M���0%�2�u� L'�������a��S��;�!-� xG���]
M�au���i���vV����\����TG���ڦ+�����)I��8_"6�*�RL�t��� ��t���S���,�q���yd��ox?��1i��)���@����yp���U��t�B���E�)�z(��إ�:<�t)x��*z�A�����w�#�:���E��:KފVv+�ڳk���3��}�Ղbm�ud�����x=@��i;5�6�ꥳ/Z&�6f���PLXK^џ��솶xPY��ѦYb�UF|S�s�q�J�o޺1\�|a8m����D���6x��	��.�/Z'pJ|o�D�O�7��ik���Qp�W�#K���
ӡ�&j>�@vM�OfP���M�:��S�G|���������v�2��H�)�y�����������r���g�҇���3��Wߦ�Ie�n�/K��0��t��r����iiG������(K�s�ф';�{��sϮუ'j�K畋�k�����$��a�S�|)���HB� �R��b�����o��/�e-���oG��u�W_}m8r���aӖ�V�q��b��k$q�j�f$�ib#`jˈ�j�b�D,С{m�0���DA�kG�(�I&	|Sk��"1�F��(�٬O��w��t �k-�шN#\�:�6o�:����ႏ�Ek��Q��ac*����͈��V�d�H�����Å�ư.�mJMb^w�$��)��:=4� ��i�K��א��H�㜠O՚��|�;ót�2�csۯ	`�i'r:���h�v�iX�9�l㦍������[�!YV�s��esJ�K��il����%����u�	��tvE�U�Z_�6�3JԉK�t��Z��ԩ��;o�5��{�-k�O(ԗ}�c7��)5ZS\���c}:N�)�D���<���ڢ�����z��ű��H�C
?x�6�9����[)'��%���J���Ô�J0���)�R�(�V�꣎I8�*��2�.��h�L�mǶ�wM����t��W�����ʈGk����m�Fp�7�[��O���CG�v�h$v`��`(h�W(hmJ�"v����]����m�x9x��G
�5,(aY�;eÿ�S��}�E�m��hC	زy�p���j:AilOgE9-	��ʃ���������e��K��]p,���zEYI���W�
!�ɴ�:�r�W����	��v�N�ͲX��)��0���z�GP�:߾�FW8�q�gW�MR<�繬��v����c�ڕ�J.Kk��=���[|BY��R�eS�`�K���ww���M�ŋC�@qwB����šP,�P��C
���3�#v�~8sg��3w�z�H�����`齗Fč�6�`m��iV G�];��i~V3��:�ܚ�Kc
�}��?��VNgd��ü��������n�	�4j��wxtf���� �{�L��<���꿛�/��E��j=6��.g�u"�v*�����_���;$���1�\S� u�K���U���<{��k����l�CĘ�GN�:B�~ZL9	�����o�����\�g�D���!|�jT.S�ÕV<��+OT�h�盻���7����J���l��g2���7G��?�%6z]��$hC&�`mn6��2W��}/��鵣�m���ݞ}>{y����8��d�%��Jus�i�� ��X�ײ�>�E^��
n]Q��Hl?���3�ΚI��og�"`������?{wUUl��-J�;"9����Z�ws��e��=��a9a�� �F����^�������8��G��n��9H�m��k>t,�����LU�O`9'�J������A���a����c�F����3ǭ�����.���@QN,&�p�ZL�k���������X�S��/�_Xe�B�B���n���[A^�����N�cQZ�YT&ܨr��7�]'ă���o�����qգ�B��Z�� ؚ����-my�1��
�K�y�����!����A6jab�gQw��eL�$��P��岅<۔m��ױ�z6�N3J�qs���M�0ԋ:�:��r�6���'�:*'#�.��O�>��C�J�6��]!A@�>t���H��JE?_�8S�N28�U���<�w���P禎$�	�U
��(%O$	�WV�y�fC)<�ឯ�E6�V���,h 6F�~;�4�?�����̼�I���ݛ�a��A*�B���64�G�_�[b�o�����ką�9�d$qRd��456ݺ�
��i�D��f�b����s��:��Q�2\Q}!��3�f��{�C����i�f�<���U��/"F\� �`!�u��#C�1{�u3TOP�!$Y�Ʉ��v�F�c{\R�hP)��+��.�kѼ��K~ L/�P�������s�
-"C��hbS���S�yf����)�d����e@����浓|FCT 9��l�������7�]�a�˜��P
^P7��Z�&�n��H�Oa���T����[��b����l��H���q�ep�vۛ��n�RY&r�G+)���GZ;Xr q�{����F^�T�{�A5��ʌ�z�f�(�m2�6!w�ؽka̡�Z,5�a�7Kl��J�J�6&�|�n��O�k ��·��Dp,��Տ�����zq�6X��hG�Ȫ�n۞�������u�& E ���T�<C���`��y����/7��ݍ|~��.��z��C@w�!)��i����*|��w�b��&��h]%
����3
� �߁D���(#��]{�Ld(Q8�4�yj��".������/���]m
�����ߵ�5:AưI���F�We�D��e
�"�qv�~�8�YQ�8zM����?i��
4�vU���}ÍI[E�b̴LO-����3Y��&��.taS��Us����Oώ�����F���$���U3S�\ɠ�fT�-7�~TPS����f@/��7�K,M�&��c�����FTt�<��o��n�w=
qv'QD�CPD��4��vm����/
�k��u1IvL\}���a�D�G�&�5F���ta��r�� aoo�}4-����*
�w0�1UZ��,w�5�$�Re��9`�U��� K�UL�ܝ!!ڧ����J�����8���:��I�s���/׀�˛	��p��Zg��G;<~Ы���6qw����f�24p:B7��m�@�m��h��b��m�kI��Q�'����W��?���Ӑ��>:'��Q_��dZ�|߽,���@�0{�Q�eX�h�ͫ�oD���4F������:
z��|q��As+)l�2�uu���i���H%���y��)��Ͼ*~{� pَя+Q���Y�������X���F�T�o���Z����+!	q��07�Ւ��O~76�Tf9��tf&>ci�����E��<Rа�м��4K��>�^w�4����fgB�P�ui����� ���癙�%s�O�7�a�r=�	&�*�q���a�{���}0���&��Q�"�Is1=���ǥ?'�kP4ߚ�*if��|�,^���3�|� 
bƐ�ր4S��t�:w�t��Yo�m�~цZ4?����A:л/χ�鳯��ds��O��h�F��e�6��-kG�h�K���B~Q��J���Q)��r�� ����T��$˭��s� �nY����s���ޱC��^�l"�����!�앰Oc�T0���KQ��W55ѿ�g:�)�~�7g�؃'���ٖS��q����#W�	��ԋP�(ߩ��X9�V����_E�ҳ���$q�R|$ga��`�Օ~d'�R��VM���b4v�T(��3F�&k��mr�cE�ܹ5M����q/b�:�B�2�]B�_u�f�;����r�ˀR��d��oӠ��x�k��� �ṮI�i�GLds?�K��y�(���S��4�U��x�*�*'F��@)�R��9o0W�B�Վ_��~���3����G���p<�ͯ�4�ǟ٘Ȱ![[��C��b;�Wfa{Z�eA=;��6�'��-��=H����{*��ej�nP�/�=3����!��8K�Ȳ2M�����!V[%������|5��>����':}&O�Х�#�Y���[���h�N6+���6e�Wk'*����Jھ0!-�!2�]���H�R��Z��[��>I��8ʆW�����=�>(�m�0҆>�v��&��]�>?��t��J��(�3I���"տ�Zqj�18�1�ڮy�2YT�=�a�Z>ŗљ�$��RT���HT�D�R)䆰PT�t�$^�](� h�r�����2B&fTg���$ly�([;���.g�wF-;���H&�t��&���kF>���
�Ju\�O�,xċg�x�����\����۵��S1��O)Ι]��Bl�m���}#>wҤ+��)e���랬���IQ�o1b���!5p�P��Cب�z�a�@���<�ME��M.�����W�J�=����l�B?ׇK1:%�����osQ.�+r�>�F}�N��0 |S)h@N\�`��m�M�Q����޷j��/���n�6J6�/�m��r��eR��(�v���2DюU�q�Ӹ=K3�"���۠#}�5?_�)W�#�k���	Aa�l@�q��t"s�R��0�P*�V<r�S)ܨN��t �q�����l
���~�Xl�p�ьwQ����� �w����J��Je����i���W��5�[t��T�M�����m�����anS�ع���9a�����]�c#Տ����I6aE�W�;��I}��9A�*�C�Gx�>�B���d)���.3�����9o��̲/���h�ry ֬�j��[n׉�qj����rեwR}|֔?��KQx��R���Ϻ��zU��:G����ZEa;���I��V�{k�	�Z��=�[�3~�󃨜����K�fy���|�3L��ḙ]F��ч~u�P�/���,ޫ^�ѿ���7�k32pG���8j;'ǰ��ɸ�Z�O����8��l�Y/z= ���Y	P���S$]s�ms@Q=�Md��7,�V/
�n �s�V:�����k߁5�9��J���l��)�Pǝ�@d,;)����=��w��G~v���}�uz�܈	�� ��؂9����^���~���8��I��f1�u���Wִ$,uV�7;Y��q"bd;ۧ���Ulz�W�?* s�q�V���FXF�����'�V7�S�S�kf嬜"�_3_���ʖ������:>lcz[��ߺܰ�P_�9�b��h���9���Js��Z�5Z�dʱU$Ej����v��<ܯ�[�)F���'r��m�8B��Ð�U��� T�۶_�����CA��ᢹ�kG�"��6F�Y6����B�¡L(71����4S�r�z�:R
WZB�#�l��F&������dU��j�:��0�2���Vu#�߅=�+����6��h�qi��b��9�=�<�X�we���[�dzV#@U�̽���)[�n.�	�w���+�ݍR}w�{��|1�������ΚD���uĞ�A}��h�HVs��X�=�������2��dsʔ�$�s�[bV+�PXG�ڹ�o�IǪ���PG����/N|���T^��鰿���l�LFۺ|0�_��<(��`���[$���NC�����C�eB�� �B-�?T� vQ��#��߁#��EK`"����l�;rݍ��8��l5��[�Ƨ	�q��
�-+qkJ�o�#h ���)e�:h�m�Wy:N�(���N�薀C,Hz���U�u&���f���Ǳ�`{kX٧H�bY>� �CM@�)�y�tc�������C���Z��L+^�(4.�?�o��=)o�/��`�l�w�u	�OI
�-)�煃��6{����Zb���n�U���k��A��7C4Yrz�j�`�RҦґ�0y^�Yk����Z�� �Z�.xN��A
�1#
[��z4�����I;Oݹ����	�7@h���,7����g�|�"��"l�u¦yD�;�v-(a�����Tx{��b�J,��M��C.?I��X��8es�=�k1�����ʋL�=��ӲWd� Ӗ"&���ҚQD� l6T��hM�^"��ʐ�6���xs�*��R�����ۙ�v�@�V���a�'[��NiZǯ�Չ�����8�+�������I�R��a,B>S� ��썦������}�O4N��hGs�u�o�;�8ժ�h&P�R&�O0J�`C,����y�,b\�s�+���Fk$�Ȉ|�V
�����_�WfE[��&�s����!�Y%̴L�B��SҮ�f���pp���`)��NDIj�+B|y�FH%��1�k3l���дxm�c��� ���,A���\I�^�H��~g�ߎnܑ]':E�����9�lE���E΂#�t��P+��~{�N���h�� c8ɟ��M�����Q����M/��cKgQ�],E�<y߲�t:�F�� ��?����۪��D7�H�PD�=Ac[w2n4̕�Z��A��|�4�Vp�s�,��௱j!VDc���ʥrƣ �͒I���(R[Ǖqc�*�`�}�g'_��r[�7��5�?�w�KM2�H7�!��hGէ��x�0
,�u��s�k���-Y���q���4a4S�+�_��葻��z1�&]C�R� ��y-�/��)شU��QG����fr�,54���A�*<7��Hy׷��s�i2�[�SDy�&��d��#��v�}������2���ݏ�S�o�q܍��81�r=>4�t,�O��9}�o7�-?�+A�x��`��y�T�icX)�ܣ�ѕ�7�9a�`�,(e�x"J���1��ъ�����&I�'Es/a��'oV�����M��,@������^~Ʉ:8G��hnH�/�x�Q0j�~���+&�Q��.e�kgNn�>)�z��%����CU�j)���ŀPD.�xm3>��i��f���%r	��0;�{�]��&�9@#���B��*�2�FU��1xL�p���:G�(��8ä��ۦ��`��
�	�RDi#���v���wƹ�]j�&С:��5&ol@\�n�x���ޓ��)VA�5Y��#@`��bB�8�l^ә���K��':�,\1K�_X��%E8LԸ�}ܙ�k>����I;�9@���O��7��ʣ���.h�/h�z?�L �[ų�dq��hK��z&1,�y�ۗ.+S�`�#J��7L�Y&�UZc =��%�F�����|�3���ry���S�����);��ɂ�	玫�WH��:��$+���02ŭ�rrC:�N�l�BG��tN�狃��əՅ�n}V�LԤo*���x�n��2��m�p\�$G_9�V�(ǽ�j��.��;W(L��?�a��0'�q��Gq�-���|�ܴ���4�V4�-a���o)e5��kD/AW�Ar��b�һ�co��;!��oy+ďnV�6�w	���������G������0EQ�3Z�#�'����i9zQI��Վ�88q�	¬o���1��K��A�<�Q���_�4�j����p�d�y��3 ��c�t�ϒ�~(�?��i'�0���͸;����u��q�^l�趆8z���ɂ��"�7���^JFH+	���dUQ}��0~�}k�ea�Hߦ"$Q�Hl��#��o��^��$+�iz�m�S4���a��9�Xْ����b.�PnVl���gZ��Ic}MH��f�w��dif�a��pl�Z{�����MY�U	��Y���#EU���o��U<U���1c��G%�%���·S�7ur�oD'�z����Vϻ�ÁQ�	z��P_#��.����FoV��At�^��>˯Ƃ�p��㽱��b��]�Gi���B:������~��"�t���!K�R�H/��aG�Ͱ�*�ϝC���Ǭ�x�H(☓9/�PV�����z.�\I810�yF]�.a1hy��;z�����n�1��Ú\!�z�����8���-�Z*kEr��ju��l� ��(~Aw�qq���y��*�kƯ:-��+��)��HI��I����|������<[��ZŽ(^��-��U�ׄ��=.-�?���h.*$��i=$܏�ـ�}��
���r�#k��iu9�t�rj���$�n�[� �dj�N�z9<������Ҷ$r�ڿe��3�U:���8RjR�׍���	�P`�5~�ϰ!2I�Yv��O�3C>�.-�z����U}β�0;.�����?����2ն�~��﯍�	�`]�P�fP�!$����y�Y���O��=�5@$��y 1sv�	��R��G�{odeX5�J��S���S��y���%	�0�t��f���W�(�p"�w&5�X�e2�͗n�5,}�܉�D�m~\fo!o�|PE��DᓫO�S���BF����+�cv�Y�����YȀOL������n�@,P�:i���·�n�'��ocmF/=�&�/���f��Uh��^y��9�d��l�Y�3��$�<��AV{�l��}鳶�n������] �Y�ˊw���[�i%�<�S�=5}L�j
����=n|� 75��zsx"{�Z�l��}���T���w�̜��B���5���G�X�韬��įj
CЉu�:{��}�XzeHD�u0Ywo��xx���hR�,!qa����S�k�Yh������� ༶�U�	�yE䗛��A���I���?&�!ח6�n�cP{����WRj9V��B`�%��c2=z�Ds����~{�/8���Ϝ��n�P�Ksevi��J���*Ј���*�BP���t�َ'�1�����Ղ�~E_�W�/�7h��
t���j����`xMБ�K�6��͈��&� ���x�F����P@5b����&v��a^��3"$ӹֻ��E��ZÒL>�ϔp�7T�9v��c�/*4~��w�����F���Q{̶8�b�3�Y|��7��%�e �w������B꠿�9z�T�
�g�V�Y�tхgV�6��%�rܭu�R[�!�&�X1}��f��Z���޽!Vs���ǳ��h睄�؋g�<��Q1><��:�9�!���p�(�Q�\WR
o1V	�a{�$��C��%OlJE|�NaL2�\�H�'�'d��h�@=h����X�5i�� +nְ �gOq�R�y�oaD��x/#v�S	�Q>N1V�:8�*�ѠMǁ�4w~b�]���_:������;X5o7�+MQ�;О���%����:�b��?��
�b�G�(v"�ʲ�R����E
_��,���Ce�7��9�dξ�4 ϮVt|��f?Bl�`�M�;H���l�娰k��ҏ�2��9E����H*FJ ���_�;^�+[>���4����vj-�\=$�cГ����NJ���93�@�>o�^�"|�-�f^6�{�36����|1�	w)��cg<<��)?�G�x�(�a��z���ܤ��.f��qS��u��u�ʡڔ`���4��_j��V!��A�eUO��Q���w������רN�9IR�yx�g��&�*%N6?�ڞ[�wHl|������ɀ�7n� ��S��Y��3�_,Z_�^m�24�50`�e��񱏱<(؆���$��z�,"�s0`0xR���Y�b!n̏Z^�<������]ϟE-��B�+O��hϰ����(ޙގ7\,��7q#W���+FPՍyb/�1 ������+[�7w���Td��E��'����N��:�f����|p��^�&��C�Nі���~^{�M`����9�y5%�7�(�F�����c8O�W���;�n�Y��y�NE]��"Rɇ>t\�f��bp�ޝ=��>�d���CI��ε��a��P�7�.�h��o��������3t�?�C������իX���\��[�W�����%���PK   ��xX���A�K � /   images/f32ea318-bba9-4379-b39a-fc7186e9eddc.png�wTS[�7@��p��E��<*�4�Q�wB/�Q p鄀Hi� ���� Djh!RB%�<�����}ǽ���x[�=��\s�5�o�l�yh�s��tN���G �2t&�+@�������>�-� ��G��L�Q�x���co'��'~���� )W/w��G)o?�u����ۦ����!?E�qCx�j�A����.��'��/�$�����z���Q���OjF��˷�|�-����SIi��f~ܩNR�a��k�=�\�O{V��ѕ˟0��l�wޕ=%鼴�B�CmQb)���0u���00ng�8iDe$~c�9|x�P~\����~�h���?7����Z=	b��/����T)V+�2�A&~&$����`{�ƨ�Qi��9�5�Ѫ��*�=Id��o3�T	���Pzp�:i������YX ��<F��廟\����h��R=\�](�̆ZJ���ZԽO='�n��w;��>��גn�R��Z`5*ŏ�a�+P��]��Sjh���U�XU�f�nf�	�E��t�v��6�Фub�ʹ�na�m��R?RI;znĽk)�b�T�]�<�;ᡔxMnļ8� L���`����q|rט�A����3��M��R��W;'�������[ۆ���QZl����b�v�qV�
UO��(z�V)�$�ƉPo%BsKVLW}�\��4�EJ�����8jo�/�`I<�`i��#>����Z���bc��85)���!�Fװѷ1��gf�ج���!�R�E��X��[���~NM���٢�&(�={aY�VG� SW��$���"P���ס�vr�V>V�d��Z{pp)ޚ��s`�Ď
��!d���B�O���Ň��Y��솸'�9����%�ڂ�Z�\�3?��h��� �4Y,\�N�~,��޹}��������=:^K�j���F'�S�ɴu�dW#�"x#�F��Зm�lcl�4���Z["����d�	��\6�-"\�J�GM�6"���Q���QC4���X6�`��㎃�E��z�v���7%��w��_F�!��&��:��҂���E�>n���|,L��K����4I@���j����4�����ܙ�f"\�G���_	yr3P}�G���Eg޾��$�sԄGП�?����s�����}����5,0bX�J��=�g
Ƀ��x�~	�BY������wy���Y�vc]��$y����2n=\f�:A�,%ߜz\��xj⢳�J$]�eۤ:'|^�E���z���gf&�����]h �J@Ǡ����~���-O���<�j�y�X�z�1���,�*��OH~K�6�i9x<*�I��~?�oߑ�-M=�9[Yf��$	I9��ʤ��t������ĳ�k��P��Hj[�ő�������v6�C7���x��,i�ˎ�5�n񁪌�p�9a�����"`r�!,�3��T�oz��k�Xf~>��F���'ൢ1y�I����(0A=���|d����]
������|��  ƚ�_�Dd� �6EO�ۺN�S�#ݛ;�b�$y�cr�8���Q`L��a�B�����[�[����U!C{P5.5��`d,���'d[|m{�d�ug��vu֚�l��/ͽ~3a�8	��V�,KTZ��"�}�!4�������a�H�Xݎ��Iw7���ϥ3���7�H3�Y��kp������@���B)p��_Ttj�z��ٓk:a�������� ���2���i�� K�������V�w�u�n����2�������[�[������J���,-Zc>�@PB���'
�ڪ�,�=�C>�B|ٶ�j�V���V���'���yԯOX�!:Md �dw�B�(z������%2/26���I��_��1xBէ[sat=37�X�����g �V��ƺ�������4�U� �'jFO]��r���֬�Ԅ��`��Y��V��FVØx�wZlh���K~Іkm�߶�@���bw|�{�������c�U���[.�$j�$��~g�Ww���UM��rk\u;��d-ׄuﻖ��T_%���b!���/��(�2۹u�� �������Y�F	�4.��-d�F��"H[� p <O��I&�#��x���b�[u!�R2��:��Y��sYDW/ɑ��ՖY��������B�n�'_��f�vg��2��
�,�����Cn?�D��Lx��Ƞ���#BQ�Y���7�ZZn4��U��(e���#����p��Ƹ�e�)7͝�n��7?`�Ԝ��©�x�]?����:�I
E|}*j�B�l�`d���^��4 @0F7�v�v���-1��:Z�}i��Q*�S��YF�=��ŋW�g���sj{�i����[��nV�p7x���r9| ����|��?��q���_'� �s��IuD	H?���xeY�Y��+�	r��J���(�h<����8�D�9����|�(���z�G�vJ�R:3ЧI��ǰx:Ⲽgz�������_6z�����k������t�8�����WꢹOJ��Q@򥼬�ew��~�ί���es���}� ;*H9��B5x�2^�e0�LO_�|'� g�X���|��,��`�P�������spGs�wU��юz�2z��������Mxu�z���$���z(�O]f����^�1��^��G�ߑ~�y�{�!p��g��V=q7�obbo�aɷm;�k��yp��J�aE;>������ω�b�1���­pŞV���v�~�7'" �H�~r>!{>���^������y�N5*�������] �{�ӊ^�d��<+����о��r�S�g�%�؅OK?�Ǡȧ7Z<	7^;��~�숷�Ɵ�i�
tݾ��9]j1�]7�n�V���>�j�V�hpJ�>��/��~f �%�(����J���w^�G��5d������L��3�#l]�i�Npy1�y	ZB�3޸/˹�a����cr:C'H6�ՎF�	&mgrlck�J5�>�y4#�w�Ձ�Ӌ8�إS�Ԍg?�/y��x���{����X��VXx�s��׈�f�]�7��8aV���/��q��rj}��K�Z��G�u������/����^���s,�����B�����7��O8���<�ٞ�خۙ�x�U�� �.�Pڼ�\o^��(����Cv��TR:�Se��I��*0}Hcy_�L+��FmL��'��̊|L3����,�I��ٖ�hQ�Nx�/�W<bZ�Xj�Rv��n��	��u��.#&����3�x%U��@�h��MiB�k܄���Z�L�>�w�Z�Br���ƚt�c��\�S�-%��/��~Y"	�4��S2Z��5ټ�e�,������^�'��;�0:N�n�+Sd�D)�j���TT,���Ѯy�8����v��)���O�j@�4���Mf����`>��o}���6X*��,��e���]�M�=�>ZAO�͖ �^��}Zd�"uY��ņoe%\���ܧ���s���'IX?���I�1��A62��j϶����'�n��k�I�F5�Ϟf��¶[�Ә|������g�Z��J�t�B��GI�F�-���@������ޞ��Y�Zl�#:
臿�x���O� �OJ�Gcf�;�h�J������w���t��w�l��ZlN���!"##��A~O�6���|�uj�F�«L洈�^ ��yz��
��[z�|(��rP�Ţ�O#"ܝ��ia�Q��~/��d��d��^[1kx� ���pS��yv��kQ�Q�v��et�u�ҁ����m0`�����6���x]m9ܷ�<V�[au���\g����]���i��� �z�}H�'-$Qj�ݠ��hOgi����9��) �μy`�N�$�~O/��Xh�t�.-f}�xBB�1�Ⱖ����c���U�Y(*]��4��E"��v���s�L4Z���Q�>���L[���PX�n���: )��j�{��Լ�l�L}@�~��>�$F�#u)�2�q�=�ՕH7#H �����w"BX�f�ttXh�! ��)�����vs��8���1*�^N���+�>�wє�'��u�{���F<i�Z��SS:���2ܥK���y3dB��,�]"�R,�W���r�]x�J��vy}Z@m���+�wlcc�\��"��C�������륽�X����bdx]2ۮ*�{P��5�`��z�U|5�yq�.`;�Qx�֛Eϐ�b|��	6}���|�0����EzF����O�>� �	��jW4|́\���=��,�y5�)"?�޹`/�8@�R1a�K�]����&R��5��盻��9�8�`�h����V,(�O4P��ԗ峟C��a�����p����������s�IO�*��Ig	xFH�����N#fq�v��!����bHWHј����*��f1�3E���A�}h8�?ї7�b�d�E�aa�3Q4R�u/%��]Y��ugiO7G}W�]�!��#�j��th��n �X ��F+���4s*�HsF�	��H����XBP�	�P�\��S)�q�q�Z�ng�7��
cT�ߓ*����fU���۟[���s(8,A�X�95}'���9@ �I�W��W��S���� E1���?7��n��ς�ߕ>0�*��)��� � �2)?��5�6�cZ�jI5"���� ��ݩl#���۴���S wi<�*#��X��n]2q׉�bV�c~���tS�ݮd͙��L�}DL�M`[6���0#�D�i#��~�����\ %���{r2�*^�]1l0�W������.}�̹ �5eD�rчMf�CF /��K�V�-�,u��/׹G�����#� �s"_�~ޞ�r<s�n)e�te��rG�k���D32�31��Ǯ����,����M��b1Ӏb��^��#"�c]Z9տ�2�ŧ�y ��B&Y��i�y���dg�3D#o����ְ���hۄ ���o痵|/�$���+���2l��-8[�<9d�f��~g�ɮ0���Z����W���w�J$�[D�Ȏ]n�s L:<Av�I�.mmpI����	:���d�7��G6U�lk�|d{�'����#%9|��E�R����pKEs��F�_��k"C��(�`3K���Y�!;��H a1��e�ĥ4�.$M�P��sv�����G(��Ԗ02�j�Ȭ.ͺ%B6�*�9�o{NˢT��)�>ʛe���O��Zخ3\�/⧸Ea�D��d�X$���6hF�nK6Gu
G��$�q6����U,+[$��.@��Sc8��x�Mc_����'���9:����u�1z�-۵���:��Q�0@��4��U�jl��d��Rb˘.��'���������wp�Ɠae�F� ᗑH���71o�!�����ђ/5����������.M�C6V���S�;%��a�WQ�
W��즩��w`O�r��Bh�dW��n�-"Up�8?V����]ڿ?�J��u
Ꚓi/ADh�=u��C�NR��I.�>^�:8�y$M1zr`(�6�;K�c�Md#��(���ڻŎvY,�=���O�b!$��"�q~�u���F��F7K�k#�6ekK2��G|@�!.���0:|�6��CMv�Rం#$�ZB�"M?�@{��K�c3C��G�۵b�v�������i�R ����:��=�^��)F�q�s0/��W�,�=
Gd�H1<�k%%K�^�}�����t�n�S��yx��) 1�JGW�1ZA7܆�!]��·���s٪Np�s���#,��I�R1��X���5�t�����ҌZ�������*�>�ֹ+�Qm�
b�$Vx.eyL��cSm;��O�����n�D�����M�-a�{�d��>[�eː1eoŕT� |�[�JO��Fn���f3Љ��!}�h����F��V-�6��+UV{y��f�i3�L՝�r�F�J�2�R�C�vo2& žg�����kC0��L��u����������9o뉯#<2��Zk�2-�{YL�H�+AW�E��[JV�|�r�Q[T����<�B�0rIr�Y�M5O�D˟y,��U�J6�/����Hz��So�(0��a
WFw]C	�猚�b�����^���_���\*�� ���F?��2%�B��lŠ�X��{сt�BՓ�M\G���&��I����`hy_Gn�j��b�BR�_d&�e|��Z����y��, GN<2���{��=���Dy߀�b+6F5��k��K	�af�AT[a���'Ԑ�c
�V^*_���?0�R(��O��,��_��ekܳ*��߀e��a8����\v�����r� .W�x0z���Y<3qM��^���ݻ�r�<s/���4SL�-�M�e�~��O�l�?Xc*s�9�> �kn�jWϮ�ZtUظ�b�/�h.&�y��YR�F�w+fn8O���dX��7�3���P��f�/�+�* .*�VC�Z�VX&�2�\��#}y_���ڃb�?ށn��Z��^F߬����S6Q�j��fn������q�%��^�q�oW�:���`ζ�X���h�-`��pR<��ƫ�����2���Un�*`�Z��Ō������*А�i���ŧ�ω{�}�yx���WWP����@��+gx��;�t�s�9�.�hM�5�>�W�%8�"O����,��O3��Qn�J�p���8g1�I�߷bs�#S�7�F��?=��,��֚(}�b��%�˓Z����Y�N~�ͥ_;���w2�v��s��㥜��v?��2�j����]�o1�߁ ��w�'��qc�syb��yV�������	��D ����1Zn����ӭ���o눽�~�� �9���S��z	�����َ�P�@6�.�h�%hc��V�/\o�[��2��?�yLi���n�غ��\P1�x&s�G�R��=���߈i�1tW��|�y8lW��	���ެ'��g��� �[��E4�s�wU>��c�w�O���T�Y�+����i�w'�g%_k��Pi'~8�#��<��W	��V ֭��}�@DCZ�-�i�:)���7H	ڸ���R�i��?�@��ԕTF��5��M@���[?��|?N����d��Q�+A��؎�J�����v��&�a@Z|m"B'{C�5��ōɡ�gcق�Hf �(F[(�����r$�F�������j�C�h͡]���D<g���3�|Γu��Uh{$�ʭ%GrR�h= ���f�tcS]��'�S�7{�棇�:���XX��O#_�I�+�N��H��Q%u��1�f2��rls���*10�J}6���%7�dXH`��[�����1Y�5�� >�5C#��g,Cy�rA�I|�gb�_���i�a�b?��h��<&M����7.�vF��V�zU���
��w�S��ߩ�#����ȹ|�mb�r���FXS�Z��vȪ�J�`�f~e�ȭ���_33}m	BS���6�v�h�R�6{�cԯڞ&9����̕�y��H���Ba���P3���á�rPUX���f���ʌo��!������r�����H��Z�2���P��M�PM#�m��G#Ŵ09*��jK%^�g�rXL�D�6��VX�aԖ7�E��j�:���xa��~u�]��0�'��@�Z���)�mE�!l�,���S��5f[{�+x���t�@�7BM�pE&�� �\����E��R��dI���#�0Lr�Lv��D<���"���²�u{@�YP�WM�,���O,�b����	�w2[=��}�|c5�q\/�!(ɮFn"���t8�G#<�����K��Á@�^���Ti�T,�]��-��5:�/�w��2��a%�HDx�a�y#�-�t�,���Qd�6E�s�Ic�e�s�'��'&h+��G�"M���V����.��Oe�1:�NwQ 	��l�/�L���\�m"�Ϣ1Oeic��o����DD��5#��g�M4��c:�S�^��Iޤe���b��8�v�~�ζ�ݏv�^nF�J��Ŧ!d��&�x�oDݖ��ህ��[��Ӆ���M�á�������E��)�	���-H2�3��4������F���8�X���Œ�C g]ݶ?�e4-�����[Y��k�d2xX�.����zO��������G��jA0�C�gd�y�F��)BwK1+Ӷ[+��K�����3�:V�#�H��5���.F������@v����
�E ���vki�~D����'z�=�o��@��Q 
�W�%O�Շ��Ϥ�2jp����H)��U43���d�1�5��;��F$��)U:{
����`�G�@�e
�_?�¿�Pjx��Y��^0�g!�#���\$h_Ɣ�+�xK��o!Շ{ ��cs9أ��b}����߿EJy�ƾ��q`
��:4l>�R�0����b!n�m�u��mc��t��kj�Xo���)�\Qd�Y��h�Y����4~>�F��>Ȱ)�sF�.��\��D����=Α2d����'KޚI����Q��Knm��7!�Y��> 4x�^|J�:/��ҳk*��.���Ԅ�GB�Q	�| �_0�鎧�a�EC�[�lOR����_��J�<�)d�%�e�N�~A�;�{�Q��k��xj��;�¨����V^�C��a��P�M%�����X>O�DP�������{�F�4s8��}eۉ��4����Ogpi#���C�h�^KHJ6����Rm�MN��qOFR���b���c���P��_YĜ���C�3�b���G�7R�à3&HC��gӱ���(FKQ.��B�̱)��G>pn�;��o"g� $�wC�l��C��e'jI'���@�\�IM� hI�W�e��C�n�s��MTG1�*c'>����2-�3n\AȚ���)��7t�ke������r�ęS[|����2��� Cg*���"&��ۆ�(�Y}5xRK�o]������I\zn�q`̪�g�z���,� 9�C�e<{Ő�'Nj�{*7rm%���Y���u���w�8] ��d<���u�1����!R`E%�KZ` V4�j����Fg�������̻*�1�
;��g���!]��A2�`A�YZ�K�Õ!�σ�~qn�)�{��3�8���sQX+����)�d<T��Z[�7��d����u�D9	1��ާ_3z\<V*a���?Z^���s��E���f�KFr�?	��?������>�Vn&�}������ol��W�T�s9�X�����1��6��xT�ʌ��@%
h�Z�?��譒S�D���W�����v��s�gqڧ��P9����W)�G/!����<�\L!)uM��J���e��V��r��+7��v�dQ�;��b�m�>΄��|���0������*i��\�Л9"����f���&�~�(����-�r��t��t謲o{~CD���G��s�S	x�FqZ��Yr��"T&����Т�齤T�A���{�%@؇�t��y)���Z��2�sT��Y��J	M�S�-j�ޥJZ�Z*��ȈF.>׮���ѳE�E؜a�ey*�:����w�q?a3�$�Gyd?ZRJ���6�_���������5n||�F���;|���F,��!��8�r=�@E�,U*a6�r��U+VKW�O���#�E1eD����r�߾<�e����\vE;W�}ۉd��j	����ׅ��d��W�P��bP���_7�R�7�5C��[E}��`X�����&���=l�h�-tQ�Mh>�<�|/G#l���Rf����e���?��O�o�������VNے�èv�ick�.0�W��W�����׿r�����;1Q�'հ��avH|p-��c�}�i��HB���Y����a�i/�!y���Egg�P��G{������1�͹/����H�oǕ��EC]�Փ����"#`?gwB��>��2�/I����Vۨ�4嫓�le�@��`��I��2�FE����$!=V:Q@#T>Qc��@��6��	qz�� F|��2uX�W��.�^+���ε��mV���cO�#��+���m��������k%E9�CF`xQN�X"��K&�ˎ@������n�Q�:D8K�g @G�vz��:<����%�ʭqnux�:|�mG�w��ٱ��,�n}��~�-_�:`m��7��γ�^2�`��F-
�A�O�̴��*pj�<dl���=9[s����<����������-����D���۳��P��.
��W�2P�~gX�kA�`n�ujح���7����3ad��o_�m7ck���Z��!��2�#d�ܭ[o777�¿�U�'���bm�_'�	R��,���-�,e����ݍ�#����'����SZx����;E|�ۼY6Kɻ�%�mz(V�v/T��|s����=�� 0ذ�\�p|<���[fy���!,�#.>�i�!��J���,	'�
*'��1��V[w8db�vO��̻g��i�Ŧ#��{�B����VuNk��5.Ɗ^S�V�g=���tz�p�ɞx�#�w�}Cײ�,��XشhZ'h�g�u��%�	8~�M��n��]0z�}�T�R_�2]#�����7�6G�����3q�+�Mي�x�{r�_�m��L[�
���G#"�JN������({���3Q頳�!�OT;?s�N��k�l�l��S7����Й"`ʒ����2P<:�_�:�wI����ٛ�J� �wk�����z5��q�S����<��"��P��d�8�k����������Z�~�Z5��N��_)B�0�6Thp�ylK�ѡ	�IBV3��*���Ղ��B�;,�v�D�Ռ��2]pޥ��P��g3�N麲�S��n@��~K�۩'E�����nȢ9k�^R-z䓖���5�gk�)h�Wك�D{uZ�4~~U�b'�X�r«W�v~�'2|��T2H��̼���M��jyo'����U2�������]�c��7ˀ~yxx�~���q���c��o(�cJE�Z�!�^�į��(0�W�����?��$\#̌�C�<�ቢ ���H[��v��	��PF�
fLHg?Y9AXDDA^�foR���@�u���j$��YWgޙ�?D`y��i�9����p�6�n��5M��K1�	/�aęoԢѥEE�#s�͟n��g�Bɺ�U�要���ӧ����?!t=�5o������uxh(cË��+&�8&_���܁�����W^i�������*�&]{���`zz:�s���v^����e�J W`����X��M�(w?>��C+�^j�&�������vEEEf�;���mѶ�)]��5A��Q�%�����{	��-�ie:stp�kV�2�V���롈��s��≫�km-��^��!�Ύ����<�b��JJJt5޵�_|�.�9����X=126����KKK�rrw�����G3���z3�����j�C��1�N���ŭ�0@�B�j.x��!�[�i��Ͽ��b��������b��98٦�zs�L��ރ���׫>�URTI#��]�%����
Mc�� ���}r��s�����q�%AWZ|�t ���|t�E0
O K�b� ��N���������1���`f
Qx���	t��L}�D���8�|T"���Uv�9�q�'���+//���4V;��\]��y 7οu���~,�����}�K==��g���֦���b)�SS�
94���c�����
��� $�������m�-4�߿8?�a��zl@R����}A`0**	&��ט��Z�E{�}}{�a����r1��@��%X��W ���V[r��п~�z���s''�US���?�>M9�ywJU��^�C�&E�7;U��XxG�Y���¥7�y������h��t��߿rAP�"ȵ1!��@�?��[l�@w�f}�@[����w½�v�䤥�%���r��}n&��7,�K ���	�k6����K��#��U{"�cD/��������A{��kK;��$���){T
�/.::�^)r�����s��5�	�&<�3FWd-b�^;��ϭ�C��~���R�|��0#c֕�MKL���JLK�& �n�gmm-�~E���y�{�~����J���5���[] ��c�4��G��d��X�i"�W���l��p��ye
lR������c�Ju����M��Z� �+~TR�� ���a�"�+��Z��O<����>��C446�����N�.eqz�͔�fv��.sq)((���J�a�b�+T���)��~qc��DbX��e�CY��1+�y���>��: ����-=(R��"��7�P������)�iCag���� a��Q�E��ޟ��ࣴ��ԍ�hgK���z�����? ���D��3�	��h!� �]�\n�h6�%�ۗ5Jiy�����j��¥}?LvGg�����oߌm�}�!�V\��W)JIu�	�<��k����AUUu�۷ʍ[�p[`/�YYC��e�3������L26�.ok�ͯ�w���E�y �IGr��`ƿ����. k��|<��U�i��bU}�����
��6�N��Ɛ�%
K�7n�����n�}O��L%���n��Q���ۦ�7�[�Y ;e/qp*���ghW�5ÃuX�O��S�o�/���j���l�'�F���$�0�m�3>2�V��V�؈�K���2;+X�t�8ڎC0M�fȽL���L���U-5S������.�\������z��n��(�@�����q0�B�SSS��9Qb�"��B/ܗ�ׇc.����=��ν�rx�_�'�Zk`(���`�R��k�7�4\��u+�*�^��2��H��Z>ߙ��o�P"�Mj�5E��\k����6����a<^����N���ڗ6�삨�E�K1w��Dc�K�=���q���U��n�jՀUS����cyw^/Ԋ@��n�.�~���c��(���U�Z�b����<\s7�ݨ��c�����T �k��ؑ�������Zl�:Sּ��A���@������u5٢>1�n0�FE|p�ՂB�݊�b�M�O���OaHV��Q���ص+��A��#�=�	�{�G�?k/휸t�Z)g�k�����_�aW��4��枞+�vu��'>��i���42��1OT��k���8�������r�W7/4�j������,��(���ɘ0��M��y��wC7��O��V��_u����;I~)Ǳ�w����a���X{�2��d�q��#�c������+�D1��	���C,����&�]7��:�g��b�{Z����a�*�B�]u�xjvhZ��V�j3�@S!l����V�������f-����"�e~�3������[TGG��E�z&ʩ�Y�p�]l���i�O��m���<)����^��>������\�är��HN���ڦ��ʧ�R�=�1�y�#K/���Y�~�ȫ�� !�ϼ��d�6���9�^:u�h-�y�u}��|�$vӞ��a��s�y� �r�tg}�S&�&�S-ZR0S������I�����I�M�Y���y����l�PK[r�>��=Z�i0T�7�]�5���M*��swT��c�Z�Br�m���MƋ�ܩ�Z4ӭ�Tz�4Q�N&s&�T��(B�h��8�0] �>�9��;;��;�����$�C���վj �8��3{!�[jp�n����2���C��7a&��Ǯ�T&�	Y q�7&�b*	v�+E;�i���&�_{�i2��_!��Jm�@�DKgy��Ge�-{�3�����.����I��:w��d�\�V5zy�6El�.��T�$vh���Y(	�pg:�c���e�:����I]@�1��0�HKp���X�����j����чb�&�P%�~��_��1��.�KM8�ڝ�,����f��rՆ�A��;��Y�τV+23� _x����X|Z�8&�s�X�h~�k@l�*�B�h�!�8�}�g��;+H�OxC�TXE��%�9g����:�3�ViSW�"�e<�x�ǩ��6gb�G�� =P_߯_;?�4��h;�S��j���p����2@��X�4]���0�IDkD�Vo�
�ă������Q<�Ic��^k�:�WTH ����b.1H����}uEcn|�ǂ�+Żc!SJ*�6��0G��)�a�_�c�e�,8�B��t���&�v"/Ol�bU�ʸ��P�Y��[lc��sJ��FJ_�	�ڵcq|G�yv(VS78�H�U��ǲ �)�os���VX�+�0�S����k�u���j/�=GA������9EUn9�}�#��D���֧�mY����-�2H��]N��n˼�RKd�tԫZ:������I_A�����T�������Y�	�����Q�ǽ	��ɕ{sw��j���TgaE��1@w��*�{�͍
md}�w����X��}�xj���!�[�}�HF֣�s>Y
��B�$����X���g�� ��	r�ĆY ���R��F�����y��2����.;�({��5���^�A��X�A"k˧Z�V%�������ti[���rM=˸�/J��X�����������/w �f�,��� ����<HK`�x[Ã��;�}|�@u��Fr[^������M���rEʡs؃ۭ�`5��%=�f�#/�#h?�n�$02W3sŀ����"�y�k��Q�vEhZ-Kiys3-�҈e���Js���%~xKm~ 錄��[th�����mDE֫�����6�]0u��M�pL���D%��U7�*��e�)�Bq�sT;�'�JJӍ�
��GԒ�����=I�rh��ñw�_�<1���%�ËV��n��*��q3�ȑ�~�|���4*�Q���v&"�h�5�����&��mV��c�գHǚ����1���,��G�&_�3i�z�S�kR�Bz�F�&<r�%(�-/�%u��>+$Z�*#g_G������ο�٢E>�]b�?���\ٮ"���H1��ea������ɨ�w�.�nx�ܗ�����Ft�8=^Ut�zye8��:�Ц���aާf}u���ٝsr]26�N�����a��!����2M��ذ�/K��vj���%ZV:SΞ�����-{�(����o)��$�J�6.�e����L�Û�����3甊�3�� �=��z	��C����h`��*}q�i�%�m�n5�|4�����R�H��v����r�*��m�����d��M�L��� �]^��A��K'�c���`�@y��

G/��E�}�d�<9<т��	ߙ?WYV�e=:7�^g���b�%���}P�c� �<[���d�ȧ�/ܛ{i�&fn;Y�a�)�h�c�X�]ae3U��Ğu��@=f���C��o�O�k��9����Kx=�J<��H�?��z���+~gT����٬ ܍Ԧ�y�(fC۹�r�h�=����
/p}]��$7�1A���LtG�5=��l�uFR��V^��L��Yĸ.W�)���d�c���m�#!����y������n�F��5�T�By����̉o=;H�6���L�to+�����f�������[���Ť�<���\� ���0�$���ٱ�s�l�WA�4�T�Å\@�g��m������4v�H�Dwp~�k&	-RLF^Z��,p����6��=g��;"Ã�"��,c�I��^�$"�I?d�{¶�� ��x�3J-g��~�-�n�]�Wݜ4��+�(Գ]T��c�GL��1���-����u����ݻ$� ���l�m]h��=˙NoS�@����h�=�0�55��� ���/�1�")��=<H,+԰�r��U�Ǚo��x���V����Gd���Qp�f��� �Ȭ����CEM8�c#��V��|Gsz!��}�UU�8�P��9K[��G�"����Ӌ\LR6����%>řx/c�ZߙZ�TǱ]���r��=�]UO�<�9�gP.22�hw�����u#�t�s������ح�ds��.qt�����R�\�Nķu+s�vrr��X*���vO���~0jg}� ׋/��ľd���m����� ��5��s�PyM�k��$��Iyi�����g����#/�(�Mr4=�[�/�>1�,�-
aiUz���(,��N�ѫ�F�;3��^Q���߱���SȒ<#��Α�N�ém݉�贈�RFW%#�2�ո�JZ��ݵ�4�4���+`W�>#n�ܾeW�pF�_ $���=�H�Dʑ����Z�'��:���xb���0g8�����%��q!�q����a�g��Q熢�4���gE5�]Ii�u��c����ǹ�x��,�r�� ~X�1M�j��4q�p}p�K|���r��p�U�/�@�2��F�²��L�t���=�3��8M��4��O^�.{/�ͬ��%'Z�<��&��m����/�=xr	Z8���g��lѣ����
���o؉�=�8�Bݴ__��GR%1D:>���\����@�����n�`[U�ʹ���6��m��\�D���l�i�FpC��=�D�����7鍤k�A�)o�:[ʁM���c�"�Mږ4i�6g�z7f>Q6�{G�2�Gסӱ��E�����3Q�6���(��vz�R<1+�=N|2�h.�#ڸ[�Jkl�A�dl�[�X2�l.Z�1�C��+��Fd���_N�\��ӃT.��`�(��ҽ�!2� ��<)��=�r�T�כ�u>N��Ƈ�g뮟U�zb
fLS߂� ����
�A�����bv�-����n��-:�%F�l��v��Q{���d������7���y�ڏ�,�@�շ���@���`«�s���>��g;���I1'M��Q�����^V��}M��RJ��4�t� HKwwwK�HK�������t���;����<�<�q�̞=k��֜9]q��A��-���^ܼ})E�˛e{V~�2�1���BhЃI�^�z��~Go���m�����%,�729�Z�l�if�T���"��1���9T��0�p��t��5ا�����{Jb��p��t]��g=��׉!�pd��H��w��9Z����KG�.�9�?��� T�*�S[���M��u�01o�N?�ݨ%Z[j��y�]�0m�OUa���xz�2S5���O��dPՖ�x��Fr�e����9��Ơ��(w���$M�ϩ_]�����#őBM���o@-���:62��ԛ�õ����}�'�%i-Pl~�T6�7]� H���v�ڏ�@�\��?��tl��T�<o�@eW�Q����нJ˲��w���}��Y_N�VD�<�s`�C�t�F@�Z�0�����B���,dr��e��j �U6�=8d~��0%�zD#Q5�~���X��QXN#�{��%K��5���*��>'��V?�C$N�xhl���.��z�2�N�W9�&��~�as�x��Q�uV8n_<B}�)�ީ��\vT�r)j3~V_����������s鏠|v��m_�1�jL�<�������H�S?�_؉�zK��m�nk���g�ʓ�x0����z�'�~Ml+>){Ԍ�.9%�;������"a$9�(I51��څ9�gNS��~��k��y��{���Z��4��E�C�����,M��'͖4ivA�'�E-+�!+i-��Lg�"��R��YaR�o���;q� �a��~Rid�۟�r�ݰ?�N4�LbU8��(wD���at��:d�kr��߶ed�G8N�}�b�k�ڌ��\���}��[u����ʊ[S���N��#1myy�1�3P6�I�a��x5o�5�[7�]�[�8$�h���r�e�ܳ�h����ӕT�<xN\� �<mP�t����ٷ)/�&m-[� �^ٷīH�k������n��9�&�J�p�޾��<�sR<��L��8����45�mѪ~6���ͤ�q�Œ@�B��Y��؎M�� �h�7�Q�o�^	�|�2ח47���S�T9���F�~~����k�3]n※�?Q\�6��� m�hh��9a/��i����̬^��I	~;*��~��*���  ǆy㈯��ߵ�̔(�sԲ\���D����@�a����J�"=Lc�L���>�m@��g��;��Q�=��C���.y�l���?}�z�D^��o@�����-U���w�4�U��ׂ<à�6D#�0!��������� 
�ݻ�#Na�������1�1Y��TyT�Fj�*�V�����+�9��8�۪q��8�tƁ�sn|�nM����E���{x^&�@�fN��nscd<Q��QX�aI<�)>�H�nt;����/�)��9��YnҌ?�s�)�A
q����c��ӱ��g0�q#~����n�sh�V�����k��n�!�{Jexm�H���1�c=C��~��\�!i:8�f�:'���ݻ�C�U������D�Q1n(��#ű�ζQ�(0!` ��7�+XWf���Q�H���A�T�н�gM������*}�(o;��(~CZ2�W����eӘ�밲�)M����i��U��]��<0q���X��eo<��,���㇑ǔ�?t��jÃ���o�g���&q!�t��&����b}���\��T2T?���t�3�n�ϵ�:mH�.뷽�bv2N����r<'�{�7�=EFe/PFxᢧ���W�lw����4/u�6D�ۜ�8W�*��mԬ�Ԝj���wL�n���8M�k�
�Ç�Yt1V�2�ȗ�/�~܏�N!��}�і�*?���?���'t��3[��#�!z�uR�9�3�������@����[ ˏ�,^����-U��= �z��.#iI쵌t����F�$�nn��e&֎z>��_�!���I�j�7�f)qT�k�}����z�]�}hg�nԙM�o�FNt�f�[�ġ^�J>�1�:���72�af�ǯ*}2����S�zɰ���1��˧�>\G��k&�X�mPPJ��nM�}([�jb�(�=��ͪ�T�f������X"e�l�R���]�Q���s�ٟ'1M�ʓ�uOgD�f�e3�"�����T5��[iꭇ
�W�۹�wb>���U�Z�Dk�hj�~9�q�
u^(��y��9g��s3.%�iT �\ 1��0�k�Ԧw�Yj�q�ϧ��S�+�׸�\Σָ������;b#1Ī�IVc� q<�7`�L���xLS�ٲ	BI
�[/W'/�n�:��	Ж��C��
M��u���
��Y��P��v�2ثό��a���%�\NȪPL��w���˧�B8>�:S��u��Zs�*����M~bJ�v�r�?�����2���R�z6�gC�U�N=vg�#>ޝ=|����F����$�eA>Iuv2m���`��n��M`�k��R`�U��p~ 0��76
o�[B��n)C5\rHg�,.:���n�T,N�׊Hu&J'a ������`u�6�}*J�=��>��X��pn�`�~ۗ�z���s6i�m.�p?\�)}FƁ�����c�h=��������
���6�qИ���鱋�*��5�;�Q��Ӛ֧$I���\�n�괘�)�+O0�3Wj�Q�������$%z���>7#�̠���M��F�>�n4�QH�7�N%@o��kqO�#Qaf��w��+�Xo��3��䆻gķ�����{�б�>-��u�W��;	�5SgM�#��?�ۤ3��a�	��`�'�����+ K����?^�9��;/��Y"�H������6R{��+���2:d����2��bIM;''Jo��2}�����LFU��4_Ywq���@ƅK�ӞTz�M�^�b�6�*�k~��!��ɻ��f�����䤳�_Gh=e�ӓ;�8�t�W����9m-���|w`��_ע/{"o{k���	 p,�Z��.��}Zbޚ����j���B�R*����f�s���Q�+4��H���1(P����H��1|��D����G�+V�ڨR�����Wm�P�&�$~����*��_�Fd�l���0���(ܛm��Q�ZI� �i�g?Yx�[=��X��(�� �3r�����1�
�72���Vx���n�9��A�BWj��r�2���+�dHz�][�	T3i]ѢL��x��b�ݠp�Ϸ˥�X���G�q�����������ʭ��]m 2ȱ;-W���w���Jl��<�C�L�+_i|<�x�ؔ�m�Ȗ"#>�?�7d�
{z
j"U�%�*Ԕݽ��Sx�v1�Y�v�Ԉg�;ݵ#�O�5���xE�&��%a��Ɣ�Y���pX�Lx�8�P<2�Mvϻx���Sp�:�^C�rٺ{.��W�<e�Ϟ�jl�;�l���J*
��H��wW.lP�K'R�`8�b��d]��*8C�����7vQk��-">��֘K>d��Rذ�;�� �]��xp4��k��Tq✸�1QlM"YP������=J1JU�u�%s����a����S���f�#Q5tq����#m��nl���oQ�PQ-. �M��e~\��T,+����؟{(T��H�po�s��v�̉{<�^+��>��Ih�`�}ZPƐ K�*; �֚;?L[��~sk�x#5�����9�KSoؙ�R@o��/V��x���X^�2�qOj�oL��c��j02�L�j�n��0��j�T��0f�S���]o�Rh�&�[d����=�8�E{�/=7�ec� ��Z[u�1I��HUɱ��-*�I]u;�-F]���^"�I��z�{x�ba���a�"u�T�;��q�-�*��ɵf�i%p?T`HeQ
~އ&��Zv�����J�&*�x	�� >�ϪUK�RP��L�����P�����U�.��]ޝ�������J��
��8U�����?�����/�Y���yM��f�a
�r�����`�n�m�'s��}0P?R��k*~:T�T� SoL���!���ꝶ $�O�@Z�Y�=��2丑�M���O��||w��]��U螷7U�M�����=��]S���wowe�����[8�@���࣯^�sḊ������;�`ltϳT�;�����H�]�mU�*g���K�y�<K0�H��^N�2jgw���0���,����Lg}��]O�ˏ�p�|���XQ�z1;YՋ�|AU�k �[��'7ٻ�;��'He�aV������`%�e�4��Yo�>i�`��5�.'��ּ����م��qmÀ+���&��5��
��O�8����/y@�� �۸�s¹[}���6��+�>�����ZQW��v(�_�
L
̨����=gɗ]���0��T)�-��	o9���Nf�=z��$"�pN�����l0
0�2P�-�t��� ���~��/4og��d�}�(�����9A�ί-��h��9k5��4�t�M\`�
TvR��zx�����=��(@%	*����~�6��a��e�F�����[{K��GƂw-D��eʹ)�|�Q�W�zN���X�w��g��]x�c�ٹ���vR[���e��sw	��7��a�R�8�\�*L��B� �R��`hRCd�"Զ��'0�A�X͠cj�L���U���������v��檪?��yΥ������777��P&?�o����Ny�f|u�06�p:�,�л� ����-#�G��T٩�S��t&�z�h4w~��{���P���9uo������J��h߈3��>��JW�@q�taV>~C��D'�ȣ���~���������̐\�OC��<R���%�y�ZD�ד�����;��J#[V�ܔ�t�:�\6)�?�Mt��9d�ƷyhR�ܜ*��[Xa��oq���c�t����] �=���Pp�}@�?�T�#���|FhTKJI��,��yij��g��UUxxy��i������7��Ty����% �b5U�J+�kf��:�Z7����TY�}��l�x+5�ch��O�>6��'�����K6���U�֜-aF�U�ӧ;�X��b���Ӏ������ir���G����_dy|�Y�9�'Рg�p�?�������Ui�???���#yN2f��/pٜ���T��,�F�#�/g�y�sѨ}{�8�vF��w/��DԾ=RTn8��S�5az���P�'Mx�Y���l1ʊI�����E"�����'J�w���-y~5��,�_G"��NW��������#%���Z�9*Q�*��dHw��ROhe67~>��h������d���I��"���-	��Η1��!��#`_�����2h��Sc@��R]v�k��%WcO�����졩�/H�K��
r�Vl_����¬5��m.��w:��_���g�0�A�M�?�j]��O������r;]|֤ܢ[���͉��Q�AG~��K��%M�w�n�}#E1�U%_iM���%;)����%�H�)�g���C�$���7�3-�����Z����?-��I�Ɲ��fO��o���o�/�[�DtKer�c?�>tXᖭ71�e�����q���A��JuƗَ�fV���*��a���n�V�xY1��͙,�>nx�a� �x�갥o�.��o-�r����muA�'e�؀�y��z&�э�[<��ow�JܯN9����F2�^��-����8�*�5���-Ц�ԽcY��܁E�7H��s��bc��+s1��
�{�l��� F4�s1��»Q��z+J8�d��a�)7/#��7ݚ#O��ڧ��ڙ�Jb��sf�:�wi�pA'�gְ/-�_��7�U9-P�P6E/��1�0+�[�ূ}H�z�8 ]��]>A'k�b^�K�l��Z}��ΐ�3�Ll8wQ*}�	���a[��tY{�)���y�C��|PJ�K�`8�/.%�G����������c� �� �Ami��Pֺ��r#�i#bEt�N=f�&X�s�o�7��.�|����71�m�$�e{_LC�H���",�ߜIz3��V�`E7����{����>�b}������e0��㡗eǸ�;I���`#�ݲ|q�L+H�(�$�aVp�8e�����2�o�ڄ)�K� !�P"�=9�,�eۼe�K�T·�/ӊa�u�����=�ס=�����o��)^�j�Cܛg���KE�fM���L�W�.L�2�~-_�mR\�-�@������(��8D����G��H��o�B�f�3��ҷ���FaI{>�MJ�z�8����7�2�_^�$
<�z�a��8C��> ��~L�l"Ð�(���@�R�uЉQb���ZWUU�'t��]��:{��}��{�O3�\\�.�nN�}�M�N��~p�G�s�m����k���;��P�t�"�q�%.�%n�V����t�<B�8�=�]�����"b�1�p(�S�`���y�����#���=ѕ�H2���q9�T�E�;�dLRu�Vv�z.���!���{Z�H��=��ST�M����o�����u���3Ŭ��t�<���8��&�Lr��,m��mr����eCc�1�8<�;u�mpbЙ�N�l�r't�e���~^j����Xf�y����M1�d�x�]��/+A6�>u�cE��u�ʇ�O
�Zrk��.Bፒ��2�zW©{���tS�ky�!=`��dO��%�23��!(���/V4�>%\qW>RG�V�
����sC���p�ٰ��%�՚�]t_�=p����/_��mq�6��S���H(��;d,O�;����O�LL��1���Uh�Fa�{91t),�*�;���K���V����	��kA�U ���Y�]��;�A�KC����@ڰ�=���|��}�.ϋ�U4��
!��K-�N�E���{$G��ϴ}"���=l]UF��=Td��]����� ��u6�-6z�-E��~?;�j����k$����&�@:L��̗6�X/����ب��g�������i!��Lb��L*�JP St�&��˓
��]��8�1�!��y��ݐ��B�q�(3�;K1����@��3y>ء[�?\ŅM�I�/�	݂�[�hF��}k1Ƕϲz���P��/s��b�V.�6[�:��Vlu�[�\WC�mr�z�y�||�/EK��
͠L��P>�Ψ�F�ʔ�� ���^�a1������$�G2%}����X���.��'g���L1[��W���y�Z��@|X��u��:��R�ͤ!|�[d�W�sȘ�	\ŚwI�vǢ1T#��VV%�S�����^�+�[�:��6���.�Cї}D�+zO�
I:�Nl2bӵ���3��u����C^%+�Uæ����k#�Mː	����Ar�c����@>�}ؐg�df���IqV��N���c׉���+'��oF�:1��#[�U���7�{$F��@�`�[�8H�5$/ݛp��}�Q�m8��n-�S$����e1�L@�XM���-�M-
��b�0I닔_:���ף�@\�T���s�ȽԲ�	|VK���Ɉ�ZL�.���� F��H ����(Yc�9�c�ڷ �;�Y��$���rr��7@\�$�����ȓ3��$.t�p?��ݟ��H?
�H�^���2[���F�=�s������;Q���z>yRD�	ɑ��2�(��!���s ��v�<��Mw��o<��ӳ�Ϥ����#����ؕ϶qmÐ2���j��L
���Ӻ=�:ĭ����c'�H�M��I��ð��q`p����>_Y�(^o,lll��L9����_�ɳ�&�a3�ɪ�z籜1�DKm�~�6b0113�mU��㮜��-,��J�t2�s{�?;������D zkj�q$��e섥��l�7�1𣏕y����սfl��J<��-���zdP����F^���8���o|�<�G�;n?�.�������_%�E-�?+6�P�C"�'3�sm�7�/�%Z��j,�:le٩���[I��9N:���LS
���"�����	Ѷŀe��\���/,�?�s7|V�N�#��F90'���7�{�� ���l1�3�Wǟ<�v����i[݊���:=ԑ�:�����^1̔y�̒�O��K�z�(�,�����~L5B���Sr�B�<,*I7-E�!֊�
?�v�D��L������O09[�hI�T��c8"��I�\�� ��e58?�T��<3��C'|���*�}�2jw�.Y�B�����*��4_�پb]��C-a�iB�|E'��`9_U�JRZL��vk��W���(o��#���u�5p�N���ao�]q��n�tɩ�7���q=����2fT��������K��j�(R@s9�Vx�������=/��̋0pQѣ܋̰qyu	}�u۪�nMp�+����ey2]��{y���%�xe�{�
���M����ö[>�y�C���leLf��J�
�<�$�^���r��ӸR �*���К�z�nC2��,��8��'�&|���UJ�b/z����7����m�FgfL�d���plJ�gYe�����rY�.V���<g�嗸��R��y����.��8�8�Q�����?�t+c����q��J�8��d9L�x{V/���a�G���<L�ϰ�?9�Ƨ���T�,8#���`1��_��A�[=s�\;�mQ�&AqIg�ȋ~�1=�J��+��*�mu�ʀ�q���C��M�n��4$��RG_rh���a:�\�'��k�2����V�{^�9�<d;����8�{f�b�Kߠotvq�����A�)I��qF���61���K���ɒb}J.9OY�1F_{$/�Z[|�X����^��J�PMH��r�aJ縀��M y���`��AB���DM|sSQ0th�˪k�:e۷/���\a���s�5�OK8[9efFz� �W�/p���U�����t�(�Ӫ�Q�4���ܗ#ԟE��G�jě=�:ړ�娎ѿC���VG���>�g<�on�����t��*-��@Է���>鬮([g�����^T�|�{�=Do��9z�7F|ѩ�%4mm�O���5M��*���뭢^��v�"1ҩ�1�f0b���_6̖��5����x0sD�&�2YZ�F	D��SB��v�ޘ�غ����Yu?8�����J��:�r9���p�����ЪT8�Iѐ �X��t�"�G�N�����w�{q5�1��s�����Ò4�mA2��$���tvvVWA�k��;�3. x�ܚ�A=S�a`��Χ��<OqcE&'-��ZSW��_�Sb�-N�>P�#�j����ŝA���u� ����yҢ��4������7�0U�CK+��%����e�Fj��.I��_dZ,���P����A�|�]1���o|��?K��]��8�s��#�Se������ܚ�A"�o*u��$'�O��*�:3p�����Iyqlʔ�L��\�S���L�
d�h~ʥU�e]?�J����M�cu�-V���|�r��Y�y[�V���"���^ˡ�;$�MEJ�N|��*9�	R�H���|1�6Q�7QDj�)x7����-����o~�7zSQ<�D���g,�ˏ�ڏ��Nd�{S����@��Tn�X��{*Y6t��)���L9X$7}��! T?+�,|9�9w
��w]� �E�|�!W���S�S���"�E0���[s����j��5a�,��Sd`�ӹ�����b	O�$+�k$�{T馼�v���=�2�x9�f��I��;9�H�UB�$~�	1��m�A�.}�����oR��}+���_���1���O�m� �Z��YW�W;�Tm��/-P[W0Y�`|@L�����whe�F����"%JG������Y-���Ɓ�(��St��%W٩�e�2��pX� ��d�z�{m���ޫ�aF��G��K���B\�0��}���j�P�0��tN���-���$`�r;99@Ej$�`���b��_�
�i��<���O��d~[ɯ3B�D��3����,��;�f�� �d�;;~x��X�z֟��L�	�#�/�u0��&T��Rݰ ��E|�2n��Z�[��v��ǖ� �9��7h�:v��\����f�����"�]),���i��'����c!쭆W*�+x�͒�Lң��Y!�q,A�)���TO��;6��Q�F���P5�wX�K��A_�A_�r�-�n��;GU���f|K-Ms��.�g�y��b�PQ�z?����񚰘g���&^�oD��|���ԁ��|�y�����K�ۦ4���QKb���b�ԥt�M��[��*a��V��Jb��H� �[a\�?
�>ZŪA�0b�D�����#��ȥ0$ADR��v˔B�o�	��H������/�LjA����rF�D<l竒������ݜ���1����V�Ѷ��{���>KR��0﹉���K^_�}�5f��Q�A�.Q��yn��j�o3�ʃ|~ӛŃ|辑�E&f1!җ�v7]�yW\+��2s^��l>���ә��*c�&�aQ�y����M
������e
�&ʛ����ƈ��3GMT����p��8���9��=i�[���E?�G�A�-�ͯ}�X��*�'A#�HW�3w��Z`��u����gS2m�B�W*h�2D��/��ݻk|��g|KG��kW��;jA�	����8F gSZ�U�a9$�7�'�J�`EՎI#��l@�o�o];�����J\ӫ׹��DIWHg�JN�����!,+��\ǒ�m~M�,ZJb��qR���ޙ������j
����Q�з�4�+T�I�g��ѶQ��n����o�����'�<`��7�]���wK·�B�5��O;=�É��.g�#*���o��A�[Kfzm���������e��bO�����{EDe����p���c�D*�#�tDL�)e�D�����n���̮�JI�f���`�F�~�^gA�F����s�s�����T��dF��EFB�p㹾� � %�x_���+�B����p?+:�Nj��`!�����T1�|=��5��w	B��^���6�{����d'��B=k��ETV�s?����0�t���fW��s
�D�D�DԥD��N�X��?�����w�����Am�.�X�|�4���/y�� �we�$#;�P������R-K�m*��bJu�'��_{g�u��7�÷��~Mx�4�Yp�o�`��������yvb~N�f]��F��e�;�#_)$E|4����c��ӆ�0��j��^K�4G���Ѓӟ�Vcr��l��]��U-it�@�-O�rr��d��d�O�f(d�sEvn�'x�љ��N*&��)��Љe�) �6pv߉�:�|]�!���FV���j�gL�8e�z��h�4؛F���m%Q�r�GEf�W���T��h��a�c�ե��$X��_�v#8��؝3 ����t�0'�P����=+��aä��s3(�'����G{`D�����I}8):�j��*$~�;�Ӿ	��+���p�o!������)������� d��,$xt`��<����DI��n���M����ۿZQ�� Uu��+"m���G6�o��t������E�
2��ݗ�3i����l�J��!O�k��� ɵT�u��(�o��j����{��b�khF������X�ϣ��D36���`i�����-�_���������e��A�^I{_	mW`�}����N���FЊ�:I4>��wN�w,�U�Az���A����=I��A���L��H��SIX�o��؎Y�o�ie���Rf0B����^�%�(;��rɍw����y��zp�Kp�0D|�a�KC���\����j��C�X��q[�-������߼&s�ձU�r�	V�\�J�p+NwF���r�_|>��oP�a���k�� �*�A1��v� �2�r��v ΪEF^��"��h�(�^�@%2Uad�Sb�<�?W9��e�84�+[�������2�0���AZ	]���ϐ:փ�$��4���p-X��(�̓�f�ܿWe�Id�Jb��L�kP����71�үA0Jя�ɍ�
 ؛�j M�_.i~�H{	[-�)J�	���b1�69נ׫�;�>L��ëN{�ŕP�`Vѳ�����¤C��S����_�?'fm�܁�}�]�٫�����g�9��-���^^\��X��hR��g+��&�'�!�����"�����A�ͨx�ۖ�/� O1�����	��榷����[6ݭ����M�2�c��dk-O��k���d�f��8�����4�^K��#��\�N2��e��ph��<��Vi���M׷3��" 詥gU.O���5̝bUQ��74�|��6�nl������pKv��Gy}�wp}�vE����Xũ�I�Zx����o���y{<�7�ƕS��F��&_��/6|��]�B�R�y��1��r�y���C�χ���+g��?ߴd�����b�]dE�
���֨��^X���" }�q�&�	���+I���Hf�i9�>�
��@K���?n�=r�M�Xd�i��,jH-k��~�kZ����]^5R�H� ��rVVf:���p"����l��n�/,��9�43Mv�<���H���,�F��L��.2.��gu
�g�Ħ)��o�i��bR$�v0� vF:�6K2e�ͥ	Y�%s $%�đҜe��-���ByK�݀�5C�j(���rбʩ2$�l7>��*��:}�'�5����I���Բ��Ε�^a18��dق�`T�K�Dݩ^��S4c�L�j����;R[�D�������:�����_?��\��frn��sO�
�I�{�}CIY��h��Pju�~���~q�2�ܬ�b
-��ż�Y�����{�3��)�V�AmX�>�<���jIyܮ5��vSS̀,��Sj"AcsȧR?r{��)��e�T��y4-af�� �Xd�Z%�;QP�١�}VTϞRI�*Rɽ����㝹�E�XLAOh٦�>�����q���@Ua�Qb�H�?Z��+�員=ҧ��ԥ�4n��ga��5�[�d���7���f�%��vh����t�~��+T�"�.��l�h�$�nO���2��}�N΂�\(�X�J��'�D5�D�H��C���6w����� ����WCH���h�?G�(�(�}��3��x���Y�"Ǌ�]�n��_HWa=sn��]'��i��wԦRY�	in����[w���{`��!c`�&mȗ�OT("�Ҧ�y���՝[;I�b,`OVǸ�.y���GzF�b g��ߗ�^g���I��&FF#�*V��E���Oa� �'�G��G*�,���W�*�黅��3�k��eƀb�@�~�w����F�7t��y�,v�1����@&>��l)���Ha����Y�#ʙ6��Q�M����	�Y,F���VFpt�$|)n�b�b,!�/3补
A?��t�J�̌c� /�2���<L��}�!��_��C�V�G�q��#�覦h���5�H�WRO#������^��n�c	Y$��RT���\Dg6�v��QT��b�YD˥�h��rz�Y;� �3�/�d�g� L���T�^���a.d���N�7�,P�].|m$�;w�����X���=8�T*쾉5>���_N�lkR�xb����^B���~z�l��:�S7�2��Ǒ���{ի��7*;�c�����+�B�:��y���,s��
�Cu��(�2|���<$|��C��P�ϖw,0�� �@Sqm:��^�_ҽ8LpDHj)f��5E[0������3�;`֐�+T`V�s���p@
=eWNm��#=߰O$�ߝ����L����ǝ���/��;p��I���čP[�=���K��kE���)�[0֎�B����������d�3��m5[.3�M��g����ﵝG:+/K���W�a�E|�U�+��
N��#@���]9���y�O�pw���x��(p˚;"��W��9܈��@$��]=�����֟���'� L���"@����;g<��K��A�ڞ�mȇ�.x�9����#t��߲�K:n�.)�	�1�?����*�Fﮫָ�}f�?jp���Y����Qt����;���ձ�7���>��x(o��3ډ�C�NU��i�h��V���7e��o6����8�rdb4�dS91FX�i<Y[��{�RꁵۄáZ��=a�|"����kp4*��A��s��wC���ֽ��AץP�ŉA�/�>��У�Ga�v��{q����QC��٬g
�#O��B������[9��ޯ��0�]�-{v����Ǥ_~_q������7~We��"��^x,T>J�W,�֡��9vwMd��z��c��?�_���9�|�
��Oh̰�64����by��ٟ�<��tb��2��Ѳ��(��o򟆜��Gm�s�23b}/�\y=+�V��)��Y6�8�?4wu���4���u-�����FdgS�됴f�$Ҧ3��v��2.sc��ȴ@4�
 �G�����D��
�e�p�d�I̬���v��_�	±J�NH��@�J����Gш':P��[��U�t�+&�W��h�C�|�'�F��Hj��T�#:g�dm������l��_�d��aR��!v�>�3�yI_J���jw�a��f0�#��~C�|��>G����{�����W��H&wg���u�%���3Q�v��yS�
]cj�c�h�#�/e�(n� ��)�b���S��\���t
�i����k2
�k�N�&�Q -��;��*I�~���<���J�����\tig�q����J�l�#2,*������ڡ�M,��s�����3��,��v/(��Y&nVH��l/Ny��q����Ec7&�&ڍw2Y�b{m�
����6�t��d�Y��'�:mt��iD%��������ww�HU�e(�_0R��d�	��`���/Ui���E�F���m_�0%��|ӌ�5�X�%`��0\x� �1�'m��O�ԏ���/�6+�u���BQm}�:�rC�Zef��0�~�w�c��O�߿Q7Fc�⋹��J�q���,a�@���G6��ޞ�ֲNySk�3����LG=��_Ҡ��K,��\a�k�o��0lf�ٮr��������������UX��!�~�u�͊m��1��WC /#��w�|8{:Y�$�D���p6�+��/��E _
;#���#z--a8���85좤�a] ~����ʿa�3B����K\����0X��u;&9aIظ�&r?�ry�;�yq�K��� �����T��MK��J���#��T(��F?0�7sX�� ]	�n�A]-)��^稴4����=��P�j4���T5m�g:XDP��������+�Z�6�[1�����/�*�%�U+�[���W�X6��\��Vf�D��P#�1q���'�mJ�P��M��Մ�WN�{�AN �r>�+lm%�r(c�V���c����ś�{��`�+{�FR�C� �f=�	V�u�E���8�P5n5��4t<�an��˵P�#�~;�e4c�0c'���TӨ�ȟ��j�Au�����'�uJA����F��7��g�ձwv����v]���{�2�T&�@X5��)m�M�Y�kRa����\�ZqwS���y��� �B�dRp��H�p�OҠ���D!��;�+sC	����Ed�=&��������D��θW���i��b�aJՔ�j4fO�^K�������y�P���]���z`��Xt<�Lh���`�0K!��=��V`��X�r�� �)�U6�y��8$r_���� ��~��e]��\�CSD��#�3�MKR~�TF���{��@��Qh��d$�Ur� �_��s����s�͛=`$�����)3��mB�qED��`��TA�ͽdWY��?�}m&�ua�
4Gϡ_ܱ_�/��5����8��B��Eֱx)̔M�Q�.:�-�2�%Yo@�["A��� [��6�ؗ����d�s�˒�Ŝ Դ���ܪ�g4�����b�y܄]�g�W4���p�V��&<P�x#2tشR��ɶ/� d�	��k�%8�vv������ks�����_n�C��dJ���8ϱp<�W��%��-j�nR�d���.i;��FP)%���>
���)@u��`�ȴ_�g��M�CdϤ���Q��t�H 1�ZU: �:ۻ�67`&����OƹS���d�����񨅉6����yD�f�c�\	�v����&��3�������<��ii������~�w'�CڞN��F8�cN���Ӄ��ma`��,�Y�K"���"#ك���w쨮�,�5sO��9?�!�3�3�d�F*i��~��A��.8��Y�x��Ǳo��7Yvn�t��o��ZcI�G;��A��t�;�Fx௎���`����cj�*M�X��*���,���K���ewj���(6�D��.��v�������=�h��[��խ]Sٖ�&���_���#�"t�rޟ��4lF]�!�,D�)Q�&��GJ�Qb�Yya�1�/ů��D)�'y�y��4�P�]��[W��:�� ��G��R��28�{�5̣�{ۈ�ۀ�^�����G��a�9�Fb�cM��((�gY�(M0���,<͵A��r���S�|���p�����|��0�GD@��_$��L�V��~Ϲ��; :�]����` E<��1��{������PQA:ҋ��(�H�.�/����K�,��"��tB��#�Fz �^�������y��sgn���3g�'�gϞ�9��f�8�齁2�j��:�m&�4ns��-<�A�Cu9e>g�m���9�mڣ�Yj=q��\)H�>�|�su�*qp�e�6eN�K���p(�q0�L`���-x ֒�q�W�h�UX���}�P̥w��J8��'��V��W�2l���}X�WʫQ���j��m-}��Z�$�q���1�7�Bu)>>��*��g�Ϡ��Lf��N��1Q RW���)�nC��킭ɠ"?\�h�t��\�(0���]����4+�e�9]R0�ǋI�{k'�I2[�Yv+�o��l�OF�͞>�K淵.2vt�C��@����z�7�H�/!��o�?��i�����:8r���pZ���"qI����m*�1���a@�QC��2=���Wl[k><p��"�=��q�yn��K-��K.�l����0'�`��%�
C�}{��-��O�3�_����Uً�"���œ���Ig�WW�F�t��)�3F'�S�l�ߦ�2��\�2��9չ��~,�^hQ���#ߎ6�g��^�ǘD�8���A.y�>{�4�ya�g��~���&>�O"�uZ�7�����go�������Rd(�>�^ �:Q|*�����	�봖<"�'�8���53��)�dj��	2P�lM�_������r���ւ3{@����2y]A�5�F�ZBQ�c��E1I6�∎���)l�Va�g	O����(fg�g�WV ��t~��\�<��������pO�C��~�˷�m;q�Jj.�� ᗝF-�-fߘ]B*�7ke�.�*���-�iz٥k��*��*}�A���G%o��?��Q����LH���[��0{<�O�á�7��݇~Q2/���/U9�Ip-!!�E��I̹>�ؿ1T!�?��r�C��gr���AUY}��'3��p��ȿ��WJ8�z:��[����G7=��Yw?�Ȥ�Q2����{4q����~�������ζ���ce�o�O��O݄��sD���\����+�n��\��+����D��P�ɧ��G"]�?���)&��"�W�Rt�n����$�=�D�������|����yс�[Ae���E�ǈ?���ˣ��-޸��z�v��}h�k��;W��zM�N�_1z|U���Y ���7���pU���}��0�+7������>�`�X?c���7�{�}��Y��
���k�1h���|�'��R��"5�׼o���_v3�E��@ �aB�f�pD��$��q] �L���d!�*��h�
��?j�~���%''�w�=?&��>��7'4}@�X��HV�a���L益$g�� �d��3�*i�&�+��<8��ػ8?��9��[z-yK�0�L��8�J���G/�G���ټ\��S9��j�J�Ԁ�DP�� �b�U�5|�l�ȵ�C�cQ��A�LKw��e�3����{FA�"�W�E:r���.��<Q�ȅ)>�0&5a����^��D��� ��.����e�k�l�#ɡ��q�T�W�B�F��ʥ�<+ �1HG7�t������<˘�!��T�Y>��-L�}@}A0�]��9�W�����w��{Hқ�I��kl\�7:{.y��{���7gWT�!���^�&!��ƌ���<N�5��pWk[I�ݰ�$��i���	˕�jl����)o���|��iMi�\�6�m�%��D��E�(2����ߣ�� �|fw_\Y0ݬ�;���F�J�
>Li���d��32}�ҽ��!Ū�UЎ��Kv�����?�s�*/h(�b�m��^��s���ērN~��@��ō�����-/�L��yj���&�aqЃ����S&���6y�ѣ���S�$�Ɵ�ͨYD�ĝ.�&>eV�|����;��>�iQ�10{�Օ�-�G��xFv��)O>Ha�`Q�0�N�А��i'�mQ�;ߘ���	��ԁ�U/W������o�/������Q寣c��B��'�+78���G�GCt���7{v�1ӧp����Un�]�7�u'���a�I��y����W�I����Aˤ�����l�^�2��N�����^��a����ڕ���=p��M-.�M���i�nK�7N������|V֝�ࢹ�><�흠X�^�k�զ���p�[o�-÷� ��o\����hˠ��1J��,̕�9Ι��8�����n�{]�Hj��UBKb|��^��P]m������#Q��Ź3ml�Cv"~�<�8y��S���캅rI��c�=���Xcl����BO��/���������ֿ�~�-M[���x7^_�/�6�+^r��r�e�R'}��C�j��Y�ij^FƸV��j�W[dj��<D�5w��=�̸�=�gR+kz��MsK�&*�VP��f�;E��q��5Hy�VJ��W8�,u�8s�Fl��r�8��v�3G��ۼ��˻T�<�������Er��QM�6C�I��	��51���a:��Ԏ��,��{T��7N;�KW,��L�m��Ӫ/K��|�C�6�;����5������o�r!�H����Jm��^]��-��P�_�?+.��Yw�ҏ��i�d~_�q���Ǿz���A�	�����{G۬g�e)�0�>�������Ͼ���fI	����݌S�ĺ��|C��qY.K�2O�O�Ʊ@w&K�y��ӕ����[�t��P�p<�*3���/���kb�%r��[~�X�Oڋ<n��ys�v��g�����%�ۿds�@ŀ�V�	5�k}s���m2��Ɵ��ӻ��G�e��&��0DNm;��?"�b�����9Be�ґ�X2�����mr&O�r���%>P3/zc�\��zJ3�T��ꤜ��P �M�C�/���U2ͅ'!��qf��T4��;�)�pQ��^�e|s�}:�YN�6cm��/U�Up���o-��0��HΧ6�;.G	:ӛkeQp��Ҿ�g,�*��P��R�2�Hs� �ԫw���W���I�.S����fs��.tw�0��1�Hj�_��ҬO�%}@�[����Ȱ�0��!�y@y������Ǌ�g(�F�lď.�]�%�ȿ���y�S��V�i��1�������+ٔS."�4�I���D��i5�R:��L,�OZrs����m'�ɯ�%�Pm�g"�@�P 
f8�q���\�\b���柭�äȧ�hA��5�h�_�m�\���Zf�Q��s��y���$���S�ia�zY3����B��#P8�^�o���������2�Hd��f�I�W;r��k���ū����XΕU�P@+�S8�X�����ж��b�����A�pC^���5Q�z���8����-ya��?AVbiL���9v;n��t��`����$�V�I|k�~�Y�;c����vE��̢��ڟ1���S)05,!_\�]�V�8��:e�g�G�ouZ��#��I6�-&'׾)||��~����~���e��o�ф;�^�h�c�Ԑ�oz��4�u��"fo��r2/ F ��iv=�v]^bDZ���- ��g׉��7��q��z-Jc���O?�|��d�bu@G�j���'�_3<����+��H<�E16��,@�P�ӵ�؛cK��y%�ݦr8��k�B�|��`�+�Q@����ŗ�)��J�3U�W��f&�;�Nw��]���&�:G���9TTᣄ�!9�������K��$��P�'�#'/�������R��n� �36n�t� �6,�(�{ת��5��޼�}�U僛��ol��fd �=Є钻A�¯͹���eQq�߄V_2_��ꄹ��]Y!�,���<� d�ZuJ���Pg(+m.#z]t�����$/��b��T
��?R�����gZ|s�m\&���T8�_8):5�Ԛd��N|S�uNq���S-��Ѳ��b	]�[����g���la�֯����p�]=�!� M�JȠoy�i��DɝBv�d��`�&�
���K�kZ�K�����j;7l��&q<I�)���1��g�ˉ�R4^��~|��dv�1 �p����\^��d�\ 8�$�����P6g�9�Ԏ��3�.W[�ޜ���=(�24���=�k�RQ�O��*
�e�g�y��YK�"Oo?4��:��U��oX��k'����R�������t&՞1P5�������ܸJn�� ���Ϝ��u���3���鉠��& g�x�BkăG)�O�D�2ڳ��͋��)�/��}�Y���(���v�Sj�Ãx�RI:��T9�gУ⋜��eu/�aߛc����E��NX�4��k��^�&�>�c!9q=� �.��ouXq��i���3����y��}��AilY���Kb���b�;��~��Ϭ*�i��]�:�ٍ*U��j�)�N<��}�)5xz���Ra�V������en��u�Ȣ���n�7±������T�	����{�e,u�m)�����W�Ɲ�AJ�l)xr���;=�զ�I�o(t�f�}��͋�O-�Qz�d�M�I����J�����J����Q�1�AN������'���{��R�4<�����<�G�xJ������R�U�4�j�+��Su�� H�B���c��j��^��~!����oB��N|#)y$EҲ�Ȏ��yI����Q�C�d�SV��?\��sCꝽ=Uz�D5�����[b+�����f�W�;���c�El�&#Wn�������V���͙>l��?T �M�}�������V}��	gM��k����ѺW��n
�3g=�y��
��:��v�9�.{:���?���j��qlէ��i�.�A+e_k���{�tv����;����נ�&4<]{w�?$��7GI�,d2�w����{.����f;�!��:ȵ�oR^��3�,8=��n��)�|��9���	�,���^��ʺ�����Y�#����4�}�_o׽r���1O����+��l[<�UNf�L�d�+w���'ExM@0�D:��f��7�mw�w啭��죨Xgz�RT(�����mk���O�%�TD]ۿb�2Q��c�ɘ4��@CϺ?����o�$d��}�b��~}����q)�ǽ�g��n������N�k�f���q�YY�G� �ɯ\�o�L�iQ�P�p���P�J�I��v��K���Iމ�15,�p�S��2g��1jR�긫�욫�Ӱ��t������!���S��Zl��i}������b�|��1����v�3��l�{7�[(N��rR��!~�M*�v���qjg�q��$u2.�[�G�o�ǝ}�)g��fG�iF+�>�B����[v��.�VV�+�2�OAe���I����Fx�5����G:�R�Z$p��:I��n5:7�OZ��q���X���Zh�/��r>���{��:;��<?;v���8T�1����g2������TaT=��rue%̸��>V�H'܈�AJ��q|0}�n�mG�+`��ċ��k�E�j3���[��u����#�A�u�ޤ�_�~��~�Z�V^.$.!an!� �o�m����w�zf�v:�n���K�E�Nܾ��^=���@)ZJl��X�˳g-��5��1�2w��.����w��c��|��h,���{>�Vb�^T�k�?KiF�z��6�ZU�׈��|��6�Z�al�M�ຓ��fkG���/V��ax9w�����ޡ|���.���H���,��j��ԣ��:�*�/��y�MV	��P�J�:555_SR�JKKmF���a���[��(����̡Rh�=rW`�Uv�򡇨��� *�T]0�5��☽?�t���w���C�uc͜w�Z�Ğ~�U����r�N=��־���Y#tY��C(7�m��N���sD��ɻ�6��)p.�����_E�v,>�^�;��Sc��`�{�={#�1����5����Quw����a��jQW�x���M���O��B������_f��Y�j�FR����ǳ4�A�}���9a������n�څ
����ӻ����o>e���dpt��[�y�8v�����|nH׼��6�c�ڭ9�?}M��d\%�
ɬ���R�Z��.O���+Y��G�����E�'��<��,�t���;�&��B�`�Jx�3�1��B�|�S�Q�ꕦ�@mD�8�K�^�3�Y;ރn�iՊ��H�9&7O~�5��._c�Fn����k:�[���1�{k@½�XT�[q�)�����d��Ar�V�l�c��T�t�	����kk�s��;�D�UӠ��R��	c5�S���:�����G6�����g�.��)ѺUY�ќ���� �Ӹ]~����܂.����*��>D�,����y������%(�u�V1����N�y�ͮ>Ys�Ucc+\���P.�R��l-��&豔������-�˳��>�Vg#�df�9�Y��b��H1�)}����W�X�q��^��N���^�'����ͻt��m�&b{�t������4� %_���,�~�1�2��T�(q`�@�6 ���&%���\Z�%6��k'1��3�	�}�;��E)8�Yy�'U�-MJ��N�QJp�"��;2[�z�� ���\Oċ.�ZMJ�;�"�45�]rё���3B�k���EG�~*=>��^bJ���꒬=|��d��~#��O=����\��-�	���y�4�%Y��I�8��)����]�c�w'N*Ƕ�:$�'2�s�Z���������jUg/��ɤۇƭ�Ƅ�6?���z���':��A���_M#s�V�0Dr��5��Oq�6�^Y���:4��(�>@a|[�3ǿ"�q/��10�K!�6@����Ϫ�i�?f���+r�e�L��O�XT�<G��G��s��۫&���6~�K��I�@>�+��1U�ߙ��x�� 8OP��f�f����Tt�v}�.?��[Q�Gba��4
~v~�29������J��2F���OwX�i&{	FI��/�9w�O&�T6q���LG�<o$�4���?h4�泇�(�Z[���,���}�2;5�aK&��hr�v/��(�;.)�ׯ�~�Ӵn��J9N�HIgi�I�w9pt���i�z���T^��Ҵ�<�Q�R���QV竢�6"V�V���B����Z^XH�^r�܇�mq�����:��+V�szR'k�9��f�'
�j��k�S��>�~�}B6C�Na�k0� ���Y̘�a��痔��(5�W��;�������T��0�!'ͺdhBROz�7c�2e�ۧ���<�m�\�Di�^�鵵5mcN�Z�^n�uP[�Y�8Z��������Q��x�64 �7��n���:c8a3e�Ph��}�z��ާcL�>�@}�?`;�=�Qf�92�O̪��ݏe�8~�f�0%v�>�֦�S�׸w��>���w|��M��S��E�Q�y�cׅ�������#������l� �������H��1�g�_�!B������HeK=�3/h������4��;�g��1�QԈ���������R�K�U�|^M�ʘ���{$@�1�Iҹ-�F&P����Z��������r��uSK}.�Cl�i5cT˱U
������H\w)�)����"9���g��2�87�#N�@
�{ˈ�u�F&��������F��q)ln���	�-�& ��b���k�x��v(�Ĥ��~ E�.3*�T+|�>�+��۵l�[�mf� J�<��D|#������ �����1Ac��ѭ���7��{� �祧�Ƥ��Â{�l����I6_O�hV@E�c��ڶp�$�|���^]�H��6���P�*�Ùα�&�4�yFo7"��**(8ث"$�>gsD�Ro�>
�k@$�ٳ�JI7�f�(_��f\�5l\�T�u5f�Y��n�>\�*�e��63maa�;{o�k߰2 �Vsw�j��o��%jC�5ŗ��I���e��i�4����N&�DD<q&+�~Ҹ5>G�Z��0P+�g�޿��d�3c�}ʇz��^��jE��"�B�3��8"W��Vׄ�Nֺ��ם`�4c�d�.窽t� ���5~�69p���~f��f�Y����Y���L1=ϡ�]�_Ծ(ox��g�m�m��=�����:���D�&/
�DPc �K��݌�(Q�i�BBB.[�we�u.�^��/cc�;�B�Ϸ�_Hdγq���9B�e'�[����5��"�1��/y�d1:��q�Y��b�W�����A5v�Z>�
֛��u6�!�a)㫛?g1?d��9�ڣ���q���:���';�L�7;Oidx��$�sL�^܇@�Q�٬��"fG�4���qk<E��t�|Q����������I&��4�u	+�΃s���+ާhq<�BGF׸eb�n�#?���c���Y�3�ׁU�([!�_�� *�IK0���%� }{|��7���Cūf�r��fn��uĝf�	2.F	k�'�q� ̈����d�=�'/��C�!-��<��b�Tr�;��ڸ8s�>C�(~����f�u�C�?幂=|]�T��ORI���( |M������JP˛��K����0Z������b	t�k��bI6��ծmE��JŎ�S�2(����c�_��⸷9��a�c3ҷ^�-���0W���	E�Y���^z�����r'婣���]葵�D��$������	��J  �
�C�<У��Q$�Qgc�ɚ���$�O�Q����aQ��0�#2��|Ķ�nAv6���DE������{���Hn�{��5�q�[c/6:}"�<�E:S�zݪ��(�RF�ҭ��ls{�{	=n�!���cCEG{Ϙ��?U�u���1T����G
|뭠P|%�Sٚ���Rs��%�D�&*������D���Ե�\�yS�W0E�{�Ƕ�9L"y�r��sz"�kv-2��H��$��Z�'���5/(q��{�|�r����zʯ���uC%��"&�K�H��=e:���)"$͔
7s0g���Y�zg�Ϥk\k0ku8���K�Jc��3̚�))��K�5�@�J�\r���iF�il��k��%)��]=J��gS�m ^��ҏ8�0ƹ��ۘ��i�b�B7
�����Y���4"H��xF��� ����2Q��"���9�NF���>Um��3!�g��>c/�BhQ�c�Q�Y�Q�iC >9~h$z8�W�n��_/-��zd�ɡ�%��9�dF	�JK{����G���IE���i��a�ydj_L��_�l�:f�׌��62��	Hܲ�������9�W̻�.(�+�X l+�{z�����uϿ&'#�"G(͟��C MP �ӥ�#�m~�O���.k�x�v� ��>(�~�r�^�5?~�f�X�xݼ:ϼ9���-��yԻY�+�s췰{�{=b�`�J^��2L��M��omTRj�?9�w.����܃��3Ne�Ȁ��?�g٧�U.u�&涮��t�&�H��2,�{�{;��� p�@c�Z�Q1c�jۙ�K��ԙ���z��F�&�I�b����38A���qw�f�y���e�%I(&ԡ���e������5����M�����]�����׽�.�\�oz{�,���l�u��ӞF���hE�i�#�o���XO�ӂk\����v��B^Ԡ��>Z�V����d44r@���mC+3BIUM�����_��)511",,(�a}OD�~-�c(z��V�x���F������F�>m�I���g�nC�q���n�pB��@PJ����VP4n�g��?lffv3++˞�Ҕ��2�(:���s�Ae�J�Hm� �����Z	�F��B�;��ͦ�`mEup���)�)	�
iA>H�����ʤs�@ccz�XAĸ�Qw��,Ӱ����zF)v�飈P����Z�c���Q�����پvI}0�|eOQ�P�����T �'(A`
���!�����gE+ �����x�U��Z��HWG��H3#&���}DPj���D��,�16��w�������{{��?%��j�b�[��m���A�d|�'�m8�j��mC8�i��,~-xX�or�����05'�})nn�oUU�����������;� ?�¾~� ,��h���93�	�����r��#f�Ǐ���d�]K+QK�3,qd~�B�ж�.p�f4DH��{��Ӏb�������l��.<���m����b�!���`RE�Β���4
u���5��+�� Ȑ�U�(,���x'?���۝N���~�Ō�fn�8�L��4[�⃁�����%0��c���Q���Q���%��A 3���(=  V��/s-��B ��R����i@�ǰ8�̗�_޻hpg4	��T���߿\ [- [>n�=�Z�A_',�T$�'��Ij4��K�;T�~�Ge��b�h�	<�.�ߴ�
�������ꩉ�w�.���R��w=q��4H(��a�r�������k��ݘ�6���Y�L]=��2��a���yǥ��eOp�$���I��8���H�t��V?o\����5X���o`�w�4�ۗ�?�z�u-�h�Տ&عzy�nh|���SB�����p!0 ��d�����R>ҩ�))�,-�r�qo���H�ƽ���O������W���s���Ƭ����$���fj�}�F�|<�\L�1���V t�c��2�wMm�l�F����]!W+<>>>g�V?�-H.��fQ"���? H� �i+�<�6`c!��9�	u�Y+x�Ț���bT4�Ƙ9:�/--=|�ar�:�/��V���F�ʀ{X�3���0��+ S���>S����f��ۋY[�Tʠ��9?��ɯ��X��.�mWF�0�/5��.�U^�o` ���ppu��PB�R�$(Д��ś�}ʠ?��rͿ=�2����~�Z$�7�S�Nk)�9	���BLxl7Ϳ���/�}�w.�LN� pя&�L�nL�vG䚧��%H�w�KI��e&Lrr��Gt��n����(��y� �B���ư��L?w��e�$=36�qx�S�lߢ���#���]�e줦���`����	�"�Ng2��N\W��|;�!�eHD�N~��<���O�xFa���4�����'�i"*���[�@������8����>�Q��%����j�e��)B�  �!%y�}/!i�DJ������Ti6ccc`��cH������c�r+5w���k�#��f L����q�����<FH����S�����<�l,�&�g7����q�;���~<��s�amiiѸg%}�ݹ>v�ҥo��X�ض�q빭�_($vl� �`����?�>��`l@%�1؎㪰�հI��!���
|�H�v��>�M��Ѷb�����K��gn���4'����W��@�=�h0���JvjFV�����>
�Ne�pw�B� ��,��� �](J:1#�<��"�����N�}"t&ۺ�w� ��0mf�"�S��א$�B�y�@��L���SU��O$�qv}E����񵮈�Q�������r�DX]�	�P�8O�a�f���pR[�ge��8��C ��+�hJoL2M���_�m�z���J�5��j���XJ�8äF<��On_���S����f��Z�Ox#h �k�a�!�{J�_Q�=�P5;����7t�菺�]ku(����Cd�b�ņ��ӵ�w<���؜J�����Z�+�Ha)&���+�G;�^�,�gμ��nit���"tz2?�wh��lH�܁.��O���YA,�N"~[.�#��n�����>��MJ�+����}y֛Ѣ]j��V���Xp���Pts�����ӵ�g\e����`���~v��j��kG��l���Y�{.��Α���ۥ̧��s �by��$�]�̰���ȵ��h�
���4x�,��s����yW��M���ٽ֩o����N�7��Y�8RsQ�����Gn��,�%�PF����lkƳ5۶��O�)��w�_�%��
�ln��������2�
�$u��iI�cm��H ��
u"�Wu�(�%��o�����ta��S��)c���լ���AHC3#���m+��K��՞,5W^���
[Y�\mV� ��9����7�����=U��A�����0��K��J)k��z����J���ĵ�hm)��0^���c�n��Rs�C�L�h[��hX�펒y��f_LtB��Tu��kG!l��H��^�N�Ki�S��������]�ʁ����|a8X��3�j	�DE4��㱟����������Hu!	��Ǻ�ʣ�liz@��6�1*\#EƉ��n>	Q"���?r�'���?�EFQQQ��K���oE��O:�/��K~_v�S�-B\c����`�)ԏ���¦\�Gn�+%I�D�bJ:6��������X������45/�'f�>��y=~]�aw��o�/��� ��р^ !3��tЏ~�r�z �_�UHs˼��w��ܖmɯ]z��<�|������ni�V���p�7�r�H��y`��|;b`z:y��vQqq_�Eg��ceO���q+�vB���?."Y8n�n�#��.זk�R�?_ʘf�t'w112v�\x���A5QK�g��g�܍�������(�Y �����"��A1f�'�"ȅO`y�ى>-9�л�f6�,�)x�K���X	�J�'Q�����?�/��K�7Jc��A��l� z��Z�hٟIOB���[[�]�J'.xB������/�Ǚ�r����P��`��X��w�?C
�}�|��Pw���ji-4����8��(JR�g2o�1��><��UiՓP�����$��w#��^����%I~�4�6�(R6�X�
hm{�;���owcT9~կu�����
�_EeBB����h�~�ֲx<I�53�(���IE�๠�s�~�gw�W)q�Bl5ɽH �w�n�� i<�i��_�X�s��]c5�|��y�^�����%~u0?Z��*��>Q��_�/�� Yn�� _�*e|ܿ|;o�V1�Ӈ<PQX\<��L��g��r�E��PZZ
<�aB���} 	���#�I(�"KHL,�!2
ֈ�V.�V���PsRNT+����)8:�_}�������]��7�X�������w���C������`6�㝚��_�>�X��V}��l�0����,�p���$�����]����Օ��މ��g�W.�|��r���OXtq�=��(�W�lz��ܛ	w&�A�Q�F�ʀ�#VgG� ~�����ͻ��'�	g��\r1�"�=K�����,_�@� .W�f��kjj��� ��P�������޹炸.ps��&)%{�2���ö���?�>ȍ���� ����
�&d9��b���}�W1?�~?��%�x�F��ί�4���X�gj0���)#Vqw��J���in�	=Y����)��4c����O&��d6	�{JJJ cDʝ����q���=��Q�i�k6��)�T�R�Z �>������� /Rc�ζ��U�������Y+5wY�xس�n�٨���o���(C�$�c�5��q+Z!c�c��G�z���R����(�����6��N{���!�K��d��~Mo�i��װ��N��%J��x4#?��|�!���s3`�à^�$1��yk7R�ˇ.����;I���}�=��5��� �	�АVwo/���x���@�*��S�+4�����q~zh�Cvp�/Oن��G=E��F�~�<��@\W[SS�q*~f��DD��QMG�{�Ѭ������

S���p6���KBE�'=lK��{(����[��9�-�� �mU;�	d�F��F�1$p����� �_V��AܾpҢ���yH�goZ�\}�[��q�ˀ} ��Nץ����ц�5���:B.����M�_3L�ED��{up|�	 j�!���>I`�Ǐ���ƞW�q�hv�����JV�j���35ij��K� L<�����8�� �xJxt�,q�z���]>�ؓ'��G�O�[[T�?�ǒǨX���?�mܞ+w��\��ʭ���:8��rԤ핻̶� ?9�C���u�/ �,��:v㔧��E󥝁N_�G,��,�]6DT#��f��p;��IZ�7����{松<�vt�Q%�@^S���i�E�*~����5jN��M?:�k1��}v�A����� �$}��*B;�־8�A ����S�k���<�����-��/��O���k��S�ߴ�^�r�G���ЗE�ԅ�)+++ �5r����k܋������ӳբ\T�d+�@9H�
P�zf0t��F����L_G�S�Uh]�B�Гƙ/�J�s�0-��5�����ڪ����j�;^h9�Z@+c@�{X ݿ����[)	o��=>?�j���M��"L��Ь����F2��Fس>����vƓRJv�6�WG��͔S�0�\)&��5q(_E���u%D�������]���#<j �n�<��j�;��8|�� �/N�zx��}���;W3���K���J���@��.-�*���)�?���=>tӶNK)�E�0���Rx[��7�/B����;Y(�qu�0�K����I�9�EKn���*�;;lN��n"#�.aD�_��DH@~������a\�k<ˠ96R�Τb[t�ec6��Zݥ��b)���,ؘ��爞��#��Ⱦ6����lbH~�,i�;��.�#c���b��v�9�����K��u�YW#Sz�NuL��Z���]�Z�X%��IMp��1-Io�{J<v�� �@��3��sb���� qi�{j>��»���z�z����_u�u��5Fb��T�e�����{Z�n�oE8�]V�����%:S�=��b�G��k��َJ=|R�Qo'��% �-���50lp�(h���!+d�+���o�;�,�Ea�F,��5�&u��ʵV��us���h��Hh���K�i��6T���f�be�?�(��}=9�̣^Q�H��_�]F����\�Sа�k7�C�Č�6y��Vx��o���n��݆1�>LY�a~�-���5�9Z�[�[,�ޏƽ+�k���-����zJ�z���Y�)4�s�줐_�H�SǙ8�pr���b\�o-���N�є֙�:[=u���|(�C�8f�>J�7 ��f�{��P��~�V��N��bW���6XQp	��j�4�PF���W����!W?�)���\H��n���g{Ned�G�:�v��|;�f�o���1���{���1'��	k�>��M��wn��!B�N��R���é��3��'��9��7����ߍN�������O�5����
S`�cv� q��tg����GE+����Y`�pRM<9�R�C#��g\��v���{]�7�΃�����oՓ�(�{5��Qϭ������OU4���qg���.h����X�i*�t����@ћ�4W;�k��|)�=��ݎpv��Q�`z��0X�x����g��92q�t&���l�q����j��Y� �Kz�#�(�=`Iu��W@��p��ѧ��2@u�m� 	��k�b��(0v�70V�onv^'+�:��R4��I#i�<�{���2;U0��;��un� �s���Qp�vc8���5�����#v��f��f�[���z`�N���,��7��i����D���G���'�@8M`���'el1 co�v��mN2�8�ױE�V��.EB��K�K�����ۤ�T���
���Q��!��~�,��~��j�"�;�t��	w�v�J�QsMA$.����"�R��VU�ų���(���l���gC�/�l�7�{�-7�}��=��
%1
�<(#c�>v������\�����b�VxTT(p�BB���El�II��~����8����{�c7�Ȗ� �
|��ڎ����"���K,��K_�Y�ͨ�Kϸ�+�6���`zi�ll=>�,��HL�}	6��exvt8��;�?���_�<�
�Cx����� ��Jyy������1@��8��9�Y�r#`^'�~ԁ,u3W��4�!\�L �b���p�N��� CK�E�n�ݜ���)�$f����h��f���:l��6��B�Y������k�w6@i�����Q4�xW5l�Y�(_G��[�N3��~��k��VRW!F�u�嫋d����ȼ�h�
HC ���}�~�s�5�v{�:�˵�!v�+ɛ*���\�
[�Ie����=����悢�Xdp�Ѩb��r9;)��Ya����?{{�<];�˸c^�-	���q�k��o>�}��Ɔ@q�%q�Ÿ��h8n4�;��k��:�\"+s�˶��l���Ѯ�jb�NK��ЈAf���W�EԤH�@E���,/�{�Ʈ?ZAR��qR�a8��5Ԇ#ej�jۆ+�6&t�+֋KMt�yo>e�~�,'G��7�q�ϰ��+)ލ{7�8nT::�ۏ�UoR_��o���J���JF}�����.�����l�w�e�]��S랓�4�a��H��Ə�?�'�6���^�����S0��
���%��Ժ�����GE]]�/E*&..;E��ҽ��/_������duvv�P=e���k�x��*s��*����`'�����%�v�&�˘@���m#��g�O?���׸Y[ZZ�o�[Yeݼ5Y�QWZ����u��_�ɓ��W�~IM-��q�S'qN���>Yk�^ML���qNK����������п�$pzق�Q䇆�������}���ӗ�����6���[	$dxh�s�������U�ᡡ��,%`I^QQ�=�73�$UJ��ʯ�8b�g�������X,B�p�#�4����<`�����r5G��1���'K`iN���)o&�� ���Z���JH`��+�Z+i�g��j�ߚ���=��ut�tR��d�[P?a+L%��%c���?�q�� `B���Ϻ��/��p����9�%2f��M9��_�w����m|	D�QD$�0 i�.����i�S��J��a�zh��9<�������uyy͉��^�^k��>��K�o�T+i����,U.)O�'- ���B��5&q���yo~4�y.�~b�2��`p���49���]�����V�� �D�����@X!������ŭM�G�E̯S/�V�vس	ټ�@+�@>޾ ����V����Y���$j���IOp�`耉��{�(:N<��઱�s�nڋ7�$Qֵb�/�'{IL��K���h��#����1��,���S'dS��	�h��^s֕� �!-=���M� !s���S�(�K9�q�3�9�
��$%��K��8�Q���p<䉫뙽�{�㿯P��
��M�|P�8~��V��9C�Dm�
���6��� p��ގ�l6�+�K�
}�"W� t��q]�V��:S����r��$�� 1�����
��(�4C�;gqI׬������eM±�C��-�6{ɑ�nt���@a�p�n|2����e�/�W:"�G�G��nGm}`����E}�!K�CQ��<)�Oŉ�R4	@�eC����t�_�YsP �� X1v��g����4��4���m�_<]���2����7�X��#���;	d�r��=��3,���Ab�=`�i�&=�_0�tF��Ӟ����#s8���w���W!�}H��e�iـU\�ad�o��\�L
���������n�t�Tu_�3�o�jj6�	0��ؿa�����P���z�ю9:��|��C��=�߬KOػ�\&��(�����R�t�����D٤S�OG�WM_�8&��"������30X�7��}�=x�!/,���<�>8!v�ߣ�5YV��GIn0\�`����_W};�L>&%'k:_;_�u�� ~c�l�3d�
��x↺ϧ|L��^��S�&k�&tL� ~O�GLZ�^���E�V'ǟ�/�i�j9��\U
|ۨM�+Р!2 _)�S��o~6��q:�z�Ov�W0�4b������I���2�7 �G�gupQ0�3"d�g�TX�?��$�01�'顥ח����f����̌�8j�K�\jߪ�@<A7�d����8%شY=�?�i�ߢ"������1��;�3Y�D�~E��o? 3;����A�ⷠb�`5���k���.g!���[�e�"�����F"J�2����{�5 �~�Ն#�ϝ >��Js�"�J�x2��_�X�	3�57H�X��޼���=��_��Z �t7tL�"��}�A�@6�Fܺ�^����ë�vp �`�>v5�yG�{M#��#����HӶt�i~>n�$��&ã�X�4xKj�>���o?�ί�V���`��޷�w�d�~ݎgr'"?���-2�ē��C/dF
��߷�Z����4��ǿ(�f��"?��/^sk4� �0��'���l�+̺�Bh��]g����B����?+(��a�o����2
�ƻ��)Y�1oj}����s�P�;�u�g�c�G�H6��x�����ok5X|�]8�%��I���7��?C&��m�_(��$KH�]6�G�2Fn�u ���Q������t=G�)��������$e�ܝ�!��Ϡ;7��R�b}�T�>�@���K�ڷ��@��e�މ*��Eڄ;z�.@�����Y3J����oZ"��b��h�=��E�@����ީI�q�����\��,�{j���1��25�_�:�@�w��ē�s�)�����5�Lֈ:G��+i�ږܐƯ�|���q����a�+[��5@�O �����fr��pl��/e�C���?Zv�]A�v��)�]	���|*=t�uL�/%dF�8�sP����0�K\ ��n;�a���܈�K@��o�t�c�߼�pX�J�"j<��7�,?�F�����uH۱%s�H#챏˭�ٖ��ʐ��t�/^H�1 I�$hX��"��Q���`��!xxH@ '� "]J��ǌ.����-�U�����S@��d��yRU"���(��C�=�
>���y��pxN�$�k[���?/>7ϋ#������dJHc1S߭���Z��@��<t읆�g-�����2ɏ�΋�ݔA�����d7=/ٵ;B??5�9>APC���t�����e'�������d�f��K�n�Y櫓~��m梺'̀2�?`�@��ۆmK?����;�CC"�ݼ�� |`i:�tM�(;`eg�D㼲{#�X��B �1Fu�%�id��������������oͳ���^����Z��`�ą;ڗ�ɀ�z���PIò^ r~����(��m�]�vh�L�N�,���adS��v�)�:��KP���a��z�,�M	�|�B��~R� �pc!��k�-�>��͇bb����
JJ�>>�MMM7o����3����G
��ܶ66jFF����41)\\��`��55�ZZZ9���ǚ~@N�%��(he���E蛍�{�yX)��"�Ui�hE@@��G�����쏄����ԢjU54"srs��qqw �[[k����S�ٹ�##�oJ�9EZ/���]�6�й��q��
�w%PIIɷ��\��,ץ��?������=4�����������t��Z''>�R��$��S���b���z�@��Q�+��@A��$�d�kD��񬣳S�ͭl�3(D��տEG�77��'Ŝf�<�FR��m��Y2r�%�Ӧ�E4�{���{�tk)�c���p��%���l�Y�ϛ�=�,���n-%�ِ۩ee����JDw���\�x�ֺ��圂ll���\�/���d����-a Џw�G�uhS�6f?s�{�Y```PHH��E��-5~�-��B���2 �����	�V���K+�
�B�(o~% +ޮ��[`���������}� h
se[�%��K����I���k�+?�r�=�`�4�sf�^��3�p �;̤@2���8�(���}���@�����K֕7��9���߿_�py�`!����Y��͛�tt##�����{NEEekk���Z���~!0��999
 R��^++���.�\���f�>D%�l�U��ۙ�:ѷ����* �.<���� �VV�_����(�������Y�� ��9����SV�	@�HPu�-�nr�8�V>�l9�ަ�^��Ӆ���z�
�쬟>}���R���Í-0¤� �6|��|��RC]��C�0,�p���L3�Խ��\W��H`�W<�)���k�5���}�|�I�j���S�q�곥�����wAOJ,��󪥵����i��̚�*��f���/������y������t�^]F�S��^6aA�>�K���p/נ���DÉ�Ҡ�H�Kӳhj]�g�pI
/ne*[*��B����n�IG�y��Ԓ򛚛1�V�88`-�ݓږpy�k�{�e��LF8g#���g��[�w`�㬩X�
��c5��r�<X�nUP���u�0�(�q8
(|)?J�p���(C�`0�fWk	���C+>���:`B���M.�hH g��U��U���Fy�.N�7o�}y��J�yn}��,z�{����{=����u��;�d���W��@x�Ǜr����c�� �I��gd�~)�x��u�TGD��|wa�e�<<7V�~�֑8�U������
������x@�����#����(߮}"Mq~�
@[z��Q�V��U*�F)��x����&hb�~���=`T�B���$��z�{������-���p0J�ʥξY����8V  �w��Ia+D��8�n�\�~�O���������h{H {������X<E�__�sl^WP>�c�apN�h�X`뢶������Afp>���c�Σ�����/XT��&i�?�pz��uG�yȩ	=Xow�Qyq�CH�u38	��Ϧ��ut�7F#��k;r��� ª�N�E�Z�TH~v��(�w��p��r�}��|��:�և\���.��5�tFǿ�+'��yI���gꩫ�o����Ift��� 4���]�ub��:���0�"�	 ��
)��6�O�t4I!/`��ـ��R�F��EH�`~=�o6���l���v3������~p�A%��[;�oW��[ÒK�b��$�#� Uza$����Rݒ?�l��5�A7��q��������m����FE:K��g����R8�>U�I��e�� V���DA��d:��M�8䟷�PTa�#�.��}���r�E�:ʞt�	B�	"�Kɒt>��I��i��y�Q?�[�CU�FW��D������*�����9["�tw�X?S?���v!�>�p�1}nmM;��j}�;{�=�������!�N�me��?�F�����Cp�O�|�ᡉ����wD�bf�� 5t0I�Ֆ��2# 	����	�	k=.l�\h�0�O7y��DUkY�X�н�/ x�]�4���p�c�:F�l��z��ߍ%�¼�}R�5hAww�|qQ_Fw.����3мAc�˖������_��p�G��l�!����Э<��F9����*滅r�=�+s;�k���m!��?��l�C7�d'��L�$��A��c^8�p(^J@/���sFO�dg��������|F�`��@~�u}�f�⤎�f�D��-���Y���3pI݆�ͪ�e'�qt0dM�~�����L�v���۾�����Z����A�Q�y�d���[cj�����@ D�k��݊�0r�-8ϫ�I't�Wn��n���'�ϕ2�Y��
Ȩ��	nTH3Z��.��n�M�T�b&|Y:.�#̓��+��*e�5�@i�ޝ˼����)Y%~I��vb��2(�Dl��$�*���#�]�h�oӧ�P�by+���j�P.X<X�i �����z�a<��_ߎu��}e�������h�NǕdO��}�NdaE��ut.���j4X�l���{�!�T�#�%�6�#R�S�uR�m���ߢ��Pr[!�W�%�x�(W�����<�l@��Y�c�]i��=�����@��״iAM�޴�CL­OG>^��k���Խ�_���} �gZ:et��9Q0�uH���r���⦊�w0� �:�� Ԛp��R^�H��}&�d�Vu��}��C�%«�F�v��5=f�,4�D���l�'����`�˦Z�ҫ��7A�Gq]�.�ZfB�����\\ܲ6��
�A����"~��M�䋎�c�/���ZP���Aq������;q�ZFؼ��K�5�s�~<K���Q.�3�q^ϩP��)^荠b�F��5�.� g'20S��Z��[�%�(�������	&06��G�� ��7����?��1��?��v{�~��y�JM��eЁ�ː����3X����K��.�������HɈ�{ZړY��ژ!��M��Za��{��Q�T��h�Z�ې��������S��v 
;�HkH0��^O�;_X�����m/�Bݾ���1��O��A+�[���PYG84�J�ʛ�?Ƚ@�nbS+���}��sY�3tO��'H���S�>��9��7���9����;b�l�:C_p{ו伸[���UNŝ��0�[�1�U?�]L'�E��#�G�e��P-����H�Ad�e��l�jᒇ"����p��:I�Jm{�ʬ��[��e��j���Su+�퇈���-'�d9�Ky��>#�X-/-�e���4')�ig��sa:&�i#\��2Pq���Z�<��!*��m�1 s�Œ�M"-+B�Oo<���/�����_տ�[�!�Ki�� ��)3E8xN�G�Q�{8���j	�œˣ5No*dwW ��[8
��B��U��0���c_���Թ{-��$u�5�3fi�S8pdtK���%%����T�֬|����Qf��B;t��E���@������Þ/�L�y���s�DhAp+�Z��+�N�w������Ҭ(�*��t���jݱ���ͻ[&b)�kmAa���N��"R�,��ԧ�wc�M��+9`2L��2�� KU�<ۡwۈ[�"YYyώi�m}˅�tlt�B��w&O0���N�o��j�L��r~�[�O�k�����=�4JN��?h�%
ݼ�>��W��T��{k�c��Q��E?I����A�:�����Q<� f7(�F�w��N</$,�H}:`��	>Z�z�D��ƪh�"�8m^['/NI
�ɤ�veY����6n�pG�[&�N�{�;.m�'� J�_0g~�r�����S¼=�c��3F�*�}��y��x�B�bQ���o�o�T:��N���%�T2Cqk�ސ�.nC��L���q���͡'a�B8�Q��i^�g&�-KX�`�m�)�tG&�g��r�vL=��)n��}t�%<H��UM����1�}f�����O�c�=�z�U,��y=���2�t�c�H�8���ʜW������ƽ )�sE�$��;M��͜w�(���v[�o�}R�²P�ʷ��$��Em@�����_9��d�M����7�FC�>�j���{�z���'KH]~�>^��Z�kӱmoU�-������*γ���U1<017l���ڻa?,;��y�z}W�A|��"����S늿:+u�ۄ�d[6-��lx%(hS��o�76�~1#Kxy⮬����毳X8/ȚO����%�����}�B��A����᪕�'w�n���j�,(T0��ws�SuW&P,�BV�_�r�P�/�c��2�$X}�\�=��K��:V������U�2���=��2�@DdP�HD^�����B:��ó�S-�X'�eI�M��7�O�(���<ZRn��.g����b��6\��oj��|����\��X���T�Y����Y�>߹?ɛY7`\ĳa�"cg�0b�֯t4��N�ϡ���=%�ӲJ�:Q#lB�@�;u��/����� g����.� 
������S졫��rQ�����N�M��.�죝���Pc��e���y"U	��<�� ���+~�eJ:#Q�x�����%�[��$����y�{_��O�h���i�;�C�;m"���.���To�YM.0a?Z~r���"����w�(;�����h�5�7��t>3�nZK�oa�)H�>�z����Db��a0f�'gY[��� _�G�%�N��k$WY|���T;Es⑈������D�3U�����ವ�ÒX=�
����9H�WL8`�a�<I�aky�����k�t&n����vx��a����B<+�ڣ�~�ཕ�J�Ulo�po�a6%���dh��q�z�K�[�8�GI�R��ċ�䤴����Z#\y(�Ai8�ja��Xh�V�����a��NA<	����Z -_�Okn��I��.D9.�=�8mZ��I�D��jNS�����GVa�V��S�Qu��k��q�$_LE�Ť'�3'��gr�Ze�'n�+V�������23xz���bD�$a �mLШ�0&���q̷�N��C@sRw6�W3S���R�7)��읉�xf�?~�TP�t�O�5���*�y�uqX��l��f}�ki��uW���M1��u<a���͏&�&� �hyPn���>�ʎ!��[Ϫ�Sn����^8ng�X~	^������@��6&7�!�f"��>�?��ݝ�W�H���T;1&�m�5����K���w�̎8v!�ʜ�z���kAaW4l���h{$"���躛��K��b51��Lu^ZN,���)��
Ԛ�II u��~�;�Uq�ʲB��d�|S=K8��6�l��R�����4"4}��-�;u�w-�aJ4��F9.΀pv�~�(;�И�a.`F�"��X&��נPj}���j#E���2�j͏���R(Qf��4�d1/�0��^!:�����;b	"�����E�s[F����RAIP��LX����=l��|�2���&���C!�����!��ä��?��w���h{k�b��ȧ�0l��2��݁��#��[��ܺn?�e���;�
H#�F�\[��t�57
e׏�r�N�sج֫땣*��[�*��_g]/���w z�p:�`�w��������b�m�*��y�˅3+�����@w6���_/WF,�*g��I�μ��������o��{?k��l()3D�~�U�x���)6��[m&<����H�M=ZZ����\@��& ��I�ث!���V���.�-�[n!���+��a��O��Qi�a�X/���A{=߁��G�ng�K4V?��/8�F��n&���Օ�u]�ɚ����BTYE�[K<j�b�|��:Jd8�y�Ny$,�� y��#��2w���V�.7g��
]�S�z�)���Rw�������'�m����g�TM,<>�o7��a�\[;s	;����;���m�����cE�9������r�@�-Bo�+܋rԈq�/PǞh��C�O7�+5.�N��{e4�G�빍&�ˈ�u��j[�)�;*�����pv���㈡�O � T�?�|�3�0��*T��p�H�%Kr���i�ڣ��?����|��eǉ��O ����5|$̅���Ś\%଴y�l��h�%D����h��~^��>��]�%�$�*��?�є{�5g�a;�şIH0��|	��Af���m�Jy��Q8�ZV�!��=�ul�x�V�8�������Yn5Y�
����b�e�W!r�aT�~����=WN�[�q�+Vb�I2Ƽ::���Ө�`At���_g0K(Qϸ+���V��!���,*�I(A�0�t¶� P#}�ugk���T}�����������7�)a�}�߽W���ב��K]����y{{J�!)`�(��V�+�C��𙬫�����}�)�hP���������q-�n>:rBdu����H�̐�!�)޳W-��jN�-���T#Vs뢤~O�gLMd�D��&��K���B� �6�q�:>4�;İ(6W�<�	(��w���-M���"�Ǳj}h��Y����A}qFÐ�~�js!��q��XW%�� >Wk�/2��a\����`t�Ms�#7�����)P&��D�ʰ��3���&����
�vo���i媢�:���*���֐�/w�R�q9�# N�K�[c�����U���L�� �E,���qn� �[Q�5��)��A@�����n^0� �ɽV��fOe��c����	�=�J��L�jm��0}��Ѡ����2̵�~4�ZПA~۲�&1�j�{5zac��}�d%>�ԡ���W��m��w�E�t�#��I��F	R	�~a~���,�^�>�2G�`���()7�cذW��*&��c:Ʃ��&�/(��`��"����X��+�6���W",f$=S�L��m�%�Q�B�n��z�{��������ӱ�W5�Nw2����UÍ��b��GN�Ύx��� wm�qk���F��q�L\ym�<JU��=�.�)�;��V3�tr�1��p��+��aW��m=bQ�˺��5&���M.W_��4��&��a�lMF��ᯀ�XP��*hX�B;� 6����laQ�t���Pj�.�$�_<��D�L��Ə55�5=�f�U�ackrk;���(mPn�P1�"�]՗���wKHY�N�<� �;ij���x'�{����4���"�,���v�DϢx"�ӛ���: C���2Qy2{��ŉΕ��x̃g�*Hζ���U#8BU�ͷ�:�簹RRY���FM��雤ᵬ�tocc��z��[nk�'e���.ar�Q����J=qtg���	3&7����p`a0��mS���
�8۱��XຉS�IL�5�CM�GU�lp�݇R�8]������?mV �Sf��NC�Y�'���J_r�����~���>��y���e_�S坚���:P�66�����tL~|�Q�TCe��V�W3�¯�:b�y	H�f��ĩ����o����O��[��$R	�D��˘�=EW�c]��Vݹ��/ ���.�՘���k1xԄSc�ѻ4J����G%�9傆��� ,wry��`������kў�5����3f*���IĨ�*�� v7��Oz���=#O2Re�R���#��a_o�3ޞ�t"����� �^)�U�&&��,M���[�.JR�;h��T�o��Y�;���sO]_��O����5ze�%.��	`^��+� �������wi�U�e5M���>:I���cω�gWn=�V���H)|Z�]"G�^�?{62:g�c4p�$G�Z�h���~�o�f��s3�F$cS����K�#���R��E�	ן���x�Ua˸fd5�σ��Ϊ���1e�ռ`�n�&��ȓ�Q�
�7T��u�w���6����ϝ���k&*Ğ��,1�syiA�����Ȭ=[ܘ��[��0�r&��g{��<���:���/�K�kZQu+>�p�~V~��<ݫ�P��k�'�j=$IA�[�A�$���w�\��o2}J�xb'�(w@���^�%�W@��I��T �$mm��DN
��v&ՙĢǝ�\<	�4}�4���qf?�y��i����G]�Xn"�n4};��\H������J9�f95�~r�X7��u��pԙjJ~��  ݼN�)�-��zqX���֯�3�E90����c�s�=�gC.aW��\�k� W���4���^D�Ol��M�ڍ��\��3(�3R���D��?q�op��.uJ���t��k/�?J��z�~����竛>D 罉�k��b��"��s]vm�ɴ�z����v��U�����
��/V�d�x��藐3Y�i�iq������͕����?�T_
YX�u&p.ʮ:�b��
ť�~� �{[�-b:-h/�� Z��`U�!Ϡ�0v@�0�Ԣ���1�b���|�AsҶf5�`yG����}�rqx0��V(b���P�4FB��U �w`��|�J��w���eFu2�"8b����&v��[ޖ��~翣�o�E��>�-�Vޘ};�@d�=d;�훅�(�����L��限�k�e:xvv�Y�a��o�.��K�4^Ik�-��tM��`p�x?��۹�̼?�e?Mz0'?��=��n����*�g''�%W�OP���	���=g�}j�H����$��x�e/�FN6�vHoP��|1N��$�BJ�X��>k�47Z��C������H�(}����șݒQ��K�9�ӯ�C����� ���x�==o��&Y�Y�.�����Ź�I%�p��:nI{��&���E�G���S�[�2��o��k�/x����a7=��7�ҒJ���ɸ�����3���M��c�PbV��0i�#���l.����������
2�g���I���\�Y����p?P��P���x/����� ��C:�癋���冀jÌ=j§X�Z��# *�0ܯ]�S�9����ZE���O���rj�|M��ok��U�n��;t<�!����[B�����תz[�CP��`[�?�9�{[T��ݔ���Hb#6�;Y�GCm�me�g�h���٘��٘3\<�-�[eP�Ƹeߴ��ZC|ʧ�mCGN�W�LV���$̾e��^,7%�4�+�O�۷nq0J�s���P�~?Vq?��gB��]����|��}�4Tw�Y<朙�|��/�85�~g��L��/�:��</KP�PxO�f,z��ܢ��khs.uO( X~��s��T�����z��Ε�F��b�4�\���GZ#>�w.ŭ�R>�]Ȥ%_�$%֯6�����Q���OO�%P,o��_#c��6<�f�T�9��m竔��������P�r�(�0΍��x���:vw��Q���`������ݡ��u+	��	�d� #��BV�)�6�IDl�*K����%ag7G�j�����%�D5Ɵ�?Œ�^���H�^ѳ���M�����:u[��@����=�a
���by�0��� K�m/n4O��ϞU[֤T�|�\|�#έ+�� ��"���5���nW�se$h�U*KJ�bх]�0k[�\h�oa:���nM��@����V-��Qi��c���Ɇ��|Vj�l5AU�ئ��`�n�g��l�mߊ�����9qdK����9Z�%7�_�6�J��:�|Ҷp0} p�8�'��F�%�����<9BB�&T(�$�)^R<3��,��Ry,M�d��妎��)�/������u��i;p�v<x��������eܐy��"4����uܞ)2F�j	ƎONw����^�&���Y45t�o��eL56���FwI5��oF���Z~�]�}]�.��gY�bq�0�1��6f�[�|����^���Ԛ��8�����.����qn�	sC+���[,�),��m�����������u��)3�h�W�мSc�ҳS�ҫ�GM]y:#��Q"���؞��;q�qK�32�&���S8�Ue^F�
���{|��] ��9�Y*��7mq�`�hZ�����Qu��L����W��\|�^%i���7�k����I�بL���۴�e����2�6�W��������-"�N�J߈{/7�2n��/�E �oC��6��.؏��A�.��H�E P5 a�EL�%Rhz����#�>?�U�ꮩ/���;����|~���d�t�����vN����Vm+��*���ּ-Ee�ZW�f��T���.Ƭ�o
a��bjd��V�+ ~�bJ�ӎ��/�x*'K�����opm�p��r�'a������S�q��]e�\���:�)��ũ�WBW�>�nv����P6u�O�ch��lø���p<|$P0����������1�Шid_��0���z�� ������vѻ�\+�=K���2�EWĬ��J"xb� +�ΨG
��$��m�Kiv�UM����nUڏ�{.~��P���W�=K��;�@�o��dJ��XS�+�x1��T(ٵ�"���~��� ��� ��B�g�}l�'v�������x�S���t�V����Ң�!jjm��x����m&&��nů�g]>�䝧���<���e�<�����D��L'���s�l�����O�p�����]�!�TL+z~��a+����#�4�-�QE}����#�Q�7�e�4}��bLi]�~/r��L�έj�:���
4��%�ђ��'=���j7[��G�J� 5�Ds���5�m~wF�@?�r
(���՝a��v�̵JEK��׭��7�ݑ�̂	^�;���ڡRN��Hl�K����5�i2�L����U:����L(��XN�OZ(Q����ː�=��c�����*_�g��EHU�b*J�0�Gxg������D��Y�k)�R�^��G��V�K���f���a����1P|dP��.>���uQ?��tcUT�Vm�Kx��N��|�����`������]���b�f�%�1��R3�@��Ȅm�������<��`6������c��@�J:2�]���u���D"F|��$�`̡qP���Nwkŗ\@�,'���%6�P�e�q�]�X� OL�}�7k+�P�<έú���o��(��������Yq�R-p����/�<�� ��'vbri?��x4�@��o��`v��I�s���{{&��5}��m��&��U�}x}v�'��WNv5�_8����)�ÎJ��q6I�C��C�OՆA|���XK;��>��ȍE���A�@�3Tȹ�#%�>M�_E`Q X��۩?>ѕԭR�%�����?Ҳ�i��`svӢ�˸HI���R�zm,��c����Stl"t�w�q(�$\[��7���a���~�3��ԍ�Ѻ)��Ӻ��Ű�x�����mO²���)���m���uVѪ�i�2bĉ3U��6�
d��.*ìW����Z�Jw*�#��%�M@F��%��?a����X���3K���i���I�F)�$
�����2\U�fv�2���ŕ��;��P{Ov���)A�?����� �_>���s,��ZC����˖����Ш��8�O�ӝ+�n5��;���=��ե���cGg%��wY��)��. �#���*�e�.5x�-H;хY�-��`���黴1�藈���>̇��+�|EU�Z~x�,��gIfA>�j�BV�#�k���)ҭ!}��/� �XC�Q_��SV6���B�5��S��b�k��qޖg����;�r�S�/�߻Ez�k�J8���0����}#�[Ju;�H]T������l�^W~���.I%����r��+9P�G�D���1������q!���b������o�@f��^���5�$Y]BtvA��&�>e�."�,�Mi�2?��6���v���nV�}�*�9��ȭ��2�������cL��I`����� 
�|���Z1�M(�=:��]�Y���?��2v�W?����^�U���y����-b=E�_�5��ԉ�{�J���8{��ԉK�B)(���ҹ�P���P E+�>����8�)�W��W5�����`�Gz�(�(�(kc�45��F�h~�ñ/54\B��ϰ��R�u5�c|��	O���G]r�Z��.������l�+�s�yV6�.,���W��iVO�W"��9��e�:Y�;3���:�1�y�e,,�@"d�&g�F݌��K���YgKZ��.!.@z;��fd| �?�5�|�32 aϳ����nc�����گ�E�Y����IX�ͨt��
����RwJߥW�{s,�w��غ�vW�*��a2m��!sܜ1��M��4���Ф�(>�D��?�k���(��7(�j}������Y��+��m^�����½��O4���)CE�`f�e�6��\��a�%���`���>ބo�#D�@叨[	uw�x)o`�Mo<�<9�Ӂ��&���Ė��ڕ����y,R�$i��mj!�G�x����HN���TU��?��?�R'����9R$cUe{'w�+�ikg�ë��wK2i��m�NǾ���ѫ���U�:	�1݆&��t�޲	�uV~�l��U
��:z�bFo��<�����NV�����X��ۛ��H��f��'禎�&����L߾b�*�E����z�,�����g3?����BJ4,nkh����8R<�Q���੤���cm}�+�~�߀��5軝ޯumN�]��G����}/¯!%��.����I	�b�yq����ZܡB�o��s��i��i�_R���ٻa;�3�}��:~v5vt���Z��Іa�h��C��4����%�a« ������3�rN/z}�D��!GI!ʃ�����rH����������
�^i�VU�����-�M`=�{�8;��ǀj�{d��8/�4G܉��,n�IEz4��P��㩾��qB:�G;=��k��D��O�ܧa�t���xem%m�ۦ���Q䬾�p���v4�e����S$"EΤ��-�t��>�
��������nZ�O��
��Ͳë_��<��~���K��s^K,--u���� �	�{�k�6hLi�x��v?p�n/_C�!;�/�����n#^�o!,�{<}Vc��z++	K��$���4�TZ��;�q8�"��=�d4ko�F���N�ryݷ�&�$����='��00�{de�q��8-��5sD!���<�o�QY´{[���N�5sr�����Qo.������h�0��hr5r��(��g����I�\*-����9����bn�D!c����^��I0*u�"ȧh|�z~wj�d�D���j��F4JRg���`�������ڛW�e������9�a���m�9���0�2�
I���k?����MF"�c�	�Y���
��Bɺ��.o���^3�<�����X���f�]��U	e�e�`�+K�ML4t���/��:9�H�0�Y_;�P~�m0T>~|Z�����O�0��J��L>�ߗ���:�V��r	*[x�a�N�x�ҭ��^F1�D-I�g�v�wPۍ�7c������&E�l�GI� �����'	U'=�(�yY�G�񯌧<���
����+��nw?A�g�z�_�X�]�@��nHiz��5�����t���|ݚ��/o�.�3��/���Jހv��.п�hTg)�Z
R�`�r��mB���"�/k��,���������p/�V�؂���9�W��(��R���%T[з~>���җ~ro.b�[���K�;gyi?3��8�LSM����|�xy{�e����k�'U����g� ��Yyuo�]�qÌV�T-N��x�D�F�[��쾯la~�PE��$�GM���!0�R7&y�U������EJgb[���.����v9Hxb���-)U��q��l���\�[�.�ra�G֙��5�\$ ���n�G���<����$���6�{jg:�5��S
�ʍRtԍXq�dٵ�$�˅���C��*"3���Պ;9��D.Q=l�D�quN�L��|&ֻ��b�y\Q@��Mi��lHɸY�Xۃ-��4j����p*�=|�Y��G޻yK��)V.�۰�AR���my(�$uf'��5�{0R�H�-IV�iL���<�}�&<��������z5�k�߽[�~-��32�G����t���f~njx���P��>w鍋�o'�z�(��n����|�$Ol���%�2������σ����cU��d�X�K�/��R�쉎���iԖ�.��DdpL���t�c�e%Ʃ�H�|�ϳ�F��no���A�:��=x��qݖ�EE�z��eT~S�a�̘i}���]5�|���t�\Ɣ�O���X��}�}ʷc����:mQ�T:&K�x�����m�Q��6Ḏ��s�c6*��`�[���S�ϵiZ���@����Tm��R�.�(L�!���^B[�gH��s���H��iw�uc�-�羾�����;s�3��V{��;S�c@;}��Z����ּA�X�.�I��o�FԼk��7�i[g	�f��Jh���ĄE��d�,�'I�d�հ�_k3t�����[���W%��;Ex�hQs��J�)��b��z�{��Vm#w���8������j�k�EADTDz��� ґ&M:(� =tED�w�  �K�J�z��A�� ��~��y�{��뮳�y�Yg=�d�=3{����|a�7���~$'s]ݤ���L�&&Jq03/荢�y�$����u����//�1����7>��o��� a��p��O����~	2�lz�V�Fw�lQ��|��w7���wS���� �9M�Θf�gL��ظ��v�o���,�h�rS������_{�������$f�}�O�������
��A����|��y��o���
��]��I��_���(!�_��_{���r���4;I��h�P&�(g���,w��;�kͶ��0���������������h!�"�qXm��s�:�DA�	P�A[���*�6�z�Y�d&��Z��vHV9HwaO����L�V��M'��Dd�P��������%6���?��9q̾�n�_�f4z���a-����{Nu��-��.�)jvҜA����'Ѿ@r�]6�I�
��8�ļ�4Z-׶� �F��B�S���5���X��ώ�?�s��KOe�۹�-_�v�0���=�8��4'�H!�$.����X�םD�>Y�������ڶ�1h.��is-ܮ%�JN�N�q�A|��i��@���&6oS<L����$���M�nt�/�l��b�����V�N:��]N��hc�y w5�+(ݭ`�$ݺ�h��xK���բ�!u�;2t��OZ�sy�(�"da�!}���cL&�>u�+�7���#kmAwj9]�Uj�� .��-'Ò	yzH0�'�{�9�ys��o�B���zo,e.w��p,�w|�t^������||S'p9h+��C�>�l�&�]��o���+Jڕn�ӈl�D	L��ܮ��ۗ��>���Tw��6�ҦE����Hc�H|�ď�El�r+!Zm(��4���r�tr2z�(���~�9�J{�S�TT��h�m�/6M�L��@D=a,�"ڲ"���K���A��R�kVC�	�M}��9Ri��"����Ɗ��sX:��/�6�(dbׂe��b���_J����qW,dۂ�X̛�509��ONux��|g�O5œ2�T�v\���u�z�}?fՆ�]��N�f�2��-
:����^��w��Y��$����.7�\_�*�Y^�,�u��
W|� a[ �q�n��eǞ�^YV��s��1b��zBW@�F��.s�����5,�|*m��=���-p�ԓ1R�o�^}���%�C�?C{����^�loj�Pgp�এOyľE�����4{�9_�B��Tk*�E������Mv�W/��iq�F� ��r*��N[j��b؀ü����|A�kB� ���G�?S�|�e��œ�c������No���i����X��2'��ʍ:MÂ�B�9��m�_K�?a�w�q�I�BJ�`���ef8n#�7��-G"�ࠢ����I�4f��d���mp���U/�5����ѡ��yD2i�}���c�����ծ-3�)����W�O����Ӟ�Ԇ�r��-�ѷ��Zt�n#��#(�w���KLn:��;�p��Je���y��0�1���'p�@�JC���F���ߟ����ڗ��wA�J�{�`��Ok�N]�bTv��<b��R�i��o�*ܼ�mX�kx���b
��ݖ[�3k�y�U4���y~)(�`�LvI�0Am�ϊkG]Y��:�56.bKġ�V��7?��ˉ�mN��u]�Y� �X�-#� ����>Pt�:Nb�����;9 ��G�u�1�uv̢��۶�,�z�8�|���L��U?%0����]ur�S���H:�t��Wٷ��f���,�V�K�"s%,!�G��?~��S��@}�$������,�yp�����Q
�$�P{Q]m�4�DSǱ�0�̧��!9�
m�B�sw���;�a-�͋!T��f2���4�_0��hE��ۮ� �W��4dA�?� ��x�ϝ�H���t
n �~7�.���[@�2mOM}_��hɤB�B`�#�����vЋ��<b�`��� L�p<;����i�9�#����;�������w�/.��B��}�	g[i���v��.���� �*��<��l%�_�^�9n�>;�E�q�7�*���H��~�x���?ֳ&Su��oT��vu��=��2�=�	j�
~A��w_DިŰ�r�Ѥ�� )�z/��Xu��B���A[4K8�V�J��b���DU�枆�a�\�.O/tZS�>��++܊��rvry3$^�]�,z}'S�Զ`�v�ר>\��u��51������mo�|�����v\gpZ#����l�NON�L��f�+�t�F8�OE�6�"n�t�{Z/����	ڬ ��	�*�(��x�zT����~�>�]pϿ����h�c���К�@e�E:U��X���o�6�E�X��@e]��_������<�=L7A���[���<V��^���n	��5V,��Y����:�`���:In�8�(��ߓ{��<K|��km�h�Yۆ��gXk���3J=���Cu;f�n���w'�Jz� H�u�pM�]Lѡ6���
�XR���i�����5��k���L���4�0b��1�V.��d1=}r-�8X}:N�#w�;2g���U6�.�S�ɞ�թ��T*�w�B�������'��>��fղ�C���@]�M���(�i���3K �����/��CS���a���B^�E��fTv����諾�xo=|���]|H��������:x}Y���=����M	�2����7MU'.�.�e�jh�
F ^�L�Ц�دx������;�K�o�[ ��c���H 7��.�5�SH���h~�uB��S{N��Zt`5�c��չB;h^����^#��[��./7
QC��Y���+-��]ߎV��6O,XԬ�� iWγjU,œ����t�C>���y}���8��q:^�F�\�?�v�	IE���PYiC-~���A����+��:�N�~c��'0J�Y�x�o%�Z\�9̽��1��}e[��he�}R�U/١�~\+�'%��~;>����0%;�~,�Yb�C�j�?㐗5���(�Ľ䴛�Q����QAW��ÌŔ~n��Sr�������sE��u
|�JM���e�t5��k}�a\�o&s|�273N�����Z�c�{�x��o�7�� ����-@���7n;�s��W�����gG-V�OQ�,&�^~U�փCլ�(���s��n����B�:�A�9�,{�tC�NѿZIJ6��d.d�G-��;�f谗{W�\gX�h7E�%������)�W�v�Q�m����UVG�e7�r��p})5�5%�Z������
|P>~�p��j�r��w�|A�.Y���j���^���2�w�7�fy��HӏX�@����#{�)�7���	�|�R5OM�Q��Ng�Q��q�"U�KO1�u��gp�]߲-����
�95Կf|b�Y>3z?� ��@k���v,f<�kU�;��r��./�ѿ�&tX� :�WT��o��s�y6v>����_�	V�9������̫A{��c��t�2��oo�I���*�7p��}���D�vH�74[ke�|l�Ȓ��^�C����1�z*�ZZ�Z�i���D�+���UiB��t����{����=9M/��p��w�r�ݰ�ʹ���V�=�,mb��.��x+����|�߆�.3MB�, ���{��,�H�8p���n����j�=]_ϭXY��-ǾƂ�.�����4�U��Jl�����%M�=�> ��2�λe&2-���2�^��֖=x۟������lPp������֗Ƈ�l��f����KEϝ�k��Bq��nX�֤��[��#�����V��0t�-���=��0��l ���Ŏv��24�Ő�uH�Q����RpT�Ά=�^&��7W,�<``��Z�_agu���m�d�^�&��r�]�ԊA5�`�tL|/Zˬ�jh�.�V���=����"ٹ(s�1��~8UN7�I�F��As4s��LKK��Gi9��'~8$U �RJ�37��ޡ�j�c��nD';k�!��{��C�Ld�n�ea�Om���t6Q��4�qU�;ז����ܿ#ܰ��g�~��~�t�!��XX;%��Ŝ"��,P�)Q�{��i�6\s=�����B/x�a;Z���375u�c��w\�_�\���`�g��rV���k߂�6�b�/�|`'����Ci�\����ʓ�ƻ����;]�5�V��ep�(B�+�����M$?�b(;�,[�w_׽��N���^����H�J���W�V׳���!+�2qϣ5����:��dյ�Y*�Y�=�14��nĵ�)��OJ�����'��$aH=l��%��כv��i�/�&��5?�\������WZ0"Pq��=6�uN�Z����u�*h�OQ^��, =^�L�>im���� Q 8�9���κ�O3HYO���7|��t�a��j��X\���j�!ϵ��=�i�����6��F�M��<�ʿ����n���(����4�YwP�r�iNY��d:����ux�T�(x^n5}�U�@]2M�B���q�I����e��63u<�{~��S9�ӒX�b�#��(;R��d2!ǐ����ި���3,�.��م:/@�-��8����7�'�F/pnXf�3t�	Uj��Yչʝ�ߔ�R`��U1[y�OX-��]�6C;��C�~�
}vW��<{_{uZ<���e0��!.g�ȮOv1�ׄ��F�J7��^�Uߊf�;�:�y=���٫��(/s�7�`l�ݔ�^��t���M�*@���X������͍2G�K�XaԘ>O��w] ���d��q>�-,�����қ�:��,F3�Y��AGc��KL@�^�Y��{�������e�}`�[`N�>����Q�6zԯ�8�GI�S��3�-m=}g���iw� G�t�S�rl�'k���UK����`�hK���~l�'���%΍km��r���� ���H��ZjcA� ���w<~�ڡ/�}}�{�&r �G�8�b�@=+��U�͏(~T�O��Uo�	�T4p;����8F���$1'O+��5�v7��jP�j��2��ּ��99F��E�~D�a���$�-Y[��{m��Y�[U>�:~�b6J��w�=�j�8;V�k6p�kp�e�s����Or6`�X�\}Q��m�KD�q�m��3bE�5w��p||k�(��(���"w����𱱱7!�B�I���=����	�r�-�U�w�x���{�h � A�E��D�Ԑ�{f���=W�� z�7��g{��:��
ϸΏ��~���o�[t����;��� x�����eXk����?�}���ǩ�̅.�4��0#ǝa���}9�0 �Z�*.*��]��l~@ 2s��v"N�TK�m�wZM�J��r�ӆ��8=��P�)�j�|�������B���2���JQ3�h�M�py��z�:c�ֈ���ߏ�o�Hi���<�z�a�^h�P�9z6�E�q�	^!	���Ψ�Z~�
*Y�\���w��̄��o���c��k1SUX�ز�Y�!�:Hm�q���p��/�!:N"w�Q���g_��ύ���hq�}�Y��G1;3��;Ӂ�j��`���7W�v/"��3�L`�F5�ا������
�D��O3�G1=~6��Q��7�T3��a�`����$��&�� �#E�C`���Q�Lq��k`�R@3S�#Q[�bSK1S\*�z�@��C2԰+ υFABY���񫻏l�@�a�����f�ftW�acՊJn}�fhթ�H��=���I|� (� ��aX�P^�0 �m�����o9n���D��u�1/�<j��I�����z�%�V7���:�1�Ěf�s'j���$QϬ���G4� �Û���b��ߺK�ܸ�%�~9[��h� ��fc��L�w��gv������cY��L;Ǐj4����;GA��b�i�l��'ˈ�M�}��?cL#M֔[$�8cibv�'�gy���L'z��^�ym��Z�@�k։�J7��"=��`l��ҽ_��5�����(`6���$ã,���t�"�c��g����gE��p�� 7y���؉�j�~Uñ��;z���H�g��� �6P7gY4~�3X~�UI�K'w���5��/���S"���Ǿ��9ja��TN��k�Ǒp�ø&�y��EI�\�	Z���5rg���X5Q@��:����x�kܖX���5sgI �3~��G/��s ��YB��s�@��7�R�����@?���a�d�gܘ;X8�w�G	{�v;��:⏍Q�r�����?CՊ�o���8�m��7���?�Պ,o=���x^-�Mf՟�6%�H����E�(XH쨳
��d�� 6��yuJ�U�T����g��F�2�S�/p'�� P	�%hY '4Q����8Xv��Q=NC�enɧcU`_z��u~VJ��Q"
*Lq�#����� [!j��7@>���Y����s�6`�+$Ӈd�KEp�b����H����\�J���?�S��/�q�L�q,v��n�Gx�+� RE��pRɏ8 )���7B,=��}zOp�Ǹ(�WO�1>HԆ��׊���$���G�
,.$ضp��	8Nl_�^�F���Xg���F�o_�q�e�u�e�t����+ ���Dg酡��0EY��-c�����-ͅϵi���]r��&������&��Ƀ[='s��.�·z���ݎ�PZ� ��o�П	m�y���h?��͏T9���OF ��ӎUz��ߥ�х��;��&��U{�Q���������?�[Z?��D��)|��tc*a�7]�Wx�Ys�\��k�w~o���ُ����F{�H��|��]�I�����w�2�a�W����.��@w$���he��������ii������ִ�?����Ky���\����?��ySȰ�!.�&�lP��F�i��{_�|y'M���פ�+^�A�S�$ݰz��𖻧������?���KM�E����A0��n$j��W�y)�
��f}Q���7����4Βd��X�v<d�u��۝����&�4�Y
&d�4ls�'�b��E3���B���(�Uh!%��#5P�e��|�z��kg��5�Zc7�Fө�T��| ��>���iy����D8	5�m�)��_�Cֱ��!:�æ��OҘ������846W���3g�΍��V��L��2�X�f'�⽨�}�~�ڸgw��"�r�<fhT��[���UA�g/������>�����
�"�������km�+/�!fflI�8;��@@�ҭ��N�QL"n/�7��e����$$������Gj;������m|��7�͍�())	>���T62�	�6�7�F���x^��z���� -��S�잌���o�a^3:�Yk@v��dL���ʗ[2�ƶ�΍��'�������~�5��wu4����C�G�k|w=C,C�TF�g=��D�E��\6D�o;��3�2��t�}ifd~�`�f^��४�ak��a����e���̢a�~r��>D��$��Û�̄R$�Q��u�E�B�j�[�������{|���1�\�}�b+�
z�E��S
zP9[_�R
���k�ke�o}�U����o��|����y9bOd�_cH���В���q�At ��TM��yO���{F]��0���G0^��/��B���o�NQy!�gG��rҨ.v�̸��c3��l
K�3>�s����;;4r�ˮ&0�����[J�U�sB\bNt��*^��|h�?:0�}Q}��ȇ��3��Z7�ZE�IG��B۫@�c4f�Ρϧr�AT��� �A{n!h=WM>>^#�����h�%����qZjnp��6����anB{���eƕ�k�x|�:7T�)��C�\�T+����-�3����h=d&(�I��o�j�p�������U�#z.�Cf|�Rc� ����c�V駫�|W.�ow���)jTu	̬=e��5����+��X ^+TīJ�x�Ljw� R$�>���ܶ�x�_s'�)PI�2�J�?d�v������p�/�]�!Ը	-#�t�>R�{�}4��N�qد���"������DfV�����NK+'����|������@ �xt��A�`r��9�"5ī�a�v��wf* ����ڔ Z��_������$��+"�6����G`�읧�&�,��JR�E	I�p� 5@@&�X�E�`�$��e{��WO�'�	���;�F�Q
��LN̔0X�gG�&�d���q�t����&JT8g��@����&w��E�z6��� ����%g�>Y)�_��j՜�Z�z$�k��'j�h�U%�?�ęɽH�(2d�o_��#�`�R��T��]zG� �<��P����T�WT�z��"x��fΨ�9�������H���$[$yFxN��v`h����M{�~}�e Η��Y�>��c͂�"�^�|���"����kJR��)ba$�O�N�/E���[(�w�؊	e���6Q��g���_%I���) ���_z��_:k�_�{�"�y�b�GYן�����p��:�8���"=�>���b�@���k�������8�	�5�H#�M-<�rP�)���c(�^�)2H9;��2;��7U�
L��K�c���6*�4/��<����p!rc����ht��#q����L-2|iP����g��6�Fz����%��^c�OLU�_�_���3?�f�ď��ϯ������7˸K�%�����z=���]�ܢ@��[9!Q(H6T�W���q������@ƪ�J*����~���U�:o*#��@� yQ�1$��0�� ٨��a����8����d�2�'����t\��u$�$5vP'�O���ߵ8������#*�Oq�?�Z��R����dq��$����?���x�I�+p����q�_������r�o�^9?�� �q��GW���S��%-'�W��ړ��%}ޜ�w"�a��+�3����"ڲ0�$t�����=�H� =��iP�I�jo佥�3S
Ul��y���2�{P1����Z|aLE>��_�y�Q������f�!s�u�29Xf�S����®gi�,��� $3������S�b�Y��>��h�|�p*�G�(�"�"�u�!��9+�)����������Br����.�=�`��zZ
Jsx U_�����iހ�Ƨ��u_���V�:yM�W�K�+��R4^������b�+;���f�����F��s��e��-er��tt�Ө��9?���j)t��� ��)�3��瑥�r�ן�~���S5����DE1�ݻ~��0���V������w(t'=�@ɟv}�r3z�V#���Yb��l���;�C^�2��&,��}��&L!�0	��L���Q
����u� �D��c�ȃ� Ct�T?�F62sۦ���
2�\�����G��*���c�P�{�}ξ��h���͢0+՞��m>3̨?]�5v�U�͋��h��?���W?��?c�'���-��zk�=���߃�'�'�#��k�=[����<Lxjn���X��S�Q������켾o� <�h�"$	#m�߉����!08�B����@Y
��U(F��M��5��*~@�Z�q�������*�����3aG紆zQ����G�%U�庣�<��S�%�������(�����TCC����Y}G]�@�Ȗ���לw�����aN&�������lN5�c�N9m�ci��c�$J|���:yu�Fҿ'�=����	Â�R�
�G�?�l��ii��W���&�M�u�OD^�$��\LƨZUVs��"�L���6}�G���J72�$��Q7���c�S���س��]u�n�#Kp��)��C7U�����6���^G�iכn$�71�2��̽�jS������{A���ER�<� �=�{q��ԪB.%_��gݻP���e5׮i��M�L�g��Es��<��Ӡ�A�E���˕
l��UtW
�����Φ���gQ��y�5�?��X�Рȣ����n��Ζ�f�OrYA���+�ﶍQ�k��K���d�T� ��I�uq�&�wU ��9�b�3�z}�7��V��v��O����aI�Ȩ=�^�tC�\�+�u��!9I����"&�xߐNnU��}*e<�#!��}�y��Q�~���V+�!n)U�Z� ��xf�Gy�C0~#e*�[��r�z�"$���vP����Ԟ�a(���W^7[Z9yl�:�;k�o��W�.
΢�t���Z��ᖃ[$���`�.��t�1C�-�?&dյ�>3��d&��3~-w׊�w
z�sC�)���9s�7�ܸh+�Z;�~�0+UT����p,��{B�|[����΄X�ƓJ��h��]'q^�j�
��'s-u��`���{�h'��BA�uSI�!�Osm��lR�����G�>�H,��b�Ʋ>;N�}+�u;Kmp�ï~7�m��z�}��
.\�I���h8�P�ux���W����き�r����u*	����i��-1����ӱ�c��MNxʍ����9\�1��y���{~wF��g�ɝ�s';\�v5E�2Z�%�^�&M� �	n�f�Z��\�6�6��Si
tY�OU�/(���l`??jL���4����rA<TM�f2K�����)�?b���k��d�u�j�\{�n�C��w��	F�}���)�W{Z��ЉȮ�r�l�ķ�ƉI��w�ہ�ŹO�HG�ViR�{G}�����r��s�H|HC3�<XF��:vL8U�r���M���㸐l����)���FX����ۻ*���k?��������k�ܔg8�;�?=+���:��� ��ߦ�ה����{ݨI�sfp×���Nޙ�NT���L�7�T{z���
8w�jWvm�Z��
��]y�����W�G���<k��E�|Ti���2!��g-Z���mwe^zj�t�oF�"�=���w�o��Y���?���\��]Y
`y�j�q���Yf�T�����QY�6�<O��^h珻{x��5I��[����;�c���O�S���#�"�R����E��"M#$.����wğ*�AN|��yA�B��o�:�R���l�h�w�1����B�RF���5A\:�"�D��M%���x]}{�a~���k���b��s��sz�Ǻ��Gf�E���+7eM��'ލu���[��bm�'�*�$W�a7�>���<K[bҦg8�N�N��x��=�[r��W[�.�6�ݖ��U&��1�uב-��{�bAIS�j9�����S�a�������;��"��Q ��{{	��9�J��?H��d�k{%��`	;�W��-�4�:x�O���5z[D���5KY<Kiq����4�m�U{�����1���g}�%��e�s�I�	՞���Ŏ�B����0�B�v��oκL��h^�j��==:��jq
?pTϖ���Bn�$�s�tȻu�kߐ��݌��g!�$]��O�Z������i;� Uz�����Opn����I{��2Sw���ٱ�Z�A��
˝�A�f!�z��7���5�fb?�Ň��_��d&��T)X��$�ժ$c*����_/�X6��a���$��y��#��iuW���6�M�׷��c�M���7HE��Q��b�Ɖ�r�,���:c���g7�_ιؤ���,n[�}w�$4\�K�]�I��*�)�+��-b�ު�٥����~}�M��Oj4���o��f��Ua`*�c�ccs=�RoO	�<��\6��טY����,x�{L֐�n�/8�9��{9�H�Q�6��}�����3��[��cg�$���w��&˒��������1Vo g��g�El����)u鑅3�9�����;���A��'_���G}8� F�d���Խ6���}(D��w���ڞfk�~6��Vk�)�h�.��$T����g�`^莦Q�5�W�4Zm�;;�'<�FV��� ��z)����ub��)3�#�r�׌h�9�#$�����Y�sk�g����u`�#������Yʥ7�[x~;<�rn?G8��f�gP(�|p�\t�Nv�����s�B�/Ȃ�����ڼ�I�C�R�өk�䪏�zk�O�¸��fN��휺]T���`k�q��?�g�� �g�fo����+�`�w��94�yz�W�3�^2�1����4_�$��fz|9���"/4���Y�G��դ�Ӟ�3�N�U����N�f�C0>Y��N���F��/eb�A��3"��
���ww�2���*�Ҝh�L���z�C].��q�@��"]��>u�����v9�O?�-�gFӆ��ںo>$�^l϶������;��y���4���&�>�<ds��	��4��hԬ�41޻����T�zI�\NUs��&~��O�'�e��W����hc��w���t �Ԙ����p��׼�?�eSJ���z�|�℞�ӴJ,�>���	#�%����	��~��E���9��]�֢���E��/G)5(�t�=�,�d�s�#7f7�U�P�b�|�WG���~l��v'��d#E�q1�w�&�JXf~N�az-��X�\3�`�u� ��i@ނ�b�x9%�jK�c ����T��e�J��JfS %�5ť���2�_>�F��Z	�)p��h�ɓoy7��zOEok^��NØ�����/�G���*��w!�
Dt1���R�Ȧ�W�����8~_�%o�Տ�����!�{��xd 5�$Z���s�eS�*����r���>���l��L0KEP�u��d��x�ak���?���mNL�K��$��_����&��m1���q%�%����n���k�ّ���?�Cz��H�vаV��ӎ1�s�v�B���J��Q�j@*��=\�|�l�'w��:�����P�ksC�c��CT����q^���՟{�G������l>��qy�d+��؉�u�o+L2�;�c��S�ڎ���g�
��) z��U��j��-�W�Uؤ��@�	��o��:X�>Pf�=i��5�	y�p!2X��r����olS0��ϳ^2߁�C���{�U���Rw�8�2q��c�������� �I��j��ڹ� ��v=}����ߘ����/�~���YH�'~8���ʾ�P!�[j1��Q���Lw��dA����ȱ�K�g徸c:l���|�h�K�]��c�8fi��-6n����bmuIE���,�.?�6�5"��ܡZ�>�ީiv2�S-�F[Z\S7� Y�n|5U�&`�C�[�|��"+��tN���&��`($�6��ۃW[��m�p.����y$����<�&X����L�Q��w�£��c�|×�K?<��~�1�|1��P�*��q^���IH�G�껞��2��\?U�쵾�}�U<T_�R�-�	ήD�ߑ�3X}�o�̊%U�|_9�.��zrP��>.���;������b��aC/R�F�H'�Fu:z}d���*u�<��}\�~4RftuN��[���b�X��hD=�՚
�y^\G^���x�A���R�B�߄���n�t���q����?����*�Ķ�����j��!�ص�ځ��������ʹ��n|�cE�G�]�ͨ+�FI���w)��Q���Ϲ��:�?��c��ǀ����C����lj�ꍱEc��b�Q?t&����m� ���KBd��ۛ��Rܹ�<i�e�x�$L
�^$n�Hk�x*�wۀ�^���Pk��{LJ�SVU�L�������z� %.~�^��~��MC���4=u�n'+�ov��-և$��~\�� ������T���
�����-]���)�벞Pf*�;g=`�=�b��M�K�"aR*��>5�y�ס�&�0��|e�>�#���7��@����w"���em7��������]�5����(X8�FB`3V�$��,�^�����i�Z�H�B��1�<d�|݇��!(�g��$Y����u�=p��j<�]�c5��(����Y�����"b� ��~���w0���㖛���$=j��=�U82��+:/�����ؒ=���~pb�p�[�`��+4ģ�<�ޥt����.~yG`�u�^�r�;���;�|�A�PV�1��Z4��v��F~��jH��cy܎b�P��������)'Z��>~�����p�,��dY~�C�O�}��e�[�)����<ʼGn��P!��*Ho�EEZ���O(�|�%�5�`�m�j^A*k��n��KSʠ��]����q@�c5|�Q�������`r���Y/����B|��k�A���ꍝI
�JR������-��u���Ϫ�x�l<n��]���7I޶��<u�_'%)C���_ a�)���+wA.m����	}�*������ǖ���|�B;���y�<�'E-��JeZH}��q�~ �Rl,嗂g5xʘ���}e��̀wN���ZH�(CB<��|���4B������b�"��;z|ُ����Y���I�>���O�3?�����/2���8��k+��3aX.��i�m��}�'�Ru�W�Ĝ��0?�חD)ؾ�LS=�`�~���]r�3l�����F��O�J�+N$I������!f=����`.�([���D��{�I��BH�w��;n����l�J�b;�7&�U
|�k�����MQ@ս��O��-��X��Fu����̞��2E�@��O@��YݻVڅ��6�_���+����7�O��Û��/�%���?ؘǮ����r��c�v'�c�_�c��&��Y`����R��J2ս�T.a�0��F�/Om\�������<�	T{���f�<�$F�s��gDV���n�y�����$	��|>Bm_���ϨE����#�󾧗�,�l�_{#o�%���^yi� �y���r�����C�'&`�؄j*��+�����D!񹟇�oY�,AO[��Q�wOM����WN��61|Ym?�|R�Q}FٝE����6ʺn5F�T�_�gq��	)벰�Q��w�!V|�kA�E�Z�Y�M�B�ǟ�|��� sBzY�}�le?��C�W�iP���'��-��_줤��9�m����`¡��!��b�O::IO5��j<�9�e/v��0u\Op�Fq&�z����ejdj#�bu&�����DQ,AO4��cu�,���l\�{unY�&����Iv���3+��0��x��D��!ea�/'RT��v�(��m����q���}HH���D�#�&����)���q��:aD�3p�p��j�:Z��?o��ag}���<�Ad5�1�g��'7;�ٮr�vaw̵��/#K	]��>~r�7���u!eR��o�+���F����Օ��*^��� PK   ��xX(	��I�  &�  /   images/f33b8d1d-9a3f-420c-bb18-27c74f47ec1c.png|�uP[�6�'8Žhq'8�R�����=@��ŋS�xq��bŝ ���M���~�����̙̜9g/����<k���"��M�  p�߼�  �P䵂���#����Â��w �^���Oe^ � �W/�<3�31Ԟ�]ݷ�=8��36�X�g���r6��de��O�ɡ'z�����ל���f1�.��
���E��q�\�ѡV����?�m�_���\��g6J"J �o��x�z(��+��	�p�����������訯at��:�����<3*�����0���B��U>~?9�%�# ]["2�c;�^���5��6��n�Ba�|��A���1(h�]�I����qaAbO4����^��7=Bcuv�&ۑY(�zL�$���\úҋފ����2/i�K,�>�����-���р;�����(m^�@@ c�?������8����`9F/W� g�~��se0���A�
���m��� (m�8)���||�o0]M1�_UZ�{dD�����p�;��cy�O��&2Ouc�k}�r��A�F~�s-p
B�� �oO���j߈F2�1�b���>q�i<A��N��ZC��7;�FE��⇕h����š�#� .�6����s���x=(�r{ǽ�-�P��
k��������>��k��e�ܔR�%F����+*
��0�Ȟ<W�琍��E,nsc�r'0]���^p��d��mvL-W��+'D5�W����3�"�H����O9�H�$:�qw2�-Sl��b�B[����E�LNO�����h�WÅ}Ӟ�vL��=:v|�k��������II$����_Hk�O�+�Gh{�_e�������i:>e��\�+4J��+��,�f�Gr,Xa�.���z;;u�/��4<:t�[���T�����n#5�aUN�ι0����B� WW��qqq�l��
T�󘬆�&:��X�꼁���9b���T6�Wts8}F�/v�A��X��У˃7�s��87w�.��L��Y! �`��f�PO,�/����L	�s�˦�Z3ӌ�w�=�F^�Z�yX�g<��ɱ���!�+9F1z�"�I�8���M�� \���
5��C��,��ÆÓ��w���<�_?����S���~S1
-�ΈH�Bw��R������7��,�s[Z��:�0K@i�bb��u�CG�1���(B8C�#���|��BE���:��X���ڔF����r��� ���'	�"���.W݋	գ����g�����$�'qs-��#%�p��^��h��C,��(���!�][�z���J�[3	��6���vʑ�\�)��=����w����8���'��m�C������B������D�8L�@B����!o�n��!E� �nq���4���7lzzz����%�����o�����Q�e.|5݃$�}�r;� j�&[k�}���Z�Lw|:��iV�����;��������+23A\Ibc���~�9����~��40�l~5K|/y��e��X�K5}}���ɤ���{���b�45���|)���+�T�N*�JTO��R`L�������o}0NC�:-"5��n�rDd�|O7�s��أW�����u��z����u?�Ʉ�׃�C�Fv��&	��|���{:q/tS�����]�E-�j_hA�[#�G����Z��T�}.9Ͻ]\�Z<=�H�W��K�aE}��W`�-g�Ӌ7�P��`�P��fI��?�6Wkf6�e~7�
�/s��LW�{��J��kX�)����K�x�ֲ��$W&99yr/�&(��lhh�9������&g�c�+5�_SQ�@�Ҏ�u�NVu���-oPEj]�tL�=]^�T�Qu:lg�/�`~{շq Q1�B+��@�,�GFb.n
�Ӌg�JI��CW�AP���
T�ꥊ lI%�"��9���q���2Md�Q9�Ln��h�N��)_M s�U�q��z�z��җ�f;	)zU��I�<��>����ˮ�PPTH<�9�6�S�Q�a1٬R�����E�4
�1���y����~A����[� ��$b����|q�3QTBP�p-�g�	[�_ff�9:��^X���P�{c�`�$� S�˗��GA��=���&��y��csTc��2I��Vz��xUs�wg�(�h�ԗ�3r�K,�ON�o|���ߎyE�� �-�[��/�6qU���Ui���zag�/��x�u��:�)���7���O�4��H�� ��_o���*�f�gJ�	��'�v��ZOd�_pPP���З<!�����)���RŢ�bΘ�~��L��J�7������~�����9`�~�4�c��sx;��eǘ!��d	t�xC(v}����e7���7&$O�����{����H,���BA@E�\�e_LA�����m����P�'�v��Q����w��VL�`�A�U����=�t�H�Q��5t���MV�� h)�#��An�Q��h��YB��7kIh��V����[+��ދ�-���Je��~�T��TR5
��ձ�mYRb�����%?�y'����,LC%�(��F��ы!��m����C�+
�(<�w/�4^!���5�O�yI�����u.�v�yG�Ԣ�/K�]����/�4S��٨4���v�^��V�C�w��###���?��m�FJ��5��w�'f<j. Ӎw培��WU�*��8)h^]�L�StC d��7e���7%^�E^	�v[V�[x���;�+,�������l{å����s �%8:75=�͍���L�i�ozϏ~lbɯ�/� Dni��\��I�C�hġ4��L'�A�эZ��@�b�J%���/.�b콺}FJ�50H���5�1����-+�^oE�t	?��T��Ce@f��0��?M�֤z�,gGm�[�i��Z?w��4��B�d�Wj	[�v�u��y����@N���d���js���J�j���	�[����6�rc���T[����$ಓc1�w�h:b����*:�w�dg��0�ԏ]�<�^{�_|�3g6��#^6<J���b7(�F��Y��&6ev�-<����7
�Mו���)�[7ېa�Ҧ@��o�,��_F����ռcx^R�6u�'0M�%$�5�搕 0�Ć��Ļ.6��f��o�\RH�BZ|�����`���=&t�(}~���K��K6d�b!��8�<Rxf'XхJ�|��9��h�v��W���t5����T����}�����}	(��Ii��wR��(p�/�V����"{3���M��+;2D*p��TT;ו�M^ޠU�F�Cf�Zr3߈�Ӳ*&��}�_�+G(ۧ�0�߂�Hc\ r4(���uG㗝L(N�w>���F�D:��؋��ӛ�z�IN���̜�/]�W�&�'�!�~�� �W�o���c]�;8�Db	o?H�Tp}��'��8��{���"OI!4����_���'����Mg9��-�ѝ����Av�sxhwV�1�5'�5^���v�R�����\�ZW�J��_xdw���H������s.CaaT�C"�+��9H���p�����dT�p�J����q�X;��5��'��c�����mw�h�C�jKK��1�����ld���~��x~~��b��w;Tķ����V�Ë��[.�!%k�q�B��~�Qm�~�#gD��ѽ�`�`>,-�΢��r�@�6�����{�v����'��7��o)��GDt~�����ݬ/�&.!A&)ݸœ��|���g��W�w�)ł~g���P-�C"�h�_�P,��S`E)Ӕ������}L�����)z�ž�H��(����|*X�
��}О���N�w���FgҚq4����ɷ�P;Ko//uR�f�*A�P��W�5֣�J�J�3aϟH��t���,�c��b@'W�{�\��ٝ��IO���[�٪ђb:�����Z����A&���ք��N?�m��7y ��'=R�g|�*z:��e�d���B���Jt�\�5���|��V�$�^���p�n��p>[\;w���b�`�C�2&����s V�������!�%3okJ
�RF�M�����lU�~��. �Ϣq#u^��rONj��_�U?j\F�:9����+�6�.��Q�2�ѓU�����g�ѲZ�t,�|�{CfK(F�Q�Sе~�����,?�-�(�'|ΗT,`7;+m�̦��O����j��8)**�s�k�5C'��z���A�,�ZXZ6��
ܬ��9>�>ggϏ��z�@�0���1+�`�ZW|s���\���[5�8�XjqDhT�4� ϑ
b�W9��H�F�F���i�8
 ��VWӄ6tϛ�� e�b�� �-�T�ʦ��Ю��*T�pn�rqN��.R�)|O�B�0pg���CX`,}�m�������b���'�9�C�#��M z��_�N]��>�8���AK�b6o�	��KY4:,�\��҅����e7H�1h�xm�'��/�$�^ �ߜ^�w)۹��8`y�0��A�-g"\��7�P����r��OZ��b�P�b��̂
$�I���b
���9�d(y���QQ�������A��,��B"�C�q����fig�&�J�1b&bĻ�S���m.�{��Y�?�sZH+��}�����VPP@R�՗�(��	
 ��譴�{�]�o�Ч�(�W�;�cѯiO�j͂Q!�5���������;j&&�~�?U
KY}V$�����m��-�k<h�v�Y�5b��tP�����L\v�s�7� ����N���_�NNN�@O�1�T^s �	7h�뛫���/���뷰�]:ɔ �u�RK�'T@>=�S�6,R3�D��K+r��h9&5�1<���FFeB��[�1͝��-���g��i� ��f̡s&С�<��.�%K ����pm�#ݷ�7cYu�}�R��c;
���;��t|�~hw`��?	��LH��{#�S|#BpK+���䠟���}�Ԁ�G�&��<�ha��'1mz������c��PSa���=Ay�Q��=�<���N�R���i1�XR�شݠ��ӋTK�G�h�f��D'5�����vҏT���[I�\�gfcD\���e��*�8_�٬�G��ue�cr��:��C�t�*�Ă7��^��< �z��߿�UUU}=%��c��mk0b��vL��/��#�W[��S7��&�3/��T�&G�
�c��m��:R��Cb�M���2<_5��c mݹ��tQm4~|UP�̮�C1ք�lSh�6�Z�1�Z�6�瘻x0I��A�5��������s���T�m_D%�]z��?f��h�U#�꒒�����F�n�:)�i��� �Y�	�d��q��9-C�V�5Ԃ�����..tZ	4r�����c�#���'��!W�� �
C���2��2��<�50�"N�羹LUR�t��N1C�+Or��>��+��@�O�nF�/N9��ȩC�h`ˑ���ʎ��9��糎W��� !<X^[�6�С8��M�[�q.[j��	���7�!�
'�6��C�Ǳ�֩ۼh��q݊X����D���Dz�����#�(=�0*|�z�u|�VUj�о㥧u�%������SP`�{�D�B2��01qW3 ��5SV:Z��W��yы]��r���50[��A�A����ُFL�Iv��s���r���t$�A�2@���53C)A���lI
l<R�������ִ�;!J�ݲm�B��fe{�q'�`~���Y���︬����T���0�?!�o�8���������b�|�wq�Ɋ���~����c�;�'�o���dO�"(�pӎP�>�_���g�+�̈́���g��ZIm}?sDU�|�Hk5�brk���S/���<W��;������.%��ET1��l>E�I�v��DA��3���1y��x����T@��^�mt^z���0:�Vb��h��(�;P��]b��Vy��,�)伷�I�1�6y��IR�c�m`�� nSq��Ħ"ә�Z�;����"�&�9���7#X!�*�i���FOJ2(+�a��kp���Ȝl���)�H2d����$y3��xR���F�N��h�������k���p��̓�2?H�/�f��=�WS�̖A^�/~�6Z�6�Y�]W ��m��K��	F5�����Z��b�����X�Dm��'��Z=�;?>2Lp�ay͒Z �uɤ�m���f����i��Sȣ��Q� v��vf#�%{tI�����YQڰ���D(B��������o�^�Gw�Sh)���	��ި�O���Z�M����k�N�����@�`��;�cB05��SO�=�6��5�*5Y���(���8'ъ��@���l3����KL�E\��W��<�'Mdr��*x`d��@;b�NS||S~����U֦��x�m��u�%a������қC��R�-Q;�͡�pqJ2��L����Emj���sy���D���l�����zK�6�Z�]c�����Zy�ئv��i�,e��Q����ɠ�!�q�α_R:����^��v��{���W�ul���^~~I��&ϓ���>0\KAA2S� eu\{NIt����&L�����5,X�)_^N�����;�.����������5c�ލ]s�"��ȋ���-V꿚H�u?��j�?=p�����Ǝ�v�~���
ә�sdC �����w��\��=��`ѱ^��yG�]$MN ��7[P�v��_�n�NƂ.ā(S�<�Yn��@쉊v��MV��1>A�s
���8PvzY��W��b��t�^|2���|.�I�
e�]A�!�t��^�Q�N��]C���6�*h�6\k�z[;K��sPE��C������@1�?�ڨ��ī�x�.�HMl/k�����kQjĶ��H'e�I�@����q������]�;�X �ݒV��x��Oq?|�#��U��!�%�0�
i�����}�����Xx�����P��LX��S�\��cL�GEX#��w:��������t�_�������~���R��aZ�|�w RW��j�3�#��S�3zU�94_�k�ӛ�d����?⼢䑨�Ju��P��8O�l$�.G1�Ky=\R����t�
��dB�RA(���"4�Q�J��1�Kl]A������+��֯ʰۂ���y�Obb�9V8����K�V�_�S�.Z�r�w8�"
�VH���+r�n����9Qn/	sN�[�H�����Դ!-����5=���AL2!�� �t~J����ͨo��2n:���^lTd��9����j�N�Ę���.N��6ć�����x�Fl����H0}m�l)d˭B-2����j>i����八�0�{ukԾ 0�+���{����Ov��r2�.d��A}]�n�"s�n5%�l4�ǚV�+�6F@}�=�
Ȯ����=����R�g"b�5<2π�_����� ]5L�ژ�HȈ_�E|[˂	V#?� �]���|�f	m��Сu7�!���h�[)Z/OL�rn�� �4
�f�;���)���zg�C�ww� ���@P�<���t����,��eK�1���~)����5H��tMI��a������8g�=$ @&:o�o�6���1�/�`T�,�B��0�l��[x�
j�yz,���)2�5s߰����4g�:`#H�}7��Xf�?#��oRv���'�]���U`" ;�G�hic�O%�_�wq�M��]���T ��LI�,���c�%Z��jw�+�sDLU4������)���ɨ� g��s��[�*�s	�J��P�R3:�4��.n���fro�vB��~���w�����ov�6D�O�8ꀜ;��(���n����`�΀Uk#`��Ϝ��oAAA��>'k=�����F���+([+�s��lV�E֑�I9�#��]u��E	��z4^L��4
��xe�p�-��Ӓ�ɶq���}=��1�]��AO�^��ˤ��N�?��9��oqU���C��mGӳ��F�oҠ��~�v�m��~u0�"���6�e�kk��g��0���Y��������4��o�����W�3�����a:���c��+����"0�� �<���PGr-%	�b#!'�L ���jTf/�{+e\=�eM�xc� ��(DF7�8c����<���j���+T�F��T�H9��3"}���4����;�b�VZ��^bX��Ķ��e^��<������/	�Gt��w.�ܔ(p�=�b�Vo���uY##�;%�)0��7s��zH�{�e��G��o?8箭?5�(c@E��A��<a4�8K)�H��*8+��|�(6���A��O%�Tz���`��88J��� ���ٽ��f�;�aட��-f�W#��/K,���ۗ�Tн�Il4TUt�[�fA���������]k;�J.��|��҆�O:Wc��3�V<��YdG�P9c!��S��y��~)��_o�s��X"m��DX�����y?6�\a���9Xl����V����#�������/2����͖qt�D;�씶��Hwj��u,�wC.�5�a��)�#�G��Qz�G�kx^z��� �x�7�F�Vo��k�S���2D$�l&�)�|-,���<$O.VZS���[Ldd�E&�%z�yle��N�VY[pp����l�vn����'@���U �E+�g�g�	=����~�����2���uʜ�|�����p���[I�ӏ�P����Z��������������+���BB)XP���[�LӼ	bY����>AǠ�q���ٶ�tC���gtH;�4I�ם�
�x�$h)��ﾇu��bگv�v;|� -ظ|��.�h�@|.�Q10��bn�Z�Z��?�c)��������K�:&���|>�ʂ��Z��V	�Kȏp~�MD���8�`��4�ɰ�5�(��(�4J�����;Pm�`ab�8���� *ޔ?�b`S��_�2_�PC�Z�|d��L��\��n���1f67�D)�Z
�d��)�&���1,�j���~�{)��ݕ�n��m�69�I`JpʽF9ȷ��j2���]r���������~5�3�y��օ�w�C�T�������������߭�Z<O@�14���ŎK���G˭�� ӷª� 2v&��̽��\n	�����!��΂���F��ohWm���WDf2-�5���J9����,�U��z1�B�:����B�H����b���U�/�g�xq��S��-���9ү�,��_l��V�@�w�
����|�������ih��U���4T�ȁ��r�k�� j��!�G�R@6_]brbU3m�=`�&�i<>2����?��}%/<���zg0%]P�l~VC��W�ygT�iX�X���d4
�����w�)�����6%�����{ǯ�EEk�"�#�2%�� m<渥�����0�ס�7fv�d�#t/o٭di�@���j��x[BЛ�HX�>{���ܜ~\V�JB�O����4��cφ���;�o�@ϲ����q�d�'�];O�O�@��x�1.��I� ��˚O;���e'wW����%:xB��n���Zmoq��(zF��Y��S��1�݃h�Y���ۏv(-,�2���]�E�)�-�ٻ�������;n������K"����hv��2���O�xE�J_0�[�����R�� ��ҵD� jYJT��ZԨ;���=Ũr��J-���`Ѽ�.m�ω��F�jl^�k�߽ڻ�gA?a�o!�VB�ǌ��!�H��ĝ���RR�V���X�!�	>K�["�1ʋ�����Lʌ�)�v���c&PA�3�?m$8]��Ƌ��	�G����O���0���߼����T��~��P4�?����� L�����;?X��
\���,��1���2���r�l��_�,��2aFFγ���8�y#!1���R@��|��84�?�G1����2$O����1�oyW�c��Y*�q�����\ �Q�ְC��F���?#-����#.�ia�K�31VC�(MPi�
����d~�;��>�
j�f� ��VW�!�>����iVJ���EL����{� s�������ׄ����f]�tu�wɼ���2��C�L�%_��������{:���~X�l��

��8<#|#<�O`D�z����9n�� F��yN����`}������' B!�'�5�Z���x����-����+�𓮷YK߇��T��8\j�.�R�m�G���Q�fI�h��7�ڶָ�Ju�.��wr�q�E��>�f���P�;n�R'b�t��q�T1�n�M�S���D��x���W|s��(�ȅi���!�n�5쒨ק��T�XW!��٫�_Sb>��ד}6<�q��џc�ꃘ�t�y��
�,p�4�t�,{��X����A��-H�8e>X���?���%fߢ��F���3��y��7�WPFj���/��CR��� �����MF.۾�F�)��p����F����0��c^=K�����0��1�Y9��ǉ�sq�����]�׌�V(���|���?��cV�
]��}[�A��³�����5�9/}
+�O���J�0�
T�%��%����<΅��'�n�U��'��Y;Ѝi��vv	%���qZZ��*'��m6�6��»���&��&�^��OD=���^�=t�ѽ���ꋡ���.թn�:ϕ 8lG�׬/�C������N�liS�WM/��4�[-�ڲ2������=�$�'gozz'}��f����X���<w)/�$H�(�q1���맘)��X!�$�I����sh��g�b
'�*)��ɯ$b+nŎ�Do�z#]A�^Me,��Pf٩��sP����O�^�$�-P��,�b��p%EVZ�%3������%��]|�P��9�)\���"���g�sUz'��Ǜ�TD��#�X��,i�=����$' `��4��~_���;����'���o�)�p��=�Ju�Gכꦽ�L���QJ�t��Ϻ�W�T[$}�h��:\bG���fg�/Fy?��c�q��Լ"�bl�`���="�����ݟ/�E�Վ���>����=!��ާ8m�U��X��Qc����]���b�G�]�6la�|���9l�@h�
�N=�T8�Ά��Xs`n4s4�����Y��<�s�!��by ��
/}l�8s�t���������ꟼ��s���hW�ĲUs5,F��4���x 
N.S��g�߭ ��/��Ѭr���%F�َR9h���
�4�1��^&�h�rvz����
z3tio7���s�}��o��L�n�b^R�A�ύ��}Ej��}��d�_�^?b�����i���.[#j�ڲK5CCJǗ�d/�Č\%]\\^@�HI5���q�q��-�_8΅t�R�(3@h�f)v%�At��j�;�ff�I�}�,�K'Ng�sTW$�����&z����us��~t������O�Vp�[j�tH<��󱛛��_yr�%%��}==��MM_@�m;E��vvl�������t��	hk�_!w�-��l��'�QL)�	"L�R�Z���MܫTP�7�I�R��&@�hȲ�/s�(0��B�����n����������	200((R��������𰼩���O'��<<r�Ԇ�B��d�^}(o~XÙ�s$�tE�C'V���2с�6�#i��LC�	��T��
�� )��R]M'***��5@f|���4ʍ;�Y�r{y$��V'MwU���$]��#h���P��V,pyn(د�w	2�?Hߢ��q	�8��K!���M��Y�S�]ᘬ�dy��n28�ʲ��`2Nx�g��`����{�S��w�PQQ�>1!	�7�y�=	��'����#�q�_��L�L�@,���g�y��ns�~y�{�"/D�Ɖu9sĶ�(��G�1H�٤��V,g|�rŰ�>Wj��N����|N"����qEy�d�ve�w���8ǣr�P���|�[�$:��%�.2�:^��Ja�+Ǩ���OhiG���E��*(�22(��W�/}:��&� s�k=`rQwvrn���< ҹ<ۅ�ıeK���3��<�@��-�D�OP�����C�wu>��G���V�-V_�����j�}�N��33� :!Gj�#�?�/[���/{{{�y^.E�"F�EH)�ϻ/�^�1�4z֯��y�)8���"�h]<����DoR'N�Αp����Y�J���{yb�$��XRR���#y��8m�jh�JW����OD.��.L&�t�Ugr�i�#ț����:�r�_�v�lӏ�=��4�]��Y�?��vZ6�f���.�<� �ll?Á&�g��o�vC�}�����eQa�eoϧ���`�����غ��@@��y�^Ӯ \����V�F��9S�Ϟ~�'0���wH�p�	܅W��;522�D�
u������e���u�V\z��'8)���Թ=&��:5%/����/n𣥦!�%XT��x��*�ۙ��ƧME�x��$�"�;5����ki>o��:��������*�fڟU/�����t�����bnַ���e�8!A4�+�DX�
11K� bWr����&sf��$���#���H�~����YK[������O���VR�4O_����h#9��@z�#��B�]Pȡo�9�%��1ڵEq��o�^_H��DQـ�镌������y�(|�Ή�$n�4=��G���}![W�yG44K��'�H�0"ɔ��anv��h����*�I2������ܒW��� ��1+�b|��ݷ��o$���)�[O��%T�C��R��p����Po��B�����_=�T�#ݕ�x����]�T�M�����r�s���������H����V�c]_k0_�(��6��*���Ś2�o ���!^'��$���u%�ώ%�Yv6�h��������r��ݴ~�n �m��̫��*
WW��	6����9��N��C�O%�s-a�K�z�@�4�����W�=JB
L`��Rs�Q"����A�_�8�>c2Ȳ�4�"�����0��o���`:;��M��p;����[��LXJx]i��q^!GL)�Z�g/b؊����;'A[���F�La�bH���4�<�jY]���I'�V���߉o9���d�(�Ty;OeI���g����8k�l���̿�~��?�� ����b����_S����\��b�6؈gGfX )��r�gB^G_m��S'�2}�K �4����}�[�����'l� <�D͑B{D�?&Əe�'�V5�%��-A���:��ʅ��K���(D��Df�J���2ٞ-�D�5o F�������9?/�ٓ5��#�P� �!r9�-���ڣ��1X�I"T�I���[�2[b����0�l��U��Ɩn6N����S��F�U
�/p��?_@k�QMZ�kS,V��5k�đ����c���;U`���,(����T���Si�}����p=�o��!��Ox�u~����]y?�R���/�>D�UN�"v��Cb22���>%��z�(]`��Hg9��4$z����d���yiZ���v輆3�s�#�䜄����gXM&rkA�,0x��_��cR�9����Y��u�@��<�)��>���EB��c8n#Xde��� �4H���1���̐�eDe��K��8_�c��nҚ0��ʕҰю����W�;=��kX�с)�Ұ��`��,Sx�:�ƞ�'=�o:��o
����h�G��>��z�">_��^P���>B��_��N��'���?���o��Rt��o��j�Lë�L4�憒�Rry/ﭓY�%��\��u�.]����%�V_/\���ཤ��]_4�qMi
X)����B���
�W^�7]�,'���3o�I���Eݪ�l�CBp�ա�M��e�݌����Qz��=w��d���b@u�La�55!�o��FK������ip5\9J�� R��?�q�s�X���{"�F�h�Տ�~���i�Ǆc�}� 㪨����^U�"�O�	��|��yU5��4t��ce��M>�!l�R�� ҲM_@��kB|�ic)�lH	�M1�|�#��:q}���v��p�H�s�e��ߺT���BÍ���Œ@�%��Mai��p�J,��m�ِ3�W��ۓ�-��G�{�(fp��ͱ�M��cؐ_��`}q��.e�>�\��q�����q��.�ީ�) ��K�t����ˊ�oeH��Z�S���H�S�t�6d�Y��k���{1���&�_3�_���+~4��l9��o{,�s�-��a��+��W���yix��!/{���`��{8��yr��~����8,oED!��S/�v^n�8C���sz���%�_�Ѫ#�$6�l)����	��Z��,#�'�9�
�D��qσ�Q�^�7z���Ȝ�R|EE�T)���X=<P<��ӑ���]���rG�Cc�+s�!��¹�����(d
�)@�������R��Uj��RL��>�=M'\Nfs( 	��R/f�G���#�Z�e� �����g[2��H�����Lb�W�]9���o$5��3��qo,�zh4��8/�
��v���V�� �t&�Ư2�Ծ�wa 0Cʨ�x�^(C355�_�<��+���e_4�W��թ5k�����^����[�P�e5V��6Z=Q��\w�G��bd�ߔL�m��S�D���H�������}��)ޡ������W�R����R�N���I���(;Q��{������R�q3:�ۃ��+����yUɥ|� ��+\�g�������4Z'��o'`���uK���z��j�TU�5j�AТq1��f�L���EA��\�W�
|SA_t�I 8�BQ�$)�O���t(*��3��u��ᷥ����
˘�����s�[9q��iq_��>.���w�i�ݿ�FN5�,N;C�5��F$�ewe.=v����k��o��ܛO����Z�n2|z�q$\"�#�ʑ��5+�Eo��%7%{��t�i�q�a;�v����R����:�tI*>Ml���<��q�MݖF lt�Yȳ��h�����v���	K�%n���������K/6���Zh�������>�-i�E휟�5�NO�t��%�3�O������vt�tԏ��Uf��/2`uX��԰�0.xp��͖��2�Y��R7��t���Ł�Z�S����xM���L'vG��P��ox���#Q�N��,��ߍ|���)�t<�RX�A�Y���M���7��MZ|r�+����!����.?=@��Pf�UK�v�|Cb�!y����h���j�ꤏ.W��$�6��"�cï�T0�۳0|�����kȘ\�2�	T��(J��i�v����w�`���t�����<V���w	t��'�߬�vj��=v� ����>G����7�yh� ʸ��Sū�G���M�T_b�'F9h����Ȥd;-��V�!C�y�k�`�iew夛�2��`ʎD�����O���Կ�ZhP�Q�;XP�]�6��1�  ����8�h4-gմɍpl)趾��?��yC���7�h"�Qeۍ®������*"G��S��X�8�J	<2^Ù�G�8�s�S�]:廧xq�]���P�!��g����,U�5	��l��q �iU�l��z?�[��<���^�ql��3�Y��n�"�1�*�<�:t��
��eG���)����I:�5V]�%ù»4C3�]�+J�!�l�:IgD̙
kB]o��p-�ㆨ�C�ɟ��'��j�c3�q	�g�P�rEC5��h0�ق/���H}E>Dw^jaB�|�(�=4����G2+,=��S2IE��7b�2��y�sv�hu.
P�	��w}]�jh�K��2J�^W7�7|sC��>r���܆R$ ��év��#�&6�?@�(���p�iu���!�g��<s7����7�tɯI��N˛a�`'�+���"i�z��xXw�{[���OE��u�<g�kwOH�ώ(�:M���lV�Kr'[����[k��mdS!�c��L(�/V8o���q�9l�Vʥ֎H`@Y����ʺ˘&�I\ ���������(Cmp���Rv�o�7�r�Z�n7�i����4ު��)��\p�:��a�� X dU(Wd��`�IC\_�CS]�D5���P/
�0�е�S3���{�A�>$�뙕X~!_{���d���D��ȘjEc�%�ދ1R7��e'��k3���4����Qx�W�1���P�z�#s$��Kw\����4���!���g��+?����:�ܑ�7�[o���.{�3ȓ��7�� ��&�:��&h7�����)^�x�w)V,8�Ж�N��]�MKq�[���.������ߜ3;;���<�s�٥�xHVU�uj>�	��{z�C�UW��h���$���w�\�i�m�������:`5u���)���L��1�3�j���_��g*C���ݢ�l�V= �o���Jnj���`>OR�o�-)n	
j_��ޥ�r`���OS�]�Icd�e�+��Q��� � ��`�TJM�t�u,��Ȗs���YlOg���Da����(��#����r�M5�[v7,���M�_o�3�[�*��-���8���Z&Յ?x�vb�w�L0܆ ߼�B�����q�@nW��N�n�;d_�F+_l��/� ����D��ݲ��B�tZ�6s�I��7���I�H,��W=������0�Ҷ��D�=f����1-?��G�Ș����w�MJ��)u�� ��lH}:�/|�0Gr�4e��|k�U�I�Y�6��h�aC|�wB����� K�/]\� >��P�R���`M����4y}U�MC��6���Ns�<�տ7C�p��n/Gg�B2-�.������
��ُ(����#y�@�j�.�R�?'f��;i��&S����c^�l/��2Na�\���f���Z��u��CD�W��n��	G��Xe�߆U;b�1>oe�%7�&#�}&.���-i���]E@K#��PϤab�쥌�����pO�*��+0
�qX_��ܬ�9��,�i�l��a�M�gh���і�J��B�Ue���4_q���.N󅓈��;���c-��t �|B(����P??%姞����%:�p�����W��z��E*"$�x*��e8z���w3zZ5Lnk.f�h�t���H4��ݙ�kr�1W��Z���[��ȫ��i�����X�a���Uꀑ���N#x���|w�0w�ɹ��B{���M����ѐC�/�ʐ�� .�4 �����f!?Z\I��E������Y�lZ�A��U��J3�C1Ku)Z���kX�\(����;f{�Q�oM��(Z�P�-�6��b��F1I���M}�k�g�qvI^��(WPm��=)��jq�{C�uK��L6�/�cWEf�hq5~��hI�'=*�4A�2ǶsZ+#������QD���G������?�i�U���g^���8�֞�����"�= y><���Ξ@����{�;��];ЇY��i�Vu�#?�\�.����6�T*��L���+����1Q�W��m�v���4&�)�a���D8|��c?�t���?�El�d5�**H����A�|^���ğ'n���]�[��#�K&�Y��	��ٕ�6f���j�]*U�]���������b���u�_����$�k�a*c�F�\7��7_ֱ�����O>����T�����	�Έ�l�;�Ph=x�o8�����/�⏙������b�A��9uJE����$����eY��4��7�w/,M��BC����<;	 yjYF��[.�-�����0�*�����Oۇϛ ߾�4�|�ӛ��T��G��U��O���M��E�i���M�~@?f��4���N1�MQr S�v�ڬC�r����x0��Rq���gRO� ��ׄ����HP~T����=�����eH��I:bs] ���i^��V��T;��ϻ�*��}(5M%w�]�aX[�5�n�����S�k�n|�)NJ��%�bʀ����/�"���7�$z����đ�Rz��a	Ξ��.J�­J F������Y��]�-$=Ν�����:΋�ɷ�������6�b���O΂Yi�9��S��<����`"Y�^1��-�T7^�Q�/7?Z�}�C&���^Č�3|�����BQzѻ-!��'ا��G����l�$
�(6sH �
��[g6�s����ɡ��'笙��Z��M�%+/�5�(.��	� �Z4�����x�31�F8B\^�?���DDDj��?�	
~OL�{w}������&���E#�K`eeeqwu�wo7[?Ń��Cg��3b���N�o��u����9*�M����]��Cu�DX���XQ9�����;)�d4M*�d��JD�����$�\�r����3��:8`��̋�Beł$ �$y-f���L!��W�Gҁ7Х6��ҹ7�l��!�W�+����e�:�p)�����y	��|����2@peH&ǧ.�����U����Q��?W�?4��NUL���=�熭�r��W9>���[�֖b��;lu�\��f\5>�H<���_6���\��O.~�}]�'�'�����M�a��Y��tG����K<�%��M�v��o����bCE�Ϧ���	�����B��s�o}�"l,b���!HW��Б<:� �ǻS|�&RRRJJ������J�]��冤$���7��}GV�nq�̻��F�C��1�"�2ŷuϳ#Q@�}��H�rwN.�F�f�	d��%�i�c��A��] ��~�	&9�I��t�)g�Z9/��`���+��W�W�l��å��E�4^�����2/3��h�RG�K�j�\2��͞	��nY���xsFd�Ǥ�Ȣ���$���>�m4��������c������M:^�.,�]<�Uw�'��૫'~�R?�Lh�b;��Kf%q�S�����?Z�[��}-��|o��������fn�~R��������e���A0S��P��.׫�u�0�/y|���]�V��7�	e�CɏX�B�/�p"����&��^�ä��s)$��aQOg8y�X_��8�tfl}�+�V��'��?S@�
�-�1Y�:/ �Z���M�q3���yr��m	J�0L���D]Gٱ��?�l���WK��������~6�T�HD�6���8��"'�����^��*vR�En�6p?��e�������_a�A��3͝�]<�t�'�c��w�LNk�ݙdB���gm���:��;U��__����>s�<���r۽Ei�e}RfQ���X�ܧ�A��l�K'2dO�	�� �Mp}��d��w��X��*��j�\��nol���UXUX�¤T�epP��c��������<�����27ǋ�j��֊��n$X�L8WϹ���Ԭ�w�>
��7݀W���BU��f���&)ا����4Pq��������G����7Ç�1�@��6(��+���*#����p2�	G������R��ͩ(��"��I?�l��}8p��c��B�%[��ɕSΕ݌�F-�Fȉ�s�Ś�Y�Ǵr����"�S��l��R�k��K�5�D��ո���Mm0)�^��6E��߿
o�ؐ����Jy.����v�e�˨��8OOO�c�P}WG-�pP��J�}�Ù#;��Eჱ�!��sb8�ծ�-c��؜w�k��O�/P~Et�;k�j<A�w$�t�/&�V%�*�2Aw?�f� �)�K}ǣW`�W�0���0�p�ծ���1�"[�~�9JUU��ѝ����6��JcV�β���s�8����BgoB�����<�X^F�J�F�i �p�Pӎ�hb"�q�~�~ :[�n����Mz�ҟ��=p���蟢`��������>����7l(d=F�=3UWo���(H�~��o�;���l�7�j����^��8��vlFA����t)J���ꠘ\%�u*"'�*?:1���@���7{L�k��D8�(��|]yydTK��ꇗ7�Ǯg*߃i���n�쨼�X��
���zZ**1��7�c�y�?3d���F_m��w����8O����ز�4$(���f���)|�c�9�*�4�V%�ߐ��舆\���PhZM�tnnn-Sӷob��6�=���;;s9H��{������������1n�k�HsP���,�L��Wx]�Cz��!��t��Š�	���
�/)�hzx&�(�����/��YYY�#J_�+��?�!��÷/��P�nz�
Io{\��{p���R��Wh����-�C�4�7a�/N��f�m]�����M�<������~`Ց 
9�?�^,���� 
#��Z�g�M�F��=�Cb)�!{e����� ��H�K�1�a�����:y�t|Vir�'0$P"�!��	�E���!�DX[%�Qm��#]���l���o�\��	�Ì��p��80��M�<�l�,/OS�QT�~���grk�(R携$�'�7̠x�X�R�W��2��� w(�v��T��ݺY9��X�&�;^VJ����xʝ�Z�: �մ�!�U!j���>
@b�'�E�jp/�u#Z��v��<6�$��^T�Q�vG;��W���E�C�@ �K)��8��i��х�f6���3�����J#c��{�n���HA�ór���)9�U1X�h�G�}��F3[�,M�aIY2���[ng���r�nt�)�R\�g�P]S�b8�H���"��Y�'`,U��RG ���`�z�v�[m1����
��x*�6D�#-��[�X*^����_e
�����{�E2 H$N��=(B�^�z�~B㯧�'Nh>�ǲ�1���o�
Dr[�1�2���}�:?b�5{����1y�j���ВT!=����m�Nڹ�o9��NX�wr��C�ɟ5�K٭h�+X�5�e�=��G�.j,�~D�%2�m]��<Pu�N�@ʿ�?3�:�P TxNayZt[��<�פ�`.֪�q���y��Ɉ�Zu�<&�����Ub�0 ��;��ՙW�C=5���6~od~�*¿�-�����әB7{�r#�5|��}0��/�-��ѥW܄�t��;��=Q�f�\�K�f�����S�i.�D>��LM�T0Q�f!��5�)�d���;y�.�-`�jX�_Y��9�wN"��\m�ұ�\�����ʽuWѾ�p;u�]�L�i���	kz��+$5���B� 5b��u�Pa1�K/1"/D� �2�������çTo���vOxNa���R��D�e����z�ng^�T�����W1����M1�E��#EluD!��y["l��X��2��� �3S窼Y$����r)�E���yHC�������<�N��ޖ�XͽXDZ���(���/]�����4�|�ӹ���}������ �<���1Yx�P)Vg9��گ�-�V������"Ү�~f.掊�e�������?��� Af�p��pi�ᔒ|�ک���Syz��`��s��Yl�P�����ʶ�:����9�����a�H8d��gϗͥl�oG��� {�]�$%�vJ��l�FE��fl�]{�&�PM�k�1'm߸W�Rt�|�rw9e��Z�'�B���[���	���xRc� *2m�8���v��dRb��fpȣ�����f���ʙ�|TH?̑�Y|��@��I���+ݤI�}������f&��hkhbh��p�?p 6���yH�b��մ>Cї�,er��V���d���z�[����2�X)N������r��I�vBRI���^�K�lBhf����3���n���"��wܱm6�o)���f��P/�I���7�Zl�a�E\3 ��rs�&��T�%�/�X�S��:�'����onˋz<�i5�Y����PM��q(����\2���9��cϹ��{�����H�(�4zȻ��?M}��[�e���������ƴq�t��vu~/���CmR�w���s����M7����5�yo�g��Ŷ��1l���*y�$=�$���l�U�PY�Ey����W���rĔ�q��kj0/.'������:b~[�%V9�B�7���6G�-�r$�N�Z�z{�b�t��սj�,�j��6�{ ����q�l#�-i�G��3|�-L��c�Ꮢ�4� ����9�Cs���>�_�U|o��T�_�F�^q��Lz�h�Q3>_�\/�ɽ��WX�1�}U�	m���w�Am09ɬZ+H���ES �s�P�F��?��`:�#~o�߬%�~����6�>N�@�3Z��xWӈ�6�lՅ�5E��H�Ġ.�>�T%�-Y��3�9�R�������XN3 ����0j�E�/|u�8|bf9ī���x�p��]V:��c2_��9���w
bކ>g"�P�g�H�zX��������P�/]���WH. JZq0;l��5�ReH���&�&��ݗ��}O#c�ͺ�����E�4�����O�f��I��dU3��Q��Y�����5�?��`�_���yv�)Ł���oA$i��0w�����w@B��A�p.�;hj�s�vl�M:���]��wB���sL_��b8��~� �|b.�W�z �~�R�y��L4�2�W��fp�t�`!�J>�����h�[,����7�[�	�<EiG�6a%7�:FJ5���r�=s��_g�o�T{[x���'��Q���qȝB&�o�Ų���`��z/�8��;=ץ��L����i�0n��M�{k��Ա`�E��j>r�7�	�_`�ÚN�\��q�b<hm�����O�E=����v�N�B�d����ڐs�e�Q�[aʴE�DB���E����5��<�8jSy�k�b~ҵ`�Ԝ��$/�?V@X;��W�s
��}��� $�O�Ց���v�m����U�biz[-U���;�&�����:[tw��C��l�����'j��Ix�h�+�X�J�1�2уP[�fxmX��Gw��o�0B�ozn��D[/B�Cl�+G��j	�5�pl��^��������j���h��폗�����g؎7aY�D�,��7T���I�����S9�,�8�l�����E���o��9XN1.{�}�z�E�	�)r�,���ѫ�%3��S�R=�	��?�~�܎���B��L�\l҉��;��;'�sr�?x.N��,��>(��{��E�l-�%�)����^��O�Ǧ��d;�_�V�/��!�7�-��R�@}�]�{�}	��/�]yW�xH���N���{އ����(����������
�ɮ�8�j�����*fQ�y�������I�>��L�./1m�6�B��٧��I��,3mu�J�tޜ�鯫�nn�vqa�ǵ�i�a��1�kH�uWȊ�3nb��ȫ#Vo,u�oRan|�y��
��[#��D����$i�u iE��5&]t1��U�y4��<)42����~�//����W]���>u���H,����D.���$@�K��E��C�*�U��^��k�{��"��]��K�<^iњ3��_[��u %�l�<������������g���a�
e^�������x.���V�(p1�N�4Ê-uS��f���/�����}��-<>"�{]��.u�ܶ��̘����-����,dPN��0r0b�Dc�.��Z���!!�=�3�k����᫺@�F���鼰�׌d�e?:W����p�=�>U	ݮ��|UZ����S�r#�s�T4P�k�ltȸ���S����NWP�ݝ�"\���<�\	����T:�O3Q)Z���g 3��g���5� �F����0q#�����b�B�O�{=�嵐����M�z�F_���/�����I��^{Y��q�/�Z���������J~('���R���Sdp���׾J��q�~*O�0�Od�U�4۩G6^yi���5�c�*���
om�v��&��~iZ��Eߪ�q�$��_@����J�[7�����m�*��1��!㏦�=
L�X�kҡ���i�\��A!eˢ	��D�~ ������ �gH%�Yժ��,~~��Bs��08��<Ь�ڭ���2�"��Ǯ����[���mE��{kr�3U^K/�'�����]3�G�3❳T�͡��f�v=?�J��m���H4�z���)R�تq_3�߸�RB���ڰ�����A��m����<$�v��,����	zt�qzd���&�e���O{���%���0%��M�Ⱥ�ՠDg�-(�8fI�7Kܺ'I�x`.�?���li{�H��r3�*�Z8�cC�/�
���F��7�v�s�g�H�C���ǕT-3������6����r����8�s�lז���h0��Iv����۷��w�V�-h��X4l�e���mG^�h9Y!�,��O�}��>NʲA\s�Xg��6g�
��w�c�,NԿc��X����� ��E��8Cr�v��ւ�'m��h��3�f��,0�l�L�]��#Vv��M�A<��e�Z����ؐ��˫T|8
�5b'٬��J�7S��e��o!Օ\�t[�0�+�јed����şE]J�Tq(3�@���@�ECS�h	�C*O�tGD ���� �{	Q_:�G��_�^5� ��a#doA�!���,�f���+>/A�UE�#�
Z��,#������ �1��K��M�Q+��Q.As|/�%�R�J#s�WoC�H^#A�������'�"PQ���I��p"� ��no��r����Ă�;%�/���,�E�gxR1�/���1w�i�����[��%���_�{�yKWK��?N�x?e��~)X@��x��[~��.仳U�/k� h��ee����D��w�'u�� $ Y��p���	@*�)��[8֕��2�Z6\E�g��bL$3���x��o�3F ~��%AiT��r�)*#cx�<D}� H���Ӫ���dS F@C�j��?Ic5�8&@z���'�a�&˟��ED*��Psgb��K�P3� �4:'��l8����Ϲ!g���/��"��An��3�����?K{��l?0��̋��z�tX#��A���O����Z5���	E?��11�鸝Ey��`��g1:��6�0ג3ڝ�^T�Tu�h��Y���Hw�!|�eZ*�8�������Q���������C�0�6ʭ;�H��H�j�*@z��>�H�DnO�ʣ���{��$��N/`�8]�%�׮��l�w/2A��
fŀ� 9k��+�vp�_#T�� /9o�~IH`=�zc��yM���Q�ğ�Q�|�<���/O�s�FH��i�0��R�F���V�W�("���"����R ��O�-��}��V��OZ`�?�����R~'"��4��܆1��߿v�+"��5[(���y��H��pٍZ\6�[��U�ȜcQG�0</!�x�	���2��p���Jf��}O�3�FG�U;k��b������Yl��	�?�~6ϯy���	���7g�l�9J]n'Q����x���_�k>��K$?�y���;^v�n�{ɑ�J���峲%//C�����V�N\�L}�����ۚ-����[,�W�������~��K�-��F�y"0�A�';��!�VU�H:Q[�O�k�SWV���DgA��
�y����s8��߉!��m�Pf�<��M���}2������a������So��%URE��a9{K��/~٠_V���o�E-&�?�2�a�{fU<m�[fh�溛"wC���*Z|�Q�m?r�\M��c/Sǰ8�]
�浺�ɷ��9}�*�L���#v���Z�z5���<45G97G=��`�w����C� 6��}_k�s�?�b��m޲�����K�a7�Ca�f�{_X�(�u�Yo���a�I�;�x����Wa��a2�7e�� �c�!0�����������s0t�V�Xr1�)��ÄA��1��7Y��I�H8mo��ǒ��L[������u�Z?`yܳA.�C�p�����^:9�PY��6̤��?z�M�k���1�eB�	�P&��P�8Y�<XL�m��\�_�B)n0c,��NŰ�u�}a~���,�X����!>fCc���L���]K��f��'���aRVNXp����v�W��թ����2}��a�u��P���j(���o�U�f�8�9���$��-��*�)�_���ヶ�ﺃ�	[�q}����Z����Ѣϸ.�S�^�kJ>mNM�v�Hv����n�j���Qj-��7��<TR��i��@�]��a-�W/��[�	�5�4�+��=��DΛͺ����bQ7
�.PD�8�rƪIFT!���6]�}-.���M7)i�s[o�}<���ü���D$����	m�6����@�cmQ��q���u��%�GG#
��gQ�j���[�S��Q�d�Gpo��~sn�_3�l�� �=��ʣ��;8Z��+&}��g$��SXq���@��������]k�Vz�$���U�;�)&P��$H�<��F9���`��x���$R�4(�c{�p(`!�4R( 1�ǖ�}6q�?�D���2."���MA+��62q/�<��fV���(�2g���& ��D!�ro^�e��xV_�t	!��8S��qWqkz�EB��D����F�K!{�L�U�]���GUt��z�ߥ�1���c��C���ȫ���t��0��u��=&|D4$���ǚ�(6p~�|}?;�1d浚�x��i����1&.���v�06@��Z:����
���/�ƣ��8t��@(�Y���g���O�a�Tt�`�W�G�%S4q�Q�.��5���L��A�`X���_X�=���еq��~�L+ִCgX��5aV#>�sFG����>`�֔����
4�b��"�·AQ�WcB��ݜ�E��s��Da-H�o���w�cT�2^�d^��(��<���lòj>T����#P�%���+#q���A9�9o*K��A�V��RK�>����\Ca%�����k�j��f+�#��m[�w2�x����J�$�P�j@fݾ��,&�c��d�K�T��қ�y�M��_PnN�l/�E�uu�o�n5��g��1���m�`pΏOE�� e����r�x�u��L'�G����}�X��'Z���Y�hcm[�Β�5P��E��Q�pw]�E�E'c܋e��;ЊՊF��g�L�6*f�W�3Kh=��jY�J�O>�����G%��kӣ'�+|����T}m_j;2#��O?J���ߐ<�:9}mZ�;Md7�OB=6�>��m����Tp.N���7|AU�J1]B
(���5�P�Bk���kGeɟvN2M��R���M|�Q��)�9�g݈��.�o[؃iz�wl�ar���_̑sCߥ�����;��|�D����:K�����"4�
v�}as��@��6��{L=}1!(����$I����G�Ja���m� !��+3(AD@&���I;�k���{TtM�>$���P�=lB�]���S�U�7��=�k�"�.��� ��g�+�1'��������&ν0�Ԇ��Ə�����Yc��BG�V|J�M��&?ʥ!�z7=&N�&�~�#@�=<�ɳH^>c���j~4Z���X�e��Xo�3���ڼ��p���S	=�����6Ɔ��z=4�^�!��;t03�k7�V#�0��&�/����)���X�+vB>+�z�w�Pm&�y�J���x��.�QdW���J���6�FPR�h T���&���j�U���N��O{��YR���9c��Q��nExV ����~���`�S3p��		>{\b6���7��F�5�dk�O�O�\~�QIA��+@p�5Ɛ����,�b��G�t��ؙ>�GW��������}%���<�]���^G���^%�8�]{dH���#ڧ:a�N��UFqb��\\u��a��%��#��L���C��)ST�\�F�W�]��Sp��g�M�= I�	�P��;?��*�7:����W�+~׾xa�a&��?�-�Jx�X�$��� %/�0�F��o��?_��<rZ�$��}����:�I$ADĊO������Yq(�����0��^]w�L#(wv�t�rѷ%�ٴ'YG��s����ϻ;���_A欞,s�7��ln�W4�w��&��S#�/��@ǌ�Ir��_�d���~巙�W�a�&�r�f��^�xF����$*�*��{֕&�ɥo���$��	�l-�!�/�`Ҝ[�Y(���IS����&-�������O�l��Ou��'v�÷��c���j ����(��#����y襜�dփNPFr�Bu�~�,��"����_�=��?+͇�M�*��!���6� �)1酶�@����[0�w����V�:�L����͍���������x	��*�8��w3W���w#�*�:���s�W1^��^��k��`�X�I�����g!EO�J����Z_�KJNP?��?�:�>`�߇� ����"�IƷ����Xe)��h�����ev�~M����}��Ԝ����y+�&�HG�jE�^�nH]y�,Jd��� �����c��~�t�@@��̇j��e_�<���yD�����}t�֑�)�<��P'F�$����)�Ǟ9��z����OxJ����|+�G��(5$?dj��W�8�V .e���3#����)��K*}�f�~G %�;tRu�AW#S�n�;k��v��%��.���%GsRξ�s��	qMi�U�@��l�G�?���R��%�۲���мW��:��.Ţ�?:��j�r��ӳ�����ϲ ���˴¯Ǽ�m۾�*A9���$�@���4� �(Ԥ���}���vB�zBh�&������T@�p/��ډ�R�ק��T4׮��~�;�'�]�9��e-��A�T��5�WW�����sA��r��x�8����s AE3��b��<���2�Z*�����퍒R�x���oz�, ��<��̺���5�;2���Y�U������ ���C���4Tr������7���u���D���W�ªҊ
��sݸ[߹:��VNA܁�}��`���E�~B{=��ob4�LC���3����nnfCk�J��g4룞Y���׫o��]w'qo�O��_���؃�.ݚ8�ߥ�����\}O�&
��@�"ϙ%y�H,Ю}J���{�y��_��Z�9 �A	���}�
A��<j����0z��cM�{��7�Zf���ZI�_���Ԃ����IE@BF��������A��hw�#G��c�_{��E�e/�}k������g%�4��&��Aru��	�\��p���S�bs���&p��/����d�Vp�{W�'�'�� J{�Ӳ%�����KJ��Y�C�ȓ�-ׯ�|!	�8XX�7�]��xh�U����乤w8Kt3�<�~jx��Vx۫��޷0��`bbR�� Y,�Z?Ӑ�(����b:u�A/+3�"佹�Z-�����$�)6�n�$�&�T��}�e��[�m��y��������%��$�i;�,�3��I\HH���v|tE�rXjm�E^~��4;k0�,��t8$.(�||��R[^�����ˁ2�'q�H�KAwo{�9~dEi-p${�\��$��cdnn��=�6�
���CCQJ��$ֿ�f.�>]=^�}��xs>)�Xk�0�#���0<n�·/�G�xl��WUW����͆�Xf���ڈ�9$p�u/W�*�ܙ���#{5~r9����،ߌ�10��v�B�Ҩ?e��U3��Zt�����r����z�i���/8��I�!?���o� Lt��%҆ml|H=�IT�i����m���;��L��#Z�QW��㛿�n!,B�$��y�9��J/�#q�ю:.�}����1\;�S� w��+x� 2���O=C��=N����:����Z�����(�|�٢6J��`��P70��'X��fg��3}k�2Vg��D�qr%����"���s�ԶE4�Mj����+�/��q$W�||��������L�,���?i�ҽ��҇K�#��0��^x��*w5��'���c��oR�8M�G�����ut6<�F�ٿ ���P|R��oVu�=hv{ItRVuF��	�c�^��B�/���LMiO��x��~$X���+����e<�C�'o�����]}�WF��6��]>@�O�D^�IL.����U�W{�(��Q���.ͮ����D��|�"�Z��}��|r�>����tfp5�oΟ�����m�D"P����'h�fzlBB��"�6O^��^<�'<��m7�5�*�2;��V�Z/㥚��i=A4]��U�y�C�c����hD�D�7l�	W|����N_�
g�]WY�6���M���z=� ���%���+�%��V�䃔f���r����q�[�������������n�`e��Ȅ3�,������U�A���M�B��b�w��|\���M��G<�h���r���!�o2!bQD�]�� �qo1���.f��a:}M���SPZh�s�,�2� �:���ǈ���	:����Fɼޞn��&m^�|��5|�I�,�Ϣ���R��O��
_"�~��Di*�i��)N�R��F .��8b�K4�+zT�'zTcv{x�F!�"��9"�]#>�^ՙ�Nss������RCsR���1�qr���rZ\���3Y���3�A�UFI$�4�6=�Zj��`<ǋ['A�Y�rH����>��Q�&d1���%�1�l���2D��q����oN�|Wri��A�%����m���iԜ�zs���7ʎ�����ǯ��<q؛���~��'w��5]�����@��� .�_���)W����UWp�U��#�H������/��QN9$�|^��Xץ9�TP�[ ����z�?�����4��m͝R��1~�.ӡG��U�~G��׋�Z~K�2��G`��C�YQ�ٲ���w��ׂ���Sr�e��/Esz��4.� '���!�k�
H��~�㟹]D�ls���T}>��H���g\z˱Y��`򛟉��/-�.���$�DgS'ފKxo6ߣ!I99p:b�����/Z`�hI	G��#
G�7,&9
�����> ��l��,ƥj*\��n��Ũ%j�=�E�:Z�]���B��Mi�R���~�q���4���Z�w�\y���P�${��ޥ��Xw��*P6����P@`�"��������G�?EQ��j���cr����@����E@R�Q"=�4�Zg�,���Ro`��i�=�ΰQۈw�^y�P����0:�z���VᤨQ��k��°qO=o�/�]����lo^��'�0jL��?��X����/��C�jӌ�z�����q1C��%y����JCĘ�e;�y�3�B�n'YQ Uk����|���_�dC02[?O�̀��ݎ뿞`��#��6��-W�8��]�� �A��i{�����L�u׌��������Ű�9t�g�.[����S%��7���sx11���  ڒ�Z�6�����kp|��P�H�"ȅ�����6jA|���c�a����O_��w2ˣ�T��K�+��'����[\ }��P��pf��;��z�?o���L����g�W�K����7LD��10�ͮxv��O����Dn�+�+�V�d��e��ߞ����K�()��Լ�"�;*6�U�#J��/�[���bIE�
�#�,�5�z��%h{9�\���fÌ*�WE��ï�#[�T��\�`�����x�/�y���q'��o_�^�c�u &�T�w�6H4)��n�>�ڎ�A��Hs��Ʃ����Ϳ+a�z~��c�E��\�@��+cZ��eM�n��5c�棉ay@�?M�&@=�]$����iŦ�Վp�=�/��F�',�xo���\5��K�����cL�Gi�waω�mGϳ�1���6���&�K�?G�~��	����͢zjN��p)%3Y?�����W���GP�^͛G�|��\!��DvP��`�#�~��$pY���C�7PVu��*��cv���=�<��pP�_��1L��Qp�0�u�cx_qE�m1���ߝ�"&5�� �:|�g�Vm�4b}%����ƪ�QZ��0���b��Z��<�R\�������[}���O�m;��(AY-}��a����33����?�SS�r��l7��>�
��p�g�ggZ���:}�D@h\�|
Z��3}*���~	aa�a3&D}Zuoj��e���;������[��s7� ��s����k�����3��q�� �J����,���qPQ�W�C�*~Y�#�9�hf*�p�/菴����|�M�ĥ-���P^����E]>�/˝B1:h�t}�O�_��_�&����X�2�HZ�����ʳ �^vw|�k(� 4��E�܂��C��Ό�0"���NuG�f��z��<y�m���`�>�OkS����DR̗�?��RƳ�J4g��R�R��`�I��F�a��9�<u�(KBI3�.w�����^�
#��.�o��$�;|�R)g���Tm��l�QO�5kŨ��j�l)j�R{���+5��h�VT;v��֎��*b�W��;�=���s����s?���������k�`���������������(�J�Q6gl��_�O��.�^��skJq�Ht!XXI�A�~B��.�o\p8_it6,�C�>�|Ěrߴno;3�O���(��s��-������'�Pc�]eϭ�6��<xFN[�l�^�JAN��B���T�3`<�����Ѓ|2k�����\2���i8��igkZ��)n�����_k0+������.iF���-������ %b�����3$H���~�4�'*E3�bP�T4/��oy�7���'Qi�C�`���DU���:zK��,)^ʷ a��5�69)m����J����([/���󭣀��d�,]�\�[J�-X�g�魬R�爭,1��0�n>���pTυ�o@�d{�!��߽��,L�v��<h%��-1���/�hY�>�KGI�Z�1[e;���1,e����$7�(;�,.�q���F�d��3��IL�)y�N��`��8^gB���LV%��s;9�e����7���N!n��y�wk�s����\_��������;qR����P11��f�b������k} +(߳%2������2����"�,4�r��H䐋��:�$i%�_b���#�HZtoR��9o�Ҵ\K/�jܰ��Ⱦ}_*z���N'�b�����9@3b�!�Y�3��%�(��3+9���i�_��2o:�j	M�8��э����I�קQb�_u�Ѣ�p��I:]�����/���ɡ�qD�97�m�!o�f>*���ޅ�؎�rh��v~T�E�[U�qU'_�\�b|ٯF����ā�z�|R�t@I.��2��!����%ފ��@��j�h�_���;�9��:�K�%H�� |�-0��� ������Iɽ�ި���<�G^����6�i6%��"��v`����4���puM�w%>�������]��Y���؃�9��ң=��O�w��INob1Z§w �jP�e�3����A	��3�w�3���&ƨ��QGR��WϿ�mZGNa���ߪY]Z��N)�_ʇ:	2ᰡ�pr� �(�9P�(4ʲC�ԏW+����,����T�˂W������g�щ��q���n�s�B*�n ��MU'�����KP֧��,�4�7����:�A3��Ru=�$���Q�����p}"P"�q��B#��������0�ɶ��w��yQ}�f ��ը��!=�
(�A�h��]�t��X�+:�g�fa[��[�Q�u�<e��~�K�>�׵��������M:Xy�-�}���{��!�_v�߽�M�G.�+�Q����<dѭ�l�WŷJ�ȃ0a���������uE��[Q)�1�>��L
@���GPcw�1f�]���h���7/jUES�S�)�-���'�tq����Ef������"�r B��'��{���.�6@�g���,�@��Ʃ�MlU9�U.S?��ua1��ʇ���G��sLX 
:��=����1�<�[��_"���&�:���ӌͪ���\���A=�b�C���7%���"�:ܔ�,]��'�K�ݎ���GKT~h�14�'J�VN�2��d�3�	^�rP������;�L�dP�p�)&Dyo�J�8�ĥ�1,��#�L��\>�^{ы�zg^қ!�"4�o�
'!�%�'�@K;'�˅����y����i���};)��3�^�_�� -����|��u�}�d��T[/~@��f�8��X`�j3�!dpAe�sqѸ����\��-l��
��8��oo-�aB���~v6k�8T���v�i� .�n���Y�e6K0���0��KF���a�F{�i��[�2�h1��X���{͛�4����ד�����i�b���1l�^�4�: `&Ȏ�7͟��Z
��ٷi��\����u��)2^C,�@3� ��ev-:�Rwb�BҦƛ�a�<lVx~�(��!y0��������@6"<n��������'#)-��cO�f3�3�����]�loC8u2B��������K���-8I&����7�kx�Ǆ��� �F��Ae��:�s�T���3E���[��%m���M���i��{^�KM�yIC����|?�Bɉ�Y�d)�b��].qt�'�m.�[_��'0/�!a�2X�c'1����w/���ё̟�`���wl(���A��^����薕�^�2���(��B=�P7��c�s���ZP���?l���ƾ/e��iU��2Lj��,���]pD�F���ԊM���` kY�g��5��'~ܸAx�5���jG�ڀ�*�3�VzD�{�a�ʜ>��7%S�J�F�S����o�Xv����K�IHA����#q��wb� �v�6j��9<�(�c�����!�+�R�˯�xwL�j�"�Vu=U�Zi�/�\��^��XQ�R5�nf�=�3��_��7��ܲi�ukg��}и�s5g	��h����?ɮЏ<�O�Ľ�^ %�R��.(����\�`.�0Ր/d��5Z
."��ۻ�tmd0�Ll�MJ��t�:�+Z|X&����.#��P۲�b7"Q �?��:�B�cv��Ja7���T;r��m� N�'OV�$ı��F\�>,SF��T��!���ۺJ�a��S�@�ʔY?����ۂ��N4R�I݆��[�x]�M8?LN�'�߰����^25>��(>;�����쇏�wzZ2" ɩ�ʲƗ��^�)��#��3��۾2�Ɛq(�IW?9	H�!��xÁr�-�O�b0��oL
G"�rX�o{F禵��B�6�b��ve�`�0i�<�_�!.A�?o���xJ)�H���SكPg��>8�ƶ���ɿ:� +^U����ɬ�\�F��9��2D�g�������,)j� T{��|~��,��R�ff���Zq�X��ȇ���;�$�W�T�z�b?®3��.-~�V%�R�5A�Z<��u�?�[��԰H93r���g�/(���P�0�e���@k��I��	���VN�[���X���IqY9,T��+W�|���P�BM��`%.��Hl���8><W»R�7�k�6q�r&5���n.�M���?ҩ�w�Z�|��[fz]�ֲ^����(Pː���e60��`@�u�U/��'гR'b�\���C-���oDU0~��(QZ6$�#������7���]�Pkt�g��o��`0t�a5}�V���dU���Y�s������8��r	]ѥڒ�1~�*�����a�yiw����	)�u��,��[!"��^,1�t�\W(�-RM�Ҽo.Ƃ�l>p^�\��ؙ��
R��<�!���D�������*1(!��7����,�b:w��b|� ^O̼ٶ��)6)��y���lG�)�b_���sv�	�n�g��cʥS6Ĳxf
�qO�o
`�֖r���t�ۆP��)Gˇ#��ٗn��.( Ȕ��9�_B�G6{����`����u�*���n����/�Qy+P���AVfg[2��-s�K1���9^\�ڮ<�����ѫ,�P P���>1
�fB������{��ݢ��@��;�!O k�v}�Ģ_aI\w�ɯ�� �y��GCҔ���s��r�@�=�\}��y���g�w�ͻ�m8^&[k˵��+�~��k2��3ͻ�=�y&ϞpYVv��&ό�i>�#���� ���C���Nb��w^�����}�k�xl�Q��E[���<�<�@JC��5�#5�Gə��pwYއ]|J��L��eڸ<ӑ�nE�ꐫ����g7�ht�=���g��h��߶��b��pJ�fH[}!��1b���4O��DՋ8L�J�6[N+���*��嘮?hPn�BxF�$�ĸT���AL��u��Ե�x�(���S���NI�,����a��1�5?al��T6����=wp�zIDi֥�����MHd��W����A}a`k��f�}���w�"}my�G�r^ݑ�ƪ���N�V�0v5n`0Ť��k�Y�h���/��ut��.�~7ӌ�j�6�����J*��U����!X�6�="��d�Ȝ��`�]������3�Ȣº3�g$�}L���Bo��}�e8r����|2�V
���H�{�x�#X�7�����C���K��3{�;� D����j��C۔-F�N��1fg�b���P�V^������H��t��� %K����t��<�ZLeG��C�:�Fx�%q��=ip{�8�{�P������^��d�q^*�G�+z&sI��W����▷^ ����n�!gb\%FY�U���!�C��������A������\���Yk����^��!	>�X7y����>�XrO ��S��9\���>g�i*�{�i����3SMq��u��]�V$hE��5�Q�Ϊj~�5�2�Gb\��O����V�D&8�^؞N�!=��$�ߊ⧬�W�Vd�ܭe�W���ۚ�40R�E�(��:�˚6;�(j-�(�|�������m���If�T�GF��2���y;ߐګ���S�hJ���0%�=����@�����twl�pX�I�+h"���(�ߥ|m���A��>�q�j~�/���u��%�`�u͹q���9�A m�(s��ux]��Df@T���&�	O�����P�:q�ʂ�N��}uu��+���~�8ж�B֌�{ym��@|k��p?	�n+hD����=9W����̌�2/��߾�s���������[� �3
NJ�P�:L>�>� (6�=4����ƕ�Fa��ܮ�D��$�T���H�,��0
T�?�����U��c�<��7�ml�Xy+9Ѻ��1��`��m�qќ��Aj�BIԇ�rh�)S7oW��i}�싑E8L<7��
q���aF �Uʕv���F��l�Gw�����֫��
����
b���8�խ�E���� y�6��r�l�]�6�JC�[�yD�v�2�<�!})΂�>�$Hȿ����ëTK�� }��פ	�9�-��|��2�Ps��x����m�7h�R�)�����P\t�Q�!b�8��_�3�C]�'��D^i�}bA�D�j�tH������"@w3;�Ϗ��u�|Gx[�Q��@�uQc�X�I#zٽY�����j\v����B9�@�/#3�JD,�)���B6b(��k�P���L�ҙx %�*2���6*�2h"ӰQS����C��)�#��7}#3s�ǞkJ�]��E٬�\L�9���sd&GC�� �;�M��"&\}����Y6Ms�=߯z���/嬕����������f �����س�S0�s��\�>��'��v� ��?��l���+��~��t���N�����2E��Z��\�k�=�`��/��'��)�/�v1#ĕ�;L���F�g��<����u�>'��'��?�l�k��*��~��bEa9�ϴ|�7�xb�\�-�HOh�����r�I�(����9Q�i�!�A�Ԗ*�K͛|�nn��t����-G����j�4ǧօ59V4��%B9��tT����x�\`Eʿ(��.�?/�:%�lĎ����GJ��vnn|8ʮ�}�]��M��ۯz�¤�k������'����Nki`^���w�Q������B�JE;[���D0Iο.��g�m�y�~%z�����U�z*{�F$�*��~�)�����&�Y����Vd�sh����b��售U�2,8���Ϡ%��g�g]>�'�(����x=w_����֒�`�L���V�����X��9��_{��:S�f���P�4�U}��0�(;�*.��~�sZ;��Ī�ο�u�i�8�՘��,GVT��eE�����o�Q��o��!ehb̪�8
�ڒx�n��r��G�h����v�q�q��ϩ��: "�ʓ�����X�j��Z�*Q�
��0	�����2o�WG��1Pݝn�n�Չ�!������4���\3�k���YJ8h��*�������1�^�3
+��s��r�W����_K�����ı��i�+�?z+�(c��D�5 �*��(0��������7W���q׸�h�;n_���k��i�+<]&DN�ֻ�|�͏�]׾�)'��Þ�G��K��6��LPĝ�wQGD�x�k6�$������#
�(�Xu�T��G�?o���� �����2����_�i�<�&�����,�����RK�#r��X����ґ���S�uEɱ$��Ք����C&�>
�L^�V�J�ek�8iз����\|��N͕kݜ{EM����RKd����PN�Gt��V�����g୻>,1=]p����o�㌺��k��7s��瀛�����j�?PK   ��xX.�8��7  �8  /   images/fb58f2af-8fe7-4c12-9116-b892dd7fd909.png��sl&N�7Z۶ͭmlm��-��S۶ml�[?u���ֶ�����y�7����;��LNf2���D��|GE"B���@�����OZB@@�"���zu�s�O :��A@R~��	ٱ,@����]F�]�������
��ˋ�������ي���&�J���U^ZB�w�oj������[2W5��Ӵ�6%�Ĳ���`�R�KI
��������E�Mjd�q�JG
�G(��6<�
� =��2�ݺ�;��w�y���E/;�=f�5��s��}�u��6#���~� 8��i)��3TFP)ϡ �b�Gf@��Q'J�)�`��׈SA�� ������C5����̒�yK�$L�e
FQb�H�	-H�ׄ6U���!~`�����o�2��k�G��o0��9�zp�����p!�2�����ѩ4���MI�L.P� T��u3���0�"��%WO�!�a��fZz��%H�H���K���O�P�&�!Ζ���}ߖ/���v@.�^7���m2B) �<	�<�W�w���YT�in� 5�I�e�p��ҽ q܏�6�.3ndJ���4~G(���o}AӬ�q�Y�;�З���a0�pk���$��"�뱕= m�a�R�m�C.PJե��86B����R�y�ca�IF�4�(NC�If�m��ۑє�nDG �6��$;{��I�OAa��3�Uڇ��R/�ZhW{�CD�D�K4RGv�b�0$�0�Qe�j}=�]KZ�V��1<T���R���Y��gW�j�\�w��(� 	
��خ�VS��ak����~S��ۑ_[��>?@�O	,����5J�JAݝ#���K���P�ed�#�d�Jzj�z�.3��}�#�P�.�w����㲹9��SԚ��z{TFMɨ�a����tP�>7C%50=9�}Lb؝�t0A�^�����:���qu��{��W��<� ��G�P�
�����P�����Lh`g�~������U�O_v7���`�Ў4[+Y�~�-?D,���B����KAP���x3n�0�_����A��Ogt�|rb�:�H��SeG�v�v'�K��:\�N��{&l����ك�f�m"��|D|Er�2��N�^��Q}<�̬·{LT�V�,���ص���J~���U�������2Ҭ��mk�(�v3Ǜ�sfR�D�x��3;G�:R���b���y�L\p�Ok��Sm8���5��AD�=	���[�F:&6[��T�E�R�d���V�se-r�#�F\Q\�d�-���ְ�(��]���E��s�����µ�4*���D�T"r8\,�<���qj#��D&�E�+�{��H{C�@�	����W�0!����9�Q�@`�G܄�ac�U���?��gi
��f�r�>b�٩��E�<���,�j�L�!�O�՗gC9�F��/&D�נ����$d���۫DCm!~���!HI�mų��@��y0]]N����i��6�u��X�\��9�!�U���SE�o���8��ȁP���@Ff]�M[5��I;"q	�jGB#wr��h.���o2��tLR��YKY9�4�6bܐX����p	6���ς��Ws>(�T�:9N>���ϺE�������r�?���1�م��K�)��:ګA?�p����1�O�N������d��ީ��eu�KS��S;Q��n��X�[pYt�׀���
`�F�t�]ϧ���t�<K(MuTO��(��Ԩ��9*IV�9�n��i�Νf)H1���ta���g�RHPW��i�&f�	�~�q;���`AV#�k�αgf�ݩmߋ����9y��,\k�%3�'��Trs����5�=��Ck:����<����VfP�Q�^׻�V��N�?�ɓA��y�7�k?'��j��B������x����W����*��y�%&�l�~27�j�{�;b*f�*����>@/���WR	�WyN�(@w ���;�_S6)`/ju
,�O�?-�o���r���t5���*�跗���5UE��|+p����ᆬ3C�
pd�O�Fb�x�Iв��������ĲBh^`�ze�]:�6��~[#�qO��`@Hg��.H�u6���������bp��é�l;SC�K���������G�]��A���a���1٫���1�{Ux ���.���B���49��Gu��x,��;�@5G�W6�O� ��)�ꆄ;�|/y��K�����N�ĥ��%�*Rnn$�S������U�ѡmkk1]�e��e.�c�pcb��4������8�?�2W��j�=�;ӥ��?�G�,Vk&���omH~�JY�KJ
��G�"���PVF�<7Axv�x��K�M��ߌ�K6�ͯ�1n1c=Z�5ͅR7��x�5^���w�!�u�pw�~��aY=�ʅ5�b I�y �[M����vx]o�Kf�G����a�Y�B\���y^�R���#ri�����u�K��T��N�<��?������{��D�Kc���w�tഩ!�p�C����ω�U-��|Ga���1������?��!lSmmx��)�;-�,}j@�<LO����c@��1���~f���5�,Q��߿Q��J�7�d�T�abL]_NMN�ā���j��1{MF���[�g �7]@�F�X��Rsw��Wp3!tSc`�.|o6r�m;��l/�Kx���}�\1���F���5YO��B����]�Ã�������C2s���t��r��Į�G�.m�B�L_f����!,sSC�{�vx¾���R|��,�c�)���12�,��xSd���x��r�A.��k2v�l�р��Gʖ�R6===��
i�14y-�2Muҋ�)��3vyd�k:O@��|��%�63�HPaE�V�HW<���H�vK�#M�H���x1�� ��ڝ�O�&c��pq�G��Je>P�-K>[뱎�s�=�	E��q䉗��P0��4ip���c9۳����5>���5���Y4a�ط8����hr�h�a���E�d�KWj�^;uGG�+[�������j�g3��~�.�Ĳ�
�އ�0��ro����JSc�Q�*@n�M����F竐��Da�3�|�~=�5�Q�[&��-�}�||�O�ٍE�[EJ���Vk�!���d���?b�r��\�R�NM�u��Q��dᗆ[N|n�c$��V�#p�@7���~�c`y���%c���cS����2��_b'�v�J0Xyd0 ����Twj�b�P�+"p�Z�!���r���ų�x%��cT�bt�
FO�-�(
{?¥�@��� tVʐ1�O�k�V������eWsl�
���'��Ț�G��*l��~��ຏ�p�F�`�����l��2���M�S/DJ���4J欟�4�\�Q�����hhp��HI�~|x�ŶZd]�g�u7�V��ZGhG��F��qh��Z�2�����k���5���֨��Rח�9��Nd���j4c��.��;�m��U8���OV��Xt����K��WE�v�2�OS���Y���M���/&F�����]ı��7oqq�� B�5�@"�>��VF�F��8�є���ǟ�i8��"��$)����sfD&u����Ӎ���G��6F�E���6��u:���%S�t!��G��u�6z�nF���K��������F����L#�^4�܂����ag�.o\�)��&0ci�����M�!l��_u���pQ��⠕��i�<9���E�s���w���uͩ�x�J��R%�̧5R�������W�o�Q12&�<�X��������h�����k��
��lp��Ǖyz#�.e k���ʦt�ZAQ��;��������~Q��oI�z=�[��)z�|WK��*a�t����8�$�W���OH���P,`�P�@��e�Qw2_\�mK��`}���x��܁�76�\�w�6���H�Χ�t����VH�̜F�^T�����$���\���g������c��c��.u9�S�u�sK�� ]���0���cI�:5�-�s�U�aJ�Vq���N�>v���@��y�( �C�@uR��U�p��L��[5��w�7�ݑWW��������䐪F2,u�TuGj_�%eG#ޗ��V�w��o(��)&;w��6bl7���$)ϊ��EX��h<��������`��f?��䷧.{��l�8�T��_+p���@,WE��3�pMv.qjB��l.�d�l`��ٰ��c5�2�=iT]#�($ti̭Dq�T�9�5���X������9����J(�N��$��H�[O!�Ώ��8�FZ��p�S��Pa�DƔ.E&�R��������'��k4�'��)��y-v��m�\�������q�q"��e�~��MNM�O��U�� Mm��,��ȑ���VE�]���E�|��Y hR�*�ꂌ�������x���-m0���]sf�5Y����i�f�B���!~��a�P��m���%i��?��.wC�%�N����b=j,����\UU%d!�U8��COO�\/�H��eh'q8�cR/&B�W�sN�TӀ�.��x�v�*�������ͯ�򕗛\����Գ��J9h^����C{�G^aD��?���W�{����x�.Wr�N:�0^鎰����N�`��%�	�����A�>teV��mI��,��j���Έ��N�Ԡ��p"�j��7{}�=~����aw��ڷ&r������?R�f�Tz>��`R� ���r����3�|Y�U����"��I�-���$�e5>Y�ݜQ���;�@�=��ʜ����������)����]a�pq����Ԣѷ��M%�l,u[^��Ft��uH_�>j*��4��{ݏ���J��F��j��-���T�!��1�2�w
�(�8����wc�2li�|@�qcX�k�ժ̇������1`�����L�X��T��8ǫ�_�xBk�������DC���xu�ʙo�
��`Q3�����;�*ٓk���{�9�
����Q*�i�"���l}7(��L��ٱ��c�NK�I0E�@�XG-�t���ʽ9!qj�o�`��L�	�YZ�8��-s[qd�٘#5��|p	�ҲT�G�М�{���.��ld��ć��0N�J7��@m/>7�#V�ڌ��w�hx2��/C�v��I�-����Wz��O�����RB_�)7b���P[�U���Uj���NK͈�6!��\��lInL�#*h#uuug�>�?E7���<$Nf�P1��݃�F�I�y�
���~loNM�S� bo�c5ڜ�� ���������-�U$�ՆQ��,X��x���k�Ǳ��s��cKf��q�S)��xJ�&?�#����J ��ar��r-w{�w�����\�5OD.&K��G5���s�6aw@~$1��"�K(ٰ�������4u��B�p`a&��y�2�{���ߋ3��w�M�&ژx퇤[�d[%�[���5��a���k�,�;������H�������xt�%���pD9j��5W�G`��dD:���c­����;��z˲g@eX�Z���j�lQm�=�1�3���Ŕo���x���X[�nu��ꓠӡ���r�46����6Y��P.ͫ�zC�2��z$Kï-Q൙���,����t������׿�!��n`	��`/qs�b�[A02��8�:��j%b.ΆU�|�?;�*�[���~�AMm� mָKR���M��Irv��b榯.�i�KO��Yh�
�Z�ݥQ������OOz�<��"�����i�zک��H�{u�]��'�����7�S���-c����}yNTjjnH�N*��x|�ZkJ���]��]���.�������	���m��EH����9�_%K�(Rlm�rM��!Հ>��9Y�Vz#i�|S8����_�k��bp:I�=j^�lX�9�ED���еj��ߒ�6Zx}é�9ʉ���něGK,���0�V�jϵc�yg�JhM� o�r���&AA� S���o�t2���l[�3��rp��d��Or��	����L��n�,�:��qE݈�k�L���>K��m�%��w����>$V4���p҈Iu��)L�K��̱/pO_�n׳�p����:b~�cE�F|�O�m��)�����ј��8J�]f��Y	_!��Y�4���)/��k�Dio2�np��B����f���2�ra����(���E��'���
��+y*���!�F\@'3ώ}�-t����y1�1h!5�E��v!�/F�z��'���8'�h�Eb_�~dq��2��
�(�q)l��Jx��m;�������]�ܬ����0���٘Qք��A��%�Z��[_Fΐu��p͝闃庉u񧨫�v^��W�A2��X�Y�(���x��k��� gb��+[M�3	ä��뭀��y�P��Փ}���9)xu�lp�	���n2x���WDt��+�vk�?G����n�S�9���%���{���`z�mN��Uhqu��Â~�f����~q�����}��x�?��~7��3K�ε����[�� V�ԡ#�-�;���#6R�c]�&�w��_8��e��bE��������Z�N�B$܋{�?�$��m^�"�X
l���v
�~�B����Ҍ�?C)\��Q�:���)ӓõf9�+��#��f=i�`�/jw�?���?�qN-|�U�!5V~b.c�G�A���G��,����B����`�֏� x�_},Ш�S%ޜ��%�~�q�,T+[@K���)�F,a�Y��E �Z~�\Љ�7��a^��ȺexN�J�g?�8�U����B(>�P?Rg���I�N.���(��5��u>�I�]4����6�>\-�?;/��eB�~r {�S���0� q(y�P��{�{Di�.�"��H,9o�<p jjE�������CKn\�$3�L�����!~�G�0&�@I��Э��E4���t����0Ρ5'��wqqm�Z��;�Yq/�0�Z�v�wK���Qz�o�	��m�_��K��������}� C���e=p�M�k���K��׿\�� &3e^jU��-NI�J}��I/���ikT��(�ΔA��Ø�I�.4�l��(O����		+}F���ܩ�����ÿ���њ-C�*	�T�g�yw9�ge{�M�J�2��֖և�����Rt#�qoՒVG���k%�J=��M)xߐ�:���9�
����M�(F����JK�Ѕ�@# 퇯9`2ն����S03f+�(�{��C�סK����b<���4�Ph"י�D[� ~Y���[sa�:l��"�� ;�!B�-�cR��K\o6����q�d>��d�l���O���L�����y$Mq�eN���4J�P�7ۅ���<Z:2~��|��{����f&�m�h�a��m���QW=�s�0�)ﻄZ�A�.���Gث`�� 9n����ۓ�F"�RZF6���q̃4�E12ٌ��zvr�u�)�^Э�<}��H��=Iɶm�� [�+-�C5�>!��D��~z&��x�A���bq����B�]v��yip���Nʙ���Phm�h��;��'Jb�K��-��M� �Y�ͬ�f)n9H>$p�'�J29H�YmB^�3.|�Y��v Lދ�`3�Q�@��
�*�~��2��E�l<0p����i�v��_H2s-bEbG,|)���3�P"?���0"DOO��&/�z�ս����R�%d֜c��� �I��!:Ww��P��r�Q�dnuX��%������7;vbKɜ�7�kVX���Z�OL���U�zx��������L���5Py�
�r�������^��6�z� �h�蒑Z ��I��k)#��tdc3 @���Q�&[��ϛ	?\H��l�J��#���ʹ���7��{N��[{�a��N��ai(�<


I���=N�gCW"�rU���KXWo�~�&G�<Ys?�I��� ���~l{��"�yT�>����Ͱ�	��h�~#&�'�̸�C�6���W
:�7;�s��CF�	��^�c��I`A0�/O�!���\�ay�6ד{)nr�j!|�/V�{ٓ ����Q�P�d�42���\�٠`L�V��֛`��3��%�o������))�D,�a1k��7o�1͔�`�N�˕u�E��@��T?Y�!���n=�`�DL��&������O��8���_Ֆs��:fO�eL�ܧ�"����d��s4z�'�}�;�8Z )�{����Y&�~2T� SC�P�H�;�t��9 !�����4�P�%G�H�F��(�h~�w�1�ݐ�
Mj�{����I�x5j��zϋ'o���w�9��wZT�K*q;!u_���ԁ�l�sԶn������Կ��Lc��$��@�HX�l���D7����I�B���Ja��|ء�ʇ	/I���������X��O���Y�L������l��(��PK<��݅�=9�-S����¦;��i$)��Z����4��\ϵp+�1)4� ����{,{�M��lc�͇�Yy�ʋ*�b^
2�5]I����N��!�N�8�8_�w�g�ނ��N����*��zN!f���/Db�M��<����/g��@��&�a`a��ٰw����(��v<��L_ZPh���e����/�ۇ�顸�,�������L����]"Wz�պ����o�.�"��Dn���\����]F�z�ﱳ�#��O�d>."f�E>)��}��H�a1[�A�|�p����˹�w�Z&6M���������O����;�J�
p��%�ckbɠ;��a�d���>�������')����zҞ�!�\�4-]�DC�o	s!�o�ƽ�K��ao.����98|�2�z `��+����D^���V�IE�_0��`����'}
�	:�* ]_`1����>�D��O��5�J��7�����49_��ݳ��(�~�G�_��r0hGuBd�����z�����iz��.�]�<�����Lc�6nN-�C��]x���F�
L��96���5u��j7��^V?=�ߺ��x���m}<��g�����򯄣����J*'h�3����(E�q�"��E����oێ�8­/�|f��Y"�V,������,*g�2��@����� �N_�`���qndњ�Lk}�sg�\��h���&��+bx'o��*Mŋ=��(m���*"����Z1���������q���L�#��I�Eq���Dŧv�F��¿��'�e�y�wc�9������6Tpq�<o}���Vt4���-���v;����#"Z!�]�L|n�wU����w��.�Nk��������ȉ�Ǆ�����*��-���:F�k�J��C^����}oK�@7/��-g��{�oN
h9B��m{m����Ϝ__5o�U�e��!�M4#��_U^$S&�S�SCn	�ƟO�rCP&]��Pj�%��[�2����'\����W�"�`|#B�����z�CP�N���>.�6ng}�'V�|�Ӏ-�~> 2�f�уI.���=��H���z���`N#sz���OF�Y��/_B�3���:�k>�O�����s�Fkm�7S�/��ķg	x��ہMs�����jW~uD^
�骥 5���oA��TF��B�����S��hj&(k�{�a�x-(h��^v?{�>�����i�m��y]��&	��қ��4� Oȵ_.]b�"�l����� �'�}m���Z[>&�|͠Y���y����A��A'=X:N�{�8�`<��X�
uHF�h�_��?��*̊�-��`i����K���Չ$f�(gV��AGh�e,�>�V/\�r�9x^~����ǴQ�t��=)t�j��i4�D�~��O*�=bl��jj&@u����t忴v< ������/2�E�:�z��Ppo�s��lR1�?v�f�I3�����L�ZqyF|��@�ǅ\�������?�ֽI|o�B_֟u-.��%/a��A�����%-n>��F�s���%A#��4X����κ�#\Y��[����b�A��㢎�Sߙ8~6���	dIB��N�|$1�b�澅��`�#�8�S~?�n�Q�:���$�#�c�H$nY�|���ѥ�RW�q��.z�,����)0���ʴ;���u6ĕ{��^y�B���%q/�m���F�+�l��#iL��E��颏���'�ҌQ���<Q�<ZTfm����	Os�]�A��+�Ǽ.�o�>"��隃����6~_���w������ل��Bq!��v�_j�vq�U���yy�x�fg��s�����o�Q��7ꉷ�������Z���"8�C�ϓ�\�ǅ}oj��-|x|��o����H��ńf��3�}F��q�f��"A\���8����b�����]�P��FϪ�V��|L0r�́����ރB�_B���h[���n=���F�����Ķ�n��م�ы�h!Y�(��׶�F;@1Im��?KbѪK���2&A�͗~�{��\MYd���M�Te�滭�� �5������ �l:�j���C��*p��hɾͦ�,tS&J��?gf#�a<G8��?F�����'�-�79��^vn,��Gt�loʸ�i'c>U�[K�<�m�DJ�>�m[�N����y"��X5��d(U"��ڻ�ىa��;��f�~h��D�m��X���jZ\�=�؂��%��>��n�4k����r~秊p�����H�o�^i��Ø1'�b�>Y����iNm�g�K��}5G��'�$w���B�r�_0�%
ٻ9JM���F�p���p��*��L̩�L=(�����5I\�/�9�ڒ�e������SU���rc�wQI����?�.L\pS����Cb2R�[q?��~$���`x�V*}	7�[DƸ� 1�a���0j�U��P`oR>聄��N���ع�Fg}9Z��ve�ҩ|`�'�!�����i�]E�;��D��\a��L�M}�Lt���;��e֋�E�9��ݔ�Ɍ1,w�Q$v�XA�i����ac�"zJ��'��"�k�aZ5M��-�7��wq��+6���=�@�4��"=1qP����Hֵad�É��)(H�;oL��P �Ŝ��;�Kk��;Х��ד1�6���M���m�F�e��jP��dJ���A��Us����#�&���IRc��b�D�K�����J�i^<zolc��2��	���6��'h���i+@��Sx48F��*by��~OO,R���&��!-��B�����d�ڧݼ,���CS�gӨs|_��G|�]4�����*�{m.��;��C�7F�@�-;�/&�X�i%����;�����o�L���#	ADNF=\յ���G���Ŗ�Z[?��r�y��]D��!���<�?��^�yq��䫳.�HC�i5�Z�I�Ș�<�)_�W���'Ъ���?LcҰ��Ɲ�+���b�y��5��#&�^��1I���Au�z��tP��D>#�krЂ$���5q���0�M����JYE&q,��^�8E��%X
אT1a���&-q��~'l�Q������t�m���'��r6�K��t�,	מ�}ݪu}ȆZ>��Z�tٶ��;�K<��EL�5*�Y����u��ׅ��ڟm�@/o�[�=+tL����y�����D�{^v�Hv,�e�qw�ب�Nؙ6��U�9}�Bd�d�-(P �z�0�`�����m�{b/����t���jR~lQt���V"E�#�V9�e]��h����wr)̕��V�f�o��1���Ŕ^�T=P�'�v-�9�v|+��}-���m��X���I��E��#�^�YV�z������Q���� ��l
��.�p�M[��
�Qb�1xEV�g ���l�.fS�Ԁ�MAj�I��Å���t�ϗ���d��O���n����_a�T��U=�R|6�(g����}�#�I��ҝ&�{0���U�h-��$U����yn�T��1�C�E�>�H�X���!3Z�B4�X�hj�Yix>t��R��
9ad�.�Qɩˢ5"��/��"Q�>�)�ρ� 5a?�|���gbuV�0��ۣ@�Fh�M:����(����e�L��c�=t=G �'�?�0�h{�^�r���`!{���)!F�6h1=#���< ��yMY.�Or��+�mJ�� �	�JG�*oY�&N��:k�ы��I�D�@}�c5I�x���)O��x�Xad��X��>�m�����U�Wg#@��C����:Nݪ^�����Ӏ����x ����X�&}����!+�'s*|��cM��G������#t`�<3�XE�{Z����3�Z�n>j�`I���!-��I�U\?�yq\(�k��!��t韠�#m�̗ZmĶg*��|��� ���� 9p|f?E���ݎ�M�$&��2_ ��{�+�b?�,oat�)V���%N*�kp# ԕ:���XpU��='2K��(V�jPce�E�Dk�Ú����E)<��Y'VI*>ō����0����R�Z���3�-�L9}�|%��ڽ��jR��Y(04 ƤVV���Hb����e��$/2ِ0��r�ާ�Ҧ%�w?�wBA��
�J7������i�����1%@F���e�9\�ļb��|OD�{����1���1��L��E��&�fV�k��@!z*�h�|�N�C�NZ�>�:+Qğ���;��Eܵ����fo஦׿��m���q��HJA�A�z'����ݧ:�X*��C���O���t&4 3y��O��k9qCw8�:|n0u N��}����oW.0�Cd��1^1���U50��u;S�+�oh��E��#�|����[���J�@�&T[ϸ��20�}�V@�Ӱ {_�<�9.'��e�.�g�|���ޤkԣߩ�(~[�0to0��0��sՒX�	�?v��3�[���]m�U�9�}Y���I�q��/��I�F���F`�εs�`�4���i'6�\�+�v�=�Y�k��U۝S=�x��ks�Rv�����
�%k9}�z�yl�x�S8�S��:�������o��)�S���ePT�~{�J���$�A���=��eˡ6.����.;rAa��H�1<�jD�}ïa�%Z:�5���ɒ�p4��r������
[��K'[����	���/G��h�����ⲃ�Q�{�yױ����T��A�z�}�[^����[ѳ�Ѣ�Ly�)����i+�~��!�?+1��8�&��z��W�gբ]��N.��̅D�	�|�B����)����='5=������ֺ�#�=g7v8�>�����`u�|�{���ٖ��$�S�R��ߏb ���[#�����l2�B�T7һ ��\��w� @��6�f���{\i�OI䘖�ۿz���/�Y-AɈT��ڸ��{��Y����8�,�}����*Xم��_g�����LY:�l؍��L������ɚ+lxwoc�g�y���V^�UN�D?	/���΀�B_�~Y��$�E�S߉�B�Ȼ�qw��&8Y�R�ʭ:��>���Dr9�a��k���Rk���ԭ��L�p������zQN�0I_�dځ41#qK�����)s哇��×*J��,�x��X�
G��[l��۹�B;��X�Qȳ4�{�m?+��B���2��2���w��g��}�>?���,5bu����P鸮��Q�k(�dE~�n�Գ���0����F���*��{���'@��}¢$洐��xą[kJ����Y���~�xx��.(ƷQ�RY��h���N���L )Z������2��X#q u�j�����vA��tkkN�ۯ�m�ip,+t=���d�]���O�ﮫ�~樕�&�������c�r��g�ӡM�Z-pn�d�0a�ڽ<{<}���/
_��W�;^��J>�b���̸�Oo�y;������S^�G�.¯t�IL�q�����E�r�j�n#)�GF�!��zKW6a�z�5���_P��-!��2*����!�PK   t~�X�2�T]  (�     jsons/user_defined.json�]�r7���>y�DH��F��1��Dk���@� �w�n�ٴ���oV��T�F�\{w�����B�����v���"<;����w!��;8<�%�.����6�a��˫����������?�ݧ�����礼}�^���b�g���r�¯y�?.W���NW�7�Nnl=���2���qGu�H�R��yM��񠝶��¶-'�ү���n�v�����
�	��V�b)��R�!���ŏ�����t��~;X\}:�_^��_���}�t��Ѐ�����s�;ۀ��^#\������+l��{�^�_a����o��9�D�h8c����?2�<Z���+������
_ʹkC�������� ���Ti�E�y��g�N��Ň��i=������߽���>��`�����������?l���ڟ?�W�\��Vˋ�Z�o<���/��c�^��E���������	�R�=�M^�x�O��o��Ow�{G�0������g�����������t�����jV��_��?��Z<�m|#s�\\�������;�xb�e��n����r��2���1�\"���v��<��w�����I&M�4a҄I&M�4a҄:M8�\\]�׳ǯ_
����j������י[t���Z�.S2q�բRX�(cAKeK���8�I�j�DTܲ�Z)@)"�QD(ʉ��2�æw��B)T#)�I	�n�ͯF
��r�U~�lc�?e�8}}6B(�:ˢ��������7����� -�Qk�7*��C�z��Y|9�#�?��~J�J��v���������(��ǖD0�K����&�4����$t��MB7	�$t��MB7	�$t��MB7	�$t������u���?{�\/W����/��n�;���j�o����DF���P���0bZ
HQ`T�ZE���%匈 P'[�	s�FZ�v�h{��r�V�_c݀6�r�(Cu��a��>�1���X��2��)K7��ΥT�fl?�k���.�m�/�c���v�'.x�ʊ���vl?Uَ���wT�$�"�@��(T�W�O�_\O�j�/�]��jI��#"2J��-��4p�:�N�^������|�����[���F��Ց�-�D	�:�F	�q���*gv$��U��w@ �_B�~9̾��k�4-��Ì��R�(n8���0�M��\�F	�O��L5���;<|��	�ar<�qU���#�&��@�?i-m	�-�g-`�3y�乓�N�;y�乓�N�;y�乓�N�;y��Nk|��hF��ۅ-�&*�\�-H�A�d��#�+�bh�tDH@G��%���z�	Ӊ�w�}�J��w�v��8-<��9c�;Mo�K�j�Ri~7W�X*mj���s�Ih՜r�c)cev�K��m@(���V�w<���:k@�@�l �g�=d�M_�F�V�oE�J��g��DC�ao�Z샧y}J����������,�?@�Q���(�=�������Xn)�'vF��^��X���P�����r>{��1;[9�l֘��L�hW0Z9�i���X��� *2/t˙r�A�&Eeؐ�u��AKZn�^3��]�-/_)g2�.l����^fE�C�  ,:�Kq9*�� \k�h|�3N��9�]I�{ta)���9j�Л��bO�7~��c#{l���"11hL�EF��X�:;Km6��D�� A&�L�2d"�D�?� /�Of�p<��qF[��TD�Ȉh=�VHC�
[�\�:7v��q�e�����%�ʖؾB�.rFc��_����$���/	���#Q^�4Z5��_z0˰ e��� "�j�h�m4eZ2�x���J�K���5QH�3�Y�@�a��v�TZ(��Ml-�g��Z��>�\�NF�NF�NF�NF��	>̞��:�~�}�i���.�~����]H+�1�j��&�@���-�QZ{�܆�UZ���%к��ZK�Pu���
- ���IiО�<$�Q�p-�:d��rm��42B�]"���;t�z|��o��"����!�]�tĀA�ށ�mU��w�.~	�>Ƅ٫��+*w�
n�xg5�Hdgfj]!��H�|Q�k�ޚ�u�:��c݂�h�E:x�f[�yҫtc��p*Io6�h���)G�E�;t���|LŐ�n�������%���Z�B�5ܗt�o������T�<T��c��g
���5�ط��Pk�	���}_d��+FX�X�1jP�:$��B�Z������)�(����������u
ňkl���o�'��Z�c�#)Jv��J��������I���:,F�<�#�O(3L�����p'�݇��Hi���Ҳ0���d��j0[�@Zh��Cٖ���v'.��^|'�ն���>�����E	��!�����r������'�N��`Z�l�'�e�� m���>]���G���͉'��/aW6�CM|�)�7B'����1�6>J]��CMLY�TX1�"ڶE�� ���^[�CM)�n��/�m�U	��s�c8{�P�i(:��������2TH���+^9\r�f���l�_Ԓ��Z�9��r�D~a�0��g�	^o#�v&����5��{��p�z����jk�����Ć�������D)�$���50\�u�@�K:]�y�K<�B�tC^�3!�M�Z�%d"ϹĂ,�٭�ZF�X����Yb�f�#L�k6����N9*M|-�8�D��}�Q6~��e�\���ϳ��0~룚��Ll���(0XZ��R"Y`�a�����'�����IT��Xshm��Ў�~D���B[�9,FÒ���%���o(�^#���i1OǸmt2��F3�m��vr.9fݚ�#���u_�CIbI� � eV��箍�Ib	+��������c�;w~>7y˴R���Q6V6�J}t�������t��U�V_[�"� 8C5 *d#$����̒�S����*L�0�¤
O�
�,Q�G;k������PX�~ц�Lu �'_X�)�,���H���8���$@�[+����V��
�Qj��?�(*b"����@%����~?�N!) ��6CS#��OiK�D?� EW�s���˿���3�4����1q�	�kx�U����`�l�8�[з��V�?bo���S� ��Tt�h4��0�X�<��o#8�m˓���SNZ�4��(Nպ���tTڠ[�@u�����	K����{�i-D�c�Z��ۯ��$�(Y?G)�H' /c	k@����L	�j�9���?j��������qL�c��񡔘�0O{������0O��TXM��TXM�0�¤
�*�TaZj1-���ZLK-���R�i�����G�3��v��>��]�v�%c�0]��3�7QXJ��ę�NR�-�1�ef�;Bi�a�E��5���Z�����!1��=p�<��an-�C�Y�6r����x�������T��n�]8�j��;xY�W�o�E5|^R\�����^���R�� Tx��ŋ�c�Vk଀?�����?9}7&��w���՛���V9�������F 
)VG3 
�(SGS��{�F3��Ob��h|8)tp"��e@�����������3���^� 5x�E ���r�������Uw5_,g�nR�.�y5��%�m�Z��'�����g����B��X	����2k�h�;��0�e:@Kd���~�oAxM\��Q�ow+ş��]?�3����'|�=�-�I���g\�CF��uq��݋oG��Qw��"ljd�
���%�rU,�0&�d�
�P�%�hLf)mICl:L�V�n�g��Q�k@�x�B���.fa�#1tZ��G�q��hi���F�:�?ʏa%�<�s�#9&��:�?Rc:���#���:P��W��̓	�k��p.ސR���Yala�)^��,O*H�]������u�yZ��V��,�+�j���=�M�H�k�eU����%�	��Jhf�y���h	��Zh��Y	:�7��ֳ�{�-/8s�x�^m��
�<�@Z/���Dl���[]�ND8]	Mg�>�u����j=;+!'b]5q�~�#'^-oxy�H���(#'r�Z��2r"��%�*#'��Z��"�Hl��!�2r��Jd[FN�m���2t�v��Ь���D-t��"Q��Z�2E���:�R='Rw����*z��C�������V����}��z�2�����B���Z&r�UV��#�L�=���|q#9h��+P�ŝL��=��@�g�2�y�����[����[�D¹��_3��B%�,T��;Le������{Le��*��]�2c��.S��
�A��T�b��cP��Xɠ�e��
�A��2,��AY5$����
*��VF�|5�KLheT�׵:���VF���N,'��Q!?:��HheTȏ����Z
��X1Bk�B���DhmT(�Wby��
��Ы**z,ï����2�!XUT�w��0�**��d(V�]f2��
�.3�UE�B�eXV��<��~��&F]��'v^O7?��/f�=�m+,#��H��q]tD���:��S���;zv|���������iڅ(MoKy�E$�JG:���	!`s�@�ᾭ��3�&�EҲ�ń�B�c�p����/,e�Е�j{z�����|?����q���s��ӊS	Pi����ek�W(<�P��D�Qz������j�!�P�d�	���ր�6Px�a&�5`*��s��[m������F+M�"��d�e�.>E�.�jū
�	T���R��}�}����gŞ(�*P��FJ}Q�[��t��U���u�t_b��X�+��I��ۅU=�e��-Δ������Kd�4��OP s5~�i��:h������s�9�.L��:b[�I�:i�V[�t)�qX�Os?;v��כ�8r��&=�y�������X����0P�3u�^��4�{�����W!��:B��� ���G�W.<w���L�p/_ߛx'.��a.�;q���hM��)�V�hC+��i��C���0��2w`���U������輦���[^����΍+����s�jz�>�ows�2Kܰ�X��r�����8m<��y�$�v:>�?��?PK
   t~�X˜��[  �e                  cirkitFile.jsonPK
   � yX<��)�  �  /             \  images/04ddd2dd-6c74-41be-bfc6-e572c074e241.pngPK
   �yyXL�4A��  ��  /             ;s  images/1697c656-98e6-4bbb-a2b4-f12a22fc7906.jpgPK
   yXv��^}%  �)  /             �e images/16ad4ddc-6952-449b-a843-6c6b0f91f705.jpgPK
   t~�X@�Ǿ�@  �@  /             P� images/20309cfb-f1e5-4537-8027-12bfe73d577d.pngPK
   t~�X�u�̔� � /             F� images/266cef04-a032-4603-9423-684d401d8b46.pngPK
   �yX �Y�9� v� /             '� images/2a0872bd-f672-45e8-b778-ad7a0f52371a.pngPK
   ���X���l��  � /             �Y images/30131ebf-3f05-42a3-9ad5-e2b3b9511573.jpgPK
   �yyX���Z��  f�  /             �W images/34701e0f-fe0f-4ef5-a5e5-12bda4ce8831.jpgPK
   t~�X���!R  R  /             �M	 images/38c30459-3482-47ee-9b33-edd591009797.pngPK
   t~�X\��䓝 Wt /             c�	 images/4809d2c9-d031-4e44-9b5c-1a8b0048f1c9.pngPK
   ﴵXJ%z�� �� /             C> images/596a7037-fb63-4077-b806-d059e7ba626d.pngPK
   t~�X���  �  /             e images/5d57974f-fced-4f10-a93b-7d150e366d9f.pngPK
   �yX$�:{� � /             �2 images/5dac6161-a6f5-4ffb-b809-ec8007c48853.pngPK
   t~�X�z��kW S� /             d� images/65d233e5-7445-4b75-a6a5-2d8c2ad1af28.pngPK
   yX�%��7 �; /             % images/67e1ca3e-4bd4-4ce2-a74c-9273116ca70d.pngPK
   ��xX��MY��  �  /             ] images/6959c78f-01fd-4792-b095-b0ffc5233e8e.pngPK
   t~�Xq����� W /             e$ images/6b3c47ca-37ce-4ada-891d-054e310e4230.pngPK
   t~�X'�%( �J /             x� images/6b7f4d85-4146-49af-b1bc-6149946ceff8.pngPK
   yX�_B�   #  /             ��! images/6c59188e-af72-47f9-a95b-923959af310f.jpgPK
   � yX��{	  -  /             " images/84b7793a-00b6-41f6-9ec0-c4aab3fc9029.pngPK
   t~�X�IM��  � /             ]5" images/86917e2b-5e70-481a-b4c7-aed39e2d087b.pngPK
   t~�X����H   C   /             �/# images/8e6e9996-4250-48fd-a42c-980e5b13088a.pngPK
   ���X�O����  � /             EP# images/90427f57-b7b1-4ef6-8fbd-3930b2051391.jpgPK
   t~�X$�8  3  /             yO$ images/958920c6-b990-4f24-a78c-97ace316bd7f.pngPK
   t~�X��) oj /             �f$ images/9b962a8e-14b5-4317-8666-1954827ef6fe.pngPK
   ﴵX��ڙQ� � /             h�+ images/a16cea49-f54a-4dcc-9abe-0eb2facfbaba.pngPK
   ��xX�@M��  2�  /             $. images/a83bc8df-a6df-47fd-a18d-828755ca269b.pngPK
   qyX�u�Q�"  &  /             �. images/bf545c77-008e-432a-b90b-35b3da31b275.pngPK
   t~�Xp>r�  �  /             8�. images/c13bb491-011f-4ad1-adfa-58d33d2d83a5.pngPK
   ��xX�Rr5�  5 /             q�. images/c34e957b-2bab-4628-9db9-846c7013e8bf.pngPK
   t~�X�|�	  	  /             �/ images/e1d4e862-170d-4bac-8b1a-e4319ef50e6b.pngPK
   qyX5��<O  g  /             ^�/ images/e63eccd2-2ed2-47c9-a1d8-30adbe2258b3.pngPK
   yXO4��~� � /             ��/ images/ece94f61-988d-4529-a2db-f0bc9c1368d4.pngPK
   ��xX���A�K � /             �W4 images/f32ea318-bba9-4379-b39a-fc7186e9eddc.pngPK
   ��xX(	��I�  &�  /             ˣ5 images/f33b8d1d-9a3f-420c-bb18-27c74f47ec1c.pngPK
   ��xX.�8��7  �8  /             a@6 images/fb58f2af-8fe7-4c12-9116-b892dd7fd909.pngPK
   t~�X�2�T]  (�               �x6 jsons/user_defined.jsonPK    & & �  /�6   